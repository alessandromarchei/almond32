
--    # Datapath of Almond-32, a 32bit DLX-based CPU 
--    # Author: Capozzoli Silvia, Marchei Alessandro, Terzano Tommaso 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.myTypes.all;
use IEEE.math_real.all;
use WORK.constants.all;

entity Datapath is 
    port (
        -- Logic signals
        CLK, RST    : in std_logic;

        -- Data signals
        DATA_IN     : in std_logic_vector (31 downto 0);      --DATA FROM DRAM
        IRAM_OUT    : in std_logic_vector (31 downto 0);      --WRITE INTO IR
        IRAM_ADDR   : out std_logic_vector (31 downto 0);
        DATA_OUT    : out std_logic_vector (31 downto 0);     --DATA TO DRAM
        DATA_ADDR   : out std_logic_vector (31 downto 0);     --ADDR TO DRAM
        BMP         : inout std_logic;      -- USED TO REPORT A CASE OF MISPREDICTED BRANCH FROM THE DATAPATH
        STALL       : out std_logic_vector(1 downto 0);

       
      -- ID Control Signals
        ID_EN       : IN STD_LOGIC;
        RF_RD       : IN STD_LOGIC;
        SIGND       : IN STD_LOGIC;
        IMM_SEL     : IN STD_LOGIC;
        BPR_EN      : IN STD_LOGIC; --branch prediction register enable used to turn on the BHT
       
      -- ALU Operation Code
        ALU_OPCODE  : IN aluOp;

      -- EX Control Signals
        EX_EN       : IN STD_LOGIC;
        ALUA_SEL   : IN STD_LOGIC;
        ALUB_SEL   : IN STD_LOGIC;
        UCB_EN        : IN STD_LOGIC;

      -- MEM Control Signals
        MEM_EN      : IN STD_LOGIC;
        MEM_DATA_SEL: IN STD_LOGIC;
        LD_SEL     : IN STD_LOGIC_VECTOR(2 downto 0);    --USED TO SELECT THE PROPER CONFIGURATION AT THE MEMORY OUTPUT (DEPENDING ON TYPE OF LOAD)
        ALR2_SEL    : IN STD_LOGIC;
        CWB_SEL     : IN STD_LOGIC_VECTOR(1 downto 0);    --CONDITION WRITE BACK SELECTOR
        
      -- WB Control signals
        WB_SEL      : IN STD_LOGIC;
        RF_WR       : IN STD_LOGIC;
        RF_MUX_SEL  : IN STD_LOGIC_VECTOR(1 downto 0)
    );
end Datapath;

architecture BEHAVIORAL of Datapath is

    component REG is  
        generic(NBIT : integer := 32);
	  Port (	clk     : in std_logic;
            reset   : in std_logic;
            enable  : in std_logic;
            data_in : in std_logic_vector(NBIT-1 downto 0);
            data_out: out std_logic_vector(NBIT-1 downto 0));
    end component;
    
    component MUX2to1 is
      Generic (NBIT: integer:= 32);
	    Port (	A:	In	std_logic_vector(NBIT-1 downto 0) ;
		          B:	In	std_logic_vector(NBIT-1 downto 0);
		          SEL:	In	std_logic;
		          Y:	Out	std_logic_vector(NBIT-1 downto 0));
      end component;
    
    component MUX3to1 is  
        Generic (NBIT: integer := 32);
        Port (
          A, B, C: in std_logic_vector(NBIT-1 downto 0);
          SEL: in std_logic_vector(1 downto 0);
          Y: out std_logic_vector(NBIT-1 downto 0)
        );
    end component;

    component MUX4to1 is  
      Generic (NBIT: integer := 32);
      Port (
        A, B, C, D: in std_logic_vector(NBIT-1 downto 0);
        SEL: in std_logic_vector(1 downto 0);
        Y: out std_logic_vector(NBIT-1 downto 0)
      );
    end component;

    component MUX5to1 is  
      Generic (NBIT: integer := 32);
      Port (
        A, B, C, D, E: in std_logic_vector(NBIT-1 downto 0);
        SEL: in std_logic_vector(2 downto 0);
        Y: out std_logic_vector(NBIT-1 downto 0)
      );
    end component;

    component PC_adder is
      Port ( A, B : in STD_LOGIC_VECTOR (31 downto 0);
             Sum : out STD_LOGIC_VECTOR (31 downto 0));
    end component;
  
    component CWBU is
      port (
          CLOCK : in std_logic;
          ALU_OP : in aluOp; -- input signals to select the operation to be performed by the ALU block
          PSW : in std_logic_vector(6 downto 0);
          COND_SEL : out std_logic_vector(1 downto 0);
          CWB_SEL : in std_logic_vector(1 downto 0);
          CWB_MUW_SEL : out std_logic_vector(1 downto 0)
          );
    end component;

    component ALU is
      generic (
        NBIT : integer := 32); --# of signals the CMP can generate
      port (
        CLOCK : in std_logic;
        AluOpcode : in aluOp; -- input signals to select the operation to be performed by the ALU block
        A : in std_logic_vector(NBIT - 1 downto 0);
        B : in std_logic_vector(NBIT - 1 downto 0);
        Cin : in std_logic;
        ALU_out : out std_logic_vector(NBIT - 1 downto 0); -- 32-bit result produced from addition, subtraction, logical, etc.
        Cout : out std_logic; -- carry out generated by the adder/subtractor
        COND : out std_logic_vector(5 downto 0)
      );
    end component;

    component FWDU is
      generic(IR_SIZE : integer := 32);
      port (
          CLOCK : in std_logic;
          RESET : in std_logic;
          EN : in std_logic;
          IR : in std_logic_vector(IR_SIZE - 1 downto 0);
          FWD_A : out std_logic_vector(1 downto 0);
          FWD_B : out std_logic_vector(1 downto 0);
          FWD_B2: out std_logic;
          ZDU_SEL : out std_logic_vector(1 downto 0)
          
          );
    end component;

    component HDU is
      generic(IR_SIZE: integer:=32);
      port (
        clk   : in std_logic;      
        rst   : in std_logic;
        IR : in std_logic_vector(31 downto 0);      -- address contained by the PC
        STALL_CODE : out std_logic_vector(1 downto 0);
        IF_STALL, ID_STALL, EX_STALL, MEM_STALL, WB_STALL:   out std_logic -- stall signals
      );
  
  end component;
    
    component BHT is 
      generic (
        NBIT : integer := 32;   -- NUMBER OF BITS OF THE PROGRAM COUNTER
        N_ENTRIES : integer := 16;      -- Change this value to set the number of entries
        WORD_OFFSET : integer := 0    -- word offset bits, to be discarded by the internal memory
      );
    
      port (
        clock   : in std_logic;
        rst   : in std_logic;
        address : in std_logic_vector(NBIT - 1 downto 0);      -- address contained by the PC
        d_in    : in std_logic;                                 -- write 1 if the content of the memory should be incremented, 0 to decrement
        w_en    : in std_logic;                                 -- write enable
        d_out   : out std_logic                                 -- single bit to represent the prediction
      );
    end component;

    component FFD is
      Port (	D:	In	std_logic;
        CK:	In	std_logic;
        RESET:	In	std_logic;
        ENABLE : in std_logic;
        Q:	Out	std_logic);
    end component;
    
    component RF is
      generic(NBIT : integer := 32;
              NREG : integer := 32);
      port ( CLK: 		IN std_logic;
              RESET: 	IN std_logic;
        ENABLE: 	IN std_logic;
        RD1: 		IN std_logic;
        RD2: 		IN std_logic;
        WR: 		IN std_logic;
        ADD_WR: 	IN std_logic_vector(integer(log2(real(NREG)))-1 downto 0);
        ADD_RD1: 	IN std_logic_vector(integer(log2(real(NREG)))-1 downto 0);
        ADD_RD2: 	IN std_logic_vector(integer(log2(real(NREG)))-1 downto 0);
        DATAIN: 	IN std_logic_vector(NBIT - 1 downto 0);
              OUT1: 		OUT std_logic_vector(NBIT - 1 downto 0);
        OUT2: 		OUT std_logic_vector(NBIT - 1 downto 0));
     end component;


-- Initialization of signals to zero

signal IF_ENABLE: std_logic := '0';
signal IF_STALL: std_logic := '0';
signal PC_out: std_logic_vector(31 downto 0) := (others => '0');
signal IRAM_address: std_logic_vector(31 downto 0) := (others => '0');
signal IR_out: std_logic_vector(31 downto 0) := (others => '0');
signal NPC_in: std_logic_vector(31 downto 0) := (others => '0');
signal NPC_out: std_logic_vector(31 downto 0) := (others => '0');
signal PC_MUX_out: std_logic_vector(31 downto 0) := (others => '0');
signal STALL_CODE: std_logic_vector(1 downto 0):= "00";
signal FWDU_en : std_logic := '0';
signal jaddition : integer := 0;

-- Decode stage
signal ID_ENABLE: std_logic := '0';
signal ID_STALL: std_logic := '0';
signal PC_SEL: std_logic_vector(1 downto 0) := (others => '0');
signal PC2_out: std_logic_vector(31 downto 0) := (others => '0');
signal PC3_out: std_logic_vector(31 downto 0) := (others => '0');
signal IMM_out: std_logic_vector(31 downto 0) := (others => '0');
signal IMM_16: std_logic_vector(31 downto 0) := (others => '0');
signal IMM_26: std_logic_vector(31 downto 0) := (others => '0');
signal JADDER_out: std_logic_vector(31 downto 0) := (others => '0');
signal A_in: std_logic_vector(31 downto 0) := (others => '0');
signal B_in: std_logic_vector(31 downto 0) := (others => '0');
signal RA_out: std_logic_vector(31 downto 0) := (others => '0');
signal RB_out: std_logic_vector(31 downto 0) := (others => '0');
signal RIMM_in: std_logic_vector(31 downto 0) := (others => '0');
signal RIMM_out: std_logic_vector(31 downto 0) := (others => '0');
signal RWB1_out: std_logic_vector(31 downto 0) := (others => '0');
signal PRD_OUT: std_logic := '0';
signal BHT_in: std_logic_vector(31 downto 0) := (others => '0');
signal BHT_out: std_logic := '0';
signal NPC2_out: std_logic_vector(31 downto 0) := (others => '0');
signal ADDR_RA: std_logic_vector(4 downto 0) := (others => '0'); -- internal signal for Register File
signal ADDR_RB: std_logic_vector(4 downto 0) := (others => '0'); -- internal signal for Register File
signal IRAMMUX_SEL: std_logic;

-- Exe stage
signal EX_ENABLE: std_logic := '0';
signal EX_STALL: std_logic := '0';
signal FWDA_OUT: std_logic_vector(31 downto 0) := (others => '0');
signal FWDB_OUT: std_logic_vector(31 downto 0) := (others => '0');
signal ALR_in: std_logic_vector(31 downto 0) := (others => '0');
signal ALR_out: std_logic_vector(31 downto 0) := (others => '0');
signal JADDER2_out: std_logic_vector(31 downto 0) := (others => '0');
signal BPR_EN2: std_logic := '0';
signal FWDA_SEL: std_logic_vector(1 downto 0) := (others => '0');
signal FWDB_SEL: std_logic_vector(1 downto 0) := (others => '0');
signal PSW_in: std_logic_vector(6 downto 0) := (others => '0');
signal PSW_out: std_logic_vector(6 downto 0) := (others => '0');
signal NPC3_out: std_logic_vector(31 downto 0) := (others => '0');
signal RWB2_out: std_logic_vector(31 downto 0) := (others => '0');
signal CIN_masked: std_logic := '0';
signal CIN_ALU: std_logic := '0';
signal ALU_C_out: std_logic := '0';
signal ZDU_out: std_logic := '0';
signal BHT_update: std_logic := '0';
signal RF_RD_en : std_logic := '0';

-- Mem stage
signal MEM_ENABLE: std_logic := '0';
signal MEM_STALL: std_logic := '0';
signal ALR2_out: std_logic_vector(31 downto 0) := (others => '0');
signal LMD_out: std_logic_vector(31 downto 0) := (others => '0');
signal RWB3_out: std_logic_vector(31 downto 0) := (others => '0');
signal LW_CONF: std_logic_vector(31 downto 0) := (others => '0');
signal LB_CONF: std_logic_vector(31 downto 0) := (others => '0');
signal LBU_CONF: std_logic_vector(31 downto 0) := (others => '0');
signal LH_CONF: std_logic_vector(31 downto 0) := (others => '0');
signal LHU_CONF: std_logic_vector(31 downto 0) := (others => '0');
signal B2_out: std_logic_vector(31 downto 0) := (others => '0');
signal IMM_LHI: std_logic_vector(31 downto 0) := (others => '0');
signal CWB_out: std_logic_vector(1 downto 0) := (others => '0');
signal CWB2_SEL: std_logic_vector(1 downto 0) := (others => '0');
signal CWB_MUX_SEL: std_logic_vector(1 downto 0) := (others => '0');
signal CWB_MUX2_out: std_logic_vector(31 downto 0) := (others => '0');
signal ALR2_in: std_logic_vector(31 downto 0) := (others => '0');
signal ZDU_SEL: std_logic_vector(1 downto 0) := (others => '0');
signal ZDU_MUX_out: std_logic_vector(31 downto 0) := (others => '0');
signal FWDB2_SEL: std_logic:= '0';
signal B2_MUX_out: std_logic_vector(31 downto 0) := (others => '0');

-- WB stage
signal WB_STALL: std_logic := '0';
signal RF_MUX_out: std_logic_vector(4 downto 0) := (others => '0');
signal WB_in: std_logic_vector(31 downto 0) := (others => '0');
signal RF_WR_en: std_logic := '0';


begin

  IRAM_ADDR <= IRAM_address;

  -- REGISTERS DECLARATION

  -- FETCH STAGE
  RegPC: REG  
  generic map (32)
    port map (clk => CLK, reset => RST, enable => IF_ENABLE, data_in => NPC_in, data_out => PC_out);

  RegIR: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => IF_ENABLE, data_in => IRAM_OUT, data_out => IR_out);
  
  RegNPC: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => IF_ENABLE, data_in => NPC_in, data_out => NPC_out);
      

  -- DECODE STAGE
  
  RegPC2: REG  
  generic map (32)
    port map (clk => CLK, reset => RST, enable => ID_ENABLE, data_in => PC_out, data_out => PC2_out);

  
  RegIMM: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => ID_ENABLE, data_in => RIMM_in, data_out => RIMM_out);
    
  RegWB1: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => ID_ENABLE, data_in => IR_out, data_out => RWB1_out);
  

  F_PRD: FFD
      port map(CK => CLK, RESET => RST, ENABLE => ID_ENABLE, D => BHT_out, Q => PRD_out);

  RegNPC2: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => ID_ENABLE, data_in => NPC_out, data_out => NPC2_out);
  
  RegJADD2: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => ID_ENABLE, data_in => JADDER_out, data_out => JADDER2_out);
  

  F_JR: FFD
      port map(CK => CLK, RESET => RST, ENABLE => ID_ENABLE, D => BPR_EN, Q => BPR_EN2);


  RegPC3: REG  
  generic map (32)
    port map (clk => CLK, reset => RST, enable => EX_ENABLE, data_in => PC2_out, data_out => PC3_out);
  
  
  -- EXE STAGE
  RegWB2: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => EX_ENABLE, data_in => RWB1_out, data_out => RWB2_out);
  
  RegB2: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => EX_ENABLE, data_in => RB_out, data_out => B2_out);
  
  RegALR: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => EX_ENABLE, data_in => ALR_in, data_out => ALR_out);
 
  RegNPC3: REG  
    generic map (32)
      port map (clk => CLK, reset => RST, enable => EX_ENABLE, data_in => NPC2_out, data_out => NPC3_out);

  RegPSW: REG  
    generic map (7)
      port map (clk => CLK, reset => RST, enable => EX_ENABLE, data_in => PSW_in, data_out => PSW_out);


-- MEM STAGE
RegALR2: REG  
   generic map (32)
     port map (clk => CLK, reset => RST, enable => MEM_ENABLE, data_in => ALR2_in, data_out => ALR2_out);  

RegWB3: REG  
  generic map (32)
    port map (clk => CLK, reset => RST, enable =>MEM_ENABLE , data_in => RWB2_out, data_out => RWB3_out);
    
  --FETCH STAGE
  AdderPC: PC_adder port map(A => IRAM_address, B => "00000000000000000000000000000001", Sum => NPC_in);

  --DECODE STAGE 
  J_Adder: PC_adder port map(A => PC2_out, B => IMM_out, Sum => JADDER_out);
 


  -- MUXs DECLARATION
 
  --FETCH STAGE

  PCMUX: MUX3to1
    generic map (32)
    port map(A => PC_OUT, B => JADDER_out, C => JADDER2_out, SEL => PC_SEL , Y => PC_MUX_out);

  IRAMMUX: MUX2to1
    generic map (32)
    port map(A => PC_MUX_out, B => NPC2_out, SEL => IRAMMUX_SEL , Y => IRAM_address);
 
  --DECODE STAGE
  
  IMMMUX: MUX2to1
    generic map (32)
    port map(A => IMM_16 , B => IMM_26 , SEL => IMM_SEL , Y => IMM_out );

  BHTMUX: MUX2to1
    generic map (32)
    port map(A => PC2_out , B => PC3_out , SEL => BPR_EN2, Y => BHT_in);

  --EXE STAGE
  RegAMUX: MUX2to1 port map(A => FWDA_OUT, B=> (others =>'0'), SEL => ALUA_SEL, Y => A_in); 

  RegBMUX: MUX2to1 port map(A => FWDB_OUT, B=> RIMM_out, SEL => ALUB_SEL, Y => B_in);

  FWDA_MUX: MUX3to1
    generic map (32)
    port map(A => RA_out, B => ALR_out, C => WB_in, SEL => FWDA_SEL , Y => FWDA_OUT);

  FWDB_MUX: MUX3to1
    generic map (32)
    port map(A => RB_out, B => ALR_out, C => WB_in, SEL => FWDB_SEL , Y => FWDB_OUT);
  
  ZDU_MUX: MUX3to1 
    generic map (32)
    port map(A => RA_out, B => CWB_MUX2_out , C => WB_in, SEL => ZDU_SEL , Y => ZDU_MUX_out);
  
  --MEM STAGE
  MEMDATAMUX: MUX2to1
      generic map (32)
      port map( A => ALR2_out, B => B2_MUX_out, SEL => MEM_DATA_SEL, Y => DATA_OUT);

  LMDMUX: MUX5to1 
      generic map (32)
      port map(A => LW_CONF, B=> LB_CONF, C => LBU_CONF, D => LH_CONF, E => LHU_CONF, SEL => LD_SEL, Y => LMD_out);
  
  ALR2_MUX: MUX2to1
      generic map (32)
      port map(A => CWB_MUX2_out, B => NPC3_out, SEL => ALR2_SEL, Y => ALR2_in);

  CWB_MUX1: MUX3to1
      generic map (2)
      port map(A => "00", B => "11" ,C => CWB_out, SEL=> CWB_MUX_SEL, Y => CWB2_SEL);
  
  CWB_MUX2: MUX4to1 
      generic map (32)
      port map(A => ALR_out, B=> "00000000000000000000000000000001", C => "00000000000000000000000000000000", D => IMM_LHI, SEL => CWB2_SEL, Y => CWB_MUX2_out ); 

  B2_MUX: MUX2to1
      generic map (32)
      port map(A => B2_out, B => WB_in, SEL=> FWDB2_SEL, Y => B2_MUX_out);
  
      --WB STAGE
  WBMUX: MUX2to1
      generic map (32)
      port map(A => ALR2_out, B => LMD_out, SEL => WB_SEL, Y => WB_in);

  RF_MUX_ADDR: MUX3to1
      generic map (5)
      port map(A => RWB3_out(15 downto 11) , B => RWB3_out(20 downto 16), C=> "11111", SEL => RF_MUX_SEL, Y => RF_MUX_out);

  -- ALU DECLARATION

  ALU1: ALU port map (CLOCK => CLK, A => A_in, B => B_in, AluOpcode => ALU_OPCODE, Cin => CIN_ALU, COND => PSW_in(5 downto 0), ALU_out => ALR_in, Cout => PSW_in(6));

  -- FWD DECLARATION
  FWD1: FWDU port map (CLOCK => CLK, RESET => RST, EN => FWDU_en, IR => IR_out, FWD_A => FWDA_SEL, FWD_B => FWDB_SEL, FWD_B2 => FWDB2_SEL, ZDU_SEL => ZDU_SEL );

  --HDU DECLARATION
  HDU1: HDU generic map (32) port map (clk  => CLK, rst => RST, STALL_CODE => STALL_CODE, IR => IR_out, IF_STALL => IF_STALL, ID_STALL => ID_STALL , EX_STALL => EX_STALL , MEM_STALL => MEM_STALL, WB_STALL => WB_STALL);

  -- BHT DECLARATION
 BHT1: BHT 
 generic map(32,8,0)
 port map (clock => CLK, rst => RST, address => BHT_in, d_in => ZDU_out, w_en => BPR_EN2, d_out => BHT_out);

  -- CWBU DECLARATION
  CWBU1: CWBU port map (CLOCK => CLK, ALU_OP => ALU_OPCODE, PSW => PSW_out, COND_SEL => CWB_out, CWB_SEL => CWB_SEL, CWB_MUW_SEL => CWB_MUX_SEL); 

  -- RF declaration
  RF1: RF
  generic map(32,32) 
    port map (CLK => CLK, RESET => RST, ENABLE => '1', RD1 => RF_RD_en, RD2 => RF_RD_en, WR => RF_WR, ADD_WR => RF_MUX_out, ADD_RD1 => ADDR_RA,
  ADD_RD2 => ADDR_RB, DATAIN => WB_in, OUT1 => RA_out, OUT2 => RB_out);
  
  -- Datapath ports mapping with internal signals

  -- SIGN EXTENSION:
  RIMM_in <= "1111111111111111" & IR_out(15 downto 0) when (IR_out(15) and SIGND) = '1' else
             "0000000000000000" & IR_out(15 downto 0); 
  
  IMM_26 <= "111111" & IR_out(25 downto 0) when IR_out(25)='1' else "000000" & IR_out(25 downto 0) ;
  IMM_16   <= "1111111111111111" & IR_out(15 downto 0) when IR_out(15)='1' else "0000000000000000" & IR_out(15 downto 0) ;
  

  ADDR_RA <=IR_out(25 downto 21);
  ADDR_RB <= IR_out(20 downto 16);
  STALL <= STALL_CODE;
  DATA_ADDR <= ALR_out;


  --ENABLE SIGNALS
  IF_ENABLE <= not(IF_STALL);
  ID_ENABLE <= ID_EN and (not(ID_STALL));
  EX_ENABLE <= EX_EN and (not(EX_STALL));
  MEM_ENABLE <= MEM_EN and (not(MEM_STALL));
  RF_WR_en <= '0' when (RF_WR = '0' or WB_STALL = '1' or BHT_out = '1' or (BMP = '1' and PRD_out = '0')) else
              '1';
  RF_RD_en <= RF_RD and (not(ID_STALL)) ;
  FWDU_en <= not(ID_STALL);

  --LOAD CONFIGURATIONS
  LB_CONF <= "111111111111111111111111" & DATA_IN(7 downto 0) when DATA_IN(7) = '1' else
             "000000000000000000000000" & DATA_IN(7 downto 0);
  
  LBU_CONF <= "000000000000000000000000" & DATA_IN(7 downto 0);

  LH_CONF <= "1111111111111111" & DATA_IN(7 downto 0) & DATA_IN(15 downto 8) when DATA_IN(7) = '1' else
             "0000000000000000" & DATA_IN(7 downto 0) & DATA_IN(15 downto 8);

  LHU_CONF <= "0000000000000000" & DATA_IN(7 downto 0) & DATA_IN(15 downto 8);

  LW_CONF <= DATA_IN(7 downto 0) & DATA_IN(15 downto 8) & DATA_IN(23 downto 16) & DATA_IN(31 downto 24);

  --IMM LHI
  IMM_LHI <= ALR_out(15 downto 0) & "0000000000000000";     --USED FOR LHI instruction : ALR_OUT contains IMM16 + 0, SO MOVE IT TO MSB


  --PC_SEL = '1' when there is a J-INSTRUCTION (UCB_EN ='1') or when both BPR_EN and the output of BHT are = '1'
  PC_SEL <= "01" when ((BPR_EN = '1' and BHT_out = '1') or UCB_EN = '1') else
            "10" when (BMP = '1' and PRD_out = '0') else
            "00";
  
  --ZERO DETECTOR UNIT: DETECT IF THE 'A' REGISTER IS ZERO, FOR BRANCH INSTRUCTIONS, DEPENDING ON THE LSB OF THE OPCODE
  --BEQZ = 0x04   ==> LSB = 0
  --BNE = 0x05    ==> LSB = 1
  ZDU_out <= '1' when (to_integer(unsigned(ZDU_MUX_out)) = 0 and RWB1_out(26) = '0') 
          else '1' when (to_integer(unsigned(ZDU_MUX_out)) /= 0 and RWB1_out(26) = '1')
          else '0';

  --BMP is READY AT EX STAGE
  -- BMP = '1' when misprediction (BPR_EN = '1' and PRD_out \= ZDU_out)
  -- otherwise BMP = '0'
  BMP <= BPR_EN2 and (PRD_out xor ZDU_out);
  IRAMMUX_SEL <= BMP and PRD_OUT;

  --ADC OPERATION, ANDING THE CARRY IN WITH ADC SIGNAL FROM THE CONTROL UNIT

   CIN_ALU <= PSW_out(6);
 
end architecture BEHAVIORAL;