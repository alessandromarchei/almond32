
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_NOP, OP_ADD, OP_ADC, OP_AND, OP_SRA, OP_OR, OP_SEQ, OP_SNE, 
   OP_SLT, OP_SGT, OP_SLE, OP_SGE, OP_SLL, OP_SRL, OP_SUB, OP_XOR, OP_NOR, 
   OP_XNOR, OP_NAND, OP_MUL);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011";

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_60;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n21, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U4 : INV_X1 port map( A => n22, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n19, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_24;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n19, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_53;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_52;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_51;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_50;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_49;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_39;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n20, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_38;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n20, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_37;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_36;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_35;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_34;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_23;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n20, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_22;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n20, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_21;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_20;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_19;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_18;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n22, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U4 : INV_X1 port map( A => n19, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U6 : INV_X1 port map( A => n20, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U8 : INV_X1 port map( A => n21, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_32;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n21, ZN => Y(2));
   U2 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U3 : INV_X1 port map( A => n20, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U5 : INV_X1 port map( A => n19, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U7 : INV_X1 port map( A => SEL, ZN => n18);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_16;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n19, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U3 : INV_X1 port map( A => SEL, ZN => n18);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_46;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_45;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_42;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_31;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_30;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_29;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_28;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_26;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n19, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_15;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_14;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_13;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_12;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_41;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_25;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_9;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n19, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);
   U4 : INV_X1 port map( A => n20, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U6 : INV_X1 port map( A => n21, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U8 : INV_X1 port map( A => n22, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_5;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n22, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U8 : INV_X1 port map( A => n19, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_4;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n20, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n20);
   U4 : INV_X1 port map( A => n21, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n21);
   U6 : INV_X1 port map( A => n22, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n22);
   U8 : INV_X1 port map( A => n19, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_126 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_126;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_126 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_125 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_125;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_125 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_124 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_124;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_124 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_123 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_123;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_123 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_122 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_122;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_122 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_121 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_121;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_121 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_120 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_120;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_120 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_119 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_119;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_119 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_118 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_118;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_118 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_117 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_117;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_117 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_116 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_116;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_116 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_115 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_115;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_115 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_114 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_114;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_114 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_113 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_113;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_113 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_112 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_112;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_112 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_111 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_111;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_111 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_110 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_110;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_110 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_109 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_109;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_109 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_108 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_108;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_108 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_107 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_107;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_107 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_106 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_106;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_106 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_105 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_105;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_105 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_104 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_104;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_104 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_103 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_103;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_103 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_102 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_102;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_102 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_101 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_101;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_101 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_100 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_100;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_100 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_99 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_99;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_99 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_98 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_98;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_98 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_97 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_97;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_97 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_96 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_96;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_96 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_95 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_95;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_95 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_94 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_94;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_94 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_93 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_93;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_93 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_92 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_92;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_92 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_91 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_91;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_91 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_90 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_90;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_90 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_89 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_89;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_89 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_88 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_88;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_88 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_87 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_87;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_87 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_86 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_86;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_86 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_85 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_85;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_85 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_84 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_84;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_84 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_83 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_83;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_83 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_82 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_82;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_82 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_81 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_81;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_81 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_80 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_80;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_80 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_79 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_79;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_79 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_78 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_78;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_78 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_77 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_77;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_77 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_76 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_76;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_76 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_75 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_75;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_75 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_74 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_74;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_74 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_73 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_73;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_73 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_72 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_72;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_72 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_71 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_71;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_71 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_70 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_70;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_70 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_69 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_69;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_69 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_68 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_68;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_68 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_67 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_67;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_67 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_66 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_66;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_66 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_65 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_65;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_65 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_64 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_64;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_64 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_63;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_63 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_62;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_62 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_61;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_61 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_60;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_60 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_59;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_59 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_58;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_58 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_57;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_57 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_56;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_56 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_55;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_55 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_54;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_54 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_53;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_53 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_52;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_52 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_51;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_51 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_50;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_50 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_49;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_49 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_48;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_48 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_47;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_47 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_46;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_46 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_45;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_45 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_44;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_44 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_43;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_43 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_42;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_42 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_41;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_41 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_40;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_40 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_39;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_39 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_38;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_38 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_37;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_37 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_36;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_36 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_35;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_35 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_34;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_34 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_33;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_33 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_32;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_32 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_31;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_31 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_30;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_30 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_29;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_29 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_28;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_28 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_27;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_27 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_26;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_26 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_25;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_25 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_24;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_24 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_23;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_23 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_22;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_22 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_21;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_21 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_20;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_20 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_19;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_19 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_18;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_18 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_17;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_17 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_16;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_16 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_15;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_15 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_14;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_14 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_13;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_13 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_12;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_12 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_11;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_10;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_10 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_9;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_9 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_8;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_8 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_7;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_7 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_6;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_6 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_5;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_5 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_4;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_4 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_3;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_3 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_2;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_2 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_1;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_1 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_60;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_60 is

   component MUX2to1_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_119
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_120
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1000, n_1001 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_120 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1000);
   RCA0 : RCAN_NBIT4_119 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1001);
   MUX21 : MUX2to1_NBIT4_60 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_24;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_24 is

   component MUX2to1_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1002, n_1003 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1002);
   RCA0 : RCAN_NBIT4_47 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1003);
   MUX21 : MUX2to1_NBIT4_24 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_53;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_53 is

   component MUX2to1_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_105
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_106
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1004, n_1005 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_106 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1004);
   RCA0 : RCAN_NBIT4_105 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1005);
   MUX21 : MUX2to1_NBIT4_53 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_52;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_52 is

   component MUX2to1_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_103
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_104
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_104 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1006);
   RCA0 : RCAN_NBIT4_103 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1007);
   MUX21 : MUX2to1_NBIT4_52 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_51;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_51 is

   component MUX2to1_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_101
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_102
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_102 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1008);
   RCA0 : RCAN_NBIT4_101 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1009);
   MUX21 : MUX2to1_NBIT4_51 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_50;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_50 is

   component MUX2to1_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_99
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_100
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_100 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1010);
   RCA0 : RCAN_NBIT4_99 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1011);
   MUX21 : MUX2to1_NBIT4_50 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_49;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_49 is

   component MUX2to1_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_97
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_98
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_98 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1012);
   RCA0 : RCAN_NBIT4_97 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1013);
   MUX21 : MUX2to1_NBIT4_49 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_39;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_39 is

   component MUX2to1_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_77
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_78
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_78 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1014);
   RCA0 : RCAN_NBIT4_77 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1015);
   MUX21 : MUX2to1_NBIT4_39 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_38;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_38 is

   component MUX2to1_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_75
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_76
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1016, n_1017 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_76 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1016);
   RCA0 : RCAN_NBIT4_75 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1017);
   MUX21 : MUX2to1_NBIT4_38 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_37;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_37 is

   component MUX2to1_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_73
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_74
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1018, n_1019 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_74 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1018);
   RCA0 : RCAN_NBIT4_73 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1019);
   MUX21 : MUX2to1_NBIT4_37 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_36;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_36 is

   component MUX2to1_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_71
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_72
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1020, n_1021 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_72 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1020);
   RCA0 : RCAN_NBIT4_71 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1021);
   MUX21 : MUX2to1_NBIT4_36 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_35;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_35 is

   component MUX2to1_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_69
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_70
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1022, n_1023 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_70 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1022);
   RCA0 : RCAN_NBIT4_69 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1023);
   MUX21 : MUX2to1_NBIT4_35 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_34;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_34 is

   component MUX2to1_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_67
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_68
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1024, n_1025 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_68 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1024);
   RCA0 : RCAN_NBIT4_67 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1025);
   MUX21 : MUX2to1_NBIT4_34 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_23;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_23 is

   component MUX2to1_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1026, n_1027 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_46 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1026);
   RCA0 : RCAN_NBIT4_45 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1027);
   MUX21 : MUX2to1_NBIT4_23 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_22;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_22 is

   component MUX2to1_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1028, n_1029 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_44 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1028);
   RCA0 : RCAN_NBIT4_43 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1029);
   MUX21 : MUX2to1_NBIT4_22 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_21;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_21 is

   component MUX2to1_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1030, n_1031 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_42 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1030);
   RCA0 : RCAN_NBIT4_41 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1031);
   MUX21 : MUX2to1_NBIT4_21 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_20;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_20 is

   component MUX2to1_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1032, n_1033 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1032);
   RCA0 : RCAN_NBIT4_39 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1033);
   MUX21 : MUX2to1_NBIT4_20 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_19;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_19 is

   component MUX2to1_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1034, n_1035 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_38 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1034);
   RCA0 : RCAN_NBIT4_37 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1035);
   MUX21 : MUX2to1_NBIT4_19 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_18;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_18 is

   component MUX2to1_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1036, n_1037 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_36 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1036);
   RCA0 : RCAN_NBIT4_35 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1037);
   MUX21 : MUX2to1_NBIT4_18 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_32;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_32 is

   component MUX2to1_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_64
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1038, n_1039 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_64 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1038);
   RCA0 : RCAN_NBIT4_63 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1039);
   MUX21 : MUX2to1_NBIT4_32 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_16;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_16 is

   component MUX2to1_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1040, n_1041 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1040);
   RCA0 : RCAN_NBIT4_31 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1041);
   MUX21 : MUX2to1_NBIT4_16 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_46;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_46 is

   component MUX2to1_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_91
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_92
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1042, n_1043 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_92 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1042);
   RCA0 : RCAN_NBIT4_91 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1043);
   MUX21 : MUX2to1_NBIT4_46 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_45;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_45 is

   component MUX2to1_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_89
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_90
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1044, n_1045 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_90 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1044);
   RCA0 : RCAN_NBIT4_89 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1045);
   MUX21 : MUX2to1_NBIT4_45 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_42;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_42 is

   component MUX2to1_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_83
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_84
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1046, n_1047 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_84 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1046);
   RCA0 : RCAN_NBIT4_83 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1047);
   MUX21 : MUX2to1_NBIT4_42 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_31;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_31 is

   component MUX2to1_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1048, n_1049 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_62 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1048);
   RCA0 : RCAN_NBIT4_61 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1049);
   MUX21 : MUX2to1_NBIT4_31 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_30;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_30 is

   component MUX2to1_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1050, n_1051 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_60 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1050);
   RCA0 : RCAN_NBIT4_59 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1051);
   MUX21 : MUX2to1_NBIT4_30 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_29;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_29 is

   component MUX2to1_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1052, n_1053 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_58 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1052);
   RCA0 : RCAN_NBIT4_57 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1053);
   MUX21 : MUX2to1_NBIT4_29 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_28;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_28 is

   component MUX2to1_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1054, n_1055 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1054);
   RCA0 : RCAN_NBIT4_55 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1055);
   MUX21 : MUX2to1_NBIT4_28 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_26;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_26 is

   component MUX2to1_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1056, n_1057 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_52 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1056);
   RCA0 : RCAN_NBIT4_51 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1057);
   MUX21 : MUX2to1_NBIT4_26 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_15;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_15 is

   component MUX2to1_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1058, n_1059 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1058);
   RCA0 : RCAN_NBIT4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1059);
   MUX21 : MUX2to1_NBIT4_15 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_14;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_14 is

   component MUX2to1_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1060, n_1061 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1060);
   RCA0 : RCAN_NBIT4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1061);
   MUX21 : MUX2to1_NBIT4_14 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_13;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_13 is

   component MUX2to1_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1062, n_1063 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1062);
   RCA0 : RCAN_NBIT4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1063);
   MUX21 : MUX2to1_NBIT4_13 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_12;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_12 is

   component MUX2to1_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1064, n_1065 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1064);
   RCA0 : RCAN_NBIT4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1065);
   MUX21 : MUX2to1_NBIT4_12 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_41;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_41 is

   component MUX2to1_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_81
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_82
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1066, n_1067 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_82 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1066);
   RCA0 : RCAN_NBIT4_81 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1067);
   MUX21 : MUX2to1_NBIT4_41 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_25;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_25 is

   component MUX2to1_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1068, n_1069 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_50 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1068);
   RCA0 : RCAN_NBIT4_49 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1069);
   MUX21 : MUX2to1_NBIT4_25 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_9;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_9 is

   component MUX2to1_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1070, n_1071 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1070);
   RCA0 : RCAN_NBIT4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1071);
   MUX21 : MUX2to1_NBIT4_9 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_5;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_5 is

   component MUX2to1_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1072, n_1073 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1072);
   RCA0 : RCAN_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1073);
   MUX21 : MUX2to1_NBIT4_5 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_4;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_4 is

   component MUX2to1_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1074, n_1075 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1074);
   RCA0 : RCAN_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1075);
   MUX21 : MUX2to1_NBIT4_4 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_206 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_206;

architecture SYN_BEHAVIORAL of PG_block_206 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_174 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_174;

architecture SYN_BEHAVIORAL of PG_block_174 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_167 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_167;

architecture SYN_BEHAVIORAL of PG_block_167 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_164 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_164;

architecture SYN_BEHAVIORAL of PG_block_164 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_62 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_62;

architecture SYN_BEHAVIORAL of PG_block_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_18 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_18;

architecture SYN_BEHAVIORAL of PG_block_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_17 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_17;

architecture SYN_BEHAVIORAL of PG_block_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_213 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_213;

architecture SYN_BEHAVIORAL of PG_block_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_211 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_211;

architecture SYN_BEHAVIORAL of PG_block_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_209 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_209;

architecture SYN_BEHAVIORAL of PG_block_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_208 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_208;

architecture SYN_BEHAVIORAL of PG_block_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_207 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_207;

architecture SYN_BEHAVIORAL of PG_block_207 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_205 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_205;

architecture SYN_BEHAVIORAL of PG_block_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_204 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_204;

architecture SYN_BEHAVIORAL of PG_block_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_203 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_203;

architecture SYN_BEHAVIORAL of PG_block_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_202 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_202;

architecture SYN_BEHAVIORAL of PG_block_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_200 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_200;

architecture SYN_BEHAVIORAL of PG_block_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_199 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_199;

architecture SYN_BEHAVIORAL of PG_block_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_198 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_198;

architecture SYN_BEHAVIORAL of PG_block_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_197 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_197;

architecture SYN_BEHAVIORAL of PG_block_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_196 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_196;

architecture SYN_BEHAVIORAL of PG_block_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_195 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_195;

architecture SYN_BEHAVIORAL of PG_block_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_192 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_192;

architecture SYN_BEHAVIORAL of PG_block_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_189 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_189;

architecture SYN_BEHAVIORAL of PG_block_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_188 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_188;

architecture SYN_BEHAVIORAL of PG_block_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_187 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_187;

architecture SYN_BEHAVIORAL of PG_block_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_186 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_186;

architecture SYN_BEHAVIORAL of PG_block_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_185 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_185;

architecture SYN_BEHAVIORAL of PG_block_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_184 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_184;

architecture SYN_BEHAVIORAL of PG_block_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_182 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_182;

architecture SYN_BEHAVIORAL of PG_block_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_181 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_181;

architecture SYN_BEHAVIORAL of PG_block_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_178 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_178;

architecture SYN_BEHAVIORAL of PG_block_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_177 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_177;

architecture SYN_BEHAVIORAL of PG_block_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_173 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_173;

architecture SYN_BEHAVIORAL of PG_block_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_172 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_172;

architecture SYN_BEHAVIORAL of PG_block_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_171 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_171;

architecture SYN_BEHAVIORAL of PG_block_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_170 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_170;

architecture SYN_BEHAVIORAL of PG_block_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_169 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_169;

architecture SYN_BEHAVIORAL of PG_block_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_168 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_168;

architecture SYN_BEHAVIORAL of PG_block_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_166 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_166;

architecture SYN_BEHAVIORAL of PG_block_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_161 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_161;

architecture SYN_BEHAVIORAL of PG_block_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_160 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_160;

architecture SYN_BEHAVIORAL of PG_block_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_159 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_159;

architecture SYN_BEHAVIORAL of PG_block_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_158 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_158;

architecture SYN_BEHAVIORAL of PG_block_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_157 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_157;

architecture SYN_BEHAVIORAL of PG_block_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_156 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_156;

architecture SYN_BEHAVIORAL of PG_block_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_155 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_155;

architecture SYN_BEHAVIORAL of PG_block_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_154 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_154;

architecture SYN_BEHAVIORAL of PG_block_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_153 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_153;

architecture SYN_BEHAVIORAL of PG_block_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_152 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_152;

architecture SYN_BEHAVIORAL of PG_block_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_151 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_151;

architecture SYN_BEHAVIORAL of PG_block_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_150 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_150;

architecture SYN_BEHAVIORAL of PG_block_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_146 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_146;

architecture SYN_BEHAVIORAL of PG_block_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_145 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_145;

architecture SYN_BEHAVIORAL of PG_block_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_144 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_144;

architecture SYN_BEHAVIORAL of PG_block_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_143 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_143;

architecture SYN_BEHAVIORAL of PG_block_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_142 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_142;

architecture SYN_BEHAVIORAL of PG_block_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_141 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_141;

architecture SYN_BEHAVIORAL of PG_block_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_139 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_139;

architecture SYN_BEHAVIORAL of PG_block_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_134 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_134;

architecture SYN_BEHAVIORAL of PG_block_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_133 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_133;

architecture SYN_BEHAVIORAL of PG_block_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_132 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_132;

architecture SYN_BEHAVIORAL of PG_block_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_131 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_131;

architecture SYN_BEHAVIORAL of PG_block_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_130 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_130;

architecture SYN_BEHAVIORAL of PG_block_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_129 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_129;

architecture SYN_BEHAVIORAL of PG_block_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_128 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_128;

architecture SYN_BEHAVIORAL of PG_block_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_127 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_127;

architecture SYN_BEHAVIORAL of PG_block_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_126 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_126;

architecture SYN_BEHAVIORAL of PG_block_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_124 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_124;

architecture SYN_BEHAVIORAL of PG_block_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_123 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_123;

architecture SYN_BEHAVIORAL of PG_block_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_119 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_119;

architecture SYN_BEHAVIORAL of PG_block_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_118 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_118;

architecture SYN_BEHAVIORAL of PG_block_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_117 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_117;

architecture SYN_BEHAVIORAL of PG_block_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_116 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_116;

architecture SYN_BEHAVIORAL of PG_block_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_115 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_115;

architecture SYN_BEHAVIORAL of PG_block_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_114 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_114;

architecture SYN_BEHAVIORAL of PG_block_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_107 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_107;

architecture SYN_BEHAVIORAL of PG_block_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_106 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_106;

architecture SYN_BEHAVIORAL of PG_block_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_105 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_105;

architecture SYN_BEHAVIORAL of PG_block_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_104 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_104;

architecture SYN_BEHAVIORAL of PG_block_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_103 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_103;

architecture SYN_BEHAVIORAL of PG_block_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_102 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_102;

architecture SYN_BEHAVIORAL of PG_block_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_101 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_101;

architecture SYN_BEHAVIORAL of PG_block_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_100 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_100;

architecture SYN_BEHAVIORAL of PG_block_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_99 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_99;

architecture SYN_BEHAVIORAL of PG_block_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_98 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_98;

architecture SYN_BEHAVIORAL of PG_block_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_97 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_97;

architecture SYN_BEHAVIORAL of PG_block_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_96 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_96;

architecture SYN_BEHAVIORAL of PG_block_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_92 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_92;

architecture SYN_BEHAVIORAL of PG_block_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_91 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_91;

architecture SYN_BEHAVIORAL of PG_block_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_90 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_90;

architecture SYN_BEHAVIORAL of PG_block_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_89 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_89;

architecture SYN_BEHAVIORAL of PG_block_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_88 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_88;

architecture SYN_BEHAVIORAL of PG_block_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_87 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_87;

architecture SYN_BEHAVIORAL of PG_block_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_85 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_85;

architecture SYN_BEHAVIORAL of PG_block_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_80 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_80;

architecture SYN_BEHAVIORAL of PG_block_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_79 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_79;

architecture SYN_BEHAVIORAL of PG_block_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_78 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_78;

architecture SYN_BEHAVIORAL of PG_block_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_77 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_77;

architecture SYN_BEHAVIORAL of PG_block_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_76 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_76;

architecture SYN_BEHAVIORAL of PG_block_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_75 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_75;

architecture SYN_BEHAVIORAL of PG_block_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_74 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_74;

architecture SYN_BEHAVIORAL of PG_block_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_73 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_73;

architecture SYN_BEHAVIORAL of PG_block_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_70 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_70;

architecture SYN_BEHAVIORAL of PG_block_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_69 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_69;

architecture SYN_BEHAVIORAL of PG_block_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_65 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_65;

architecture SYN_BEHAVIORAL of PG_block_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_64 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_64;

architecture SYN_BEHAVIORAL of PG_block_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_63 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_63;

architecture SYN_BEHAVIORAL of PG_block_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_61 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_61;

architecture SYN_BEHAVIORAL of PG_block_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_60 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_60;

architecture SYN_BEHAVIORAL of PG_block_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_53 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_53;

architecture SYN_BEHAVIORAL of PG_block_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_52 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_52;

architecture SYN_BEHAVIORAL of PG_block_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_51 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_51;

architecture SYN_BEHAVIORAL of PG_block_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_50 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_50;

architecture SYN_BEHAVIORAL of PG_block_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_49 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_49;

architecture SYN_BEHAVIORAL of PG_block_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_48 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_48;

architecture SYN_BEHAVIORAL of PG_block_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_47 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_47;

architecture SYN_BEHAVIORAL of PG_block_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_46 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_46;

architecture SYN_BEHAVIORAL of PG_block_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_45 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_45;

architecture SYN_BEHAVIORAL of PG_block_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_44 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_44;

architecture SYN_BEHAVIORAL of PG_block_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_43 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_43;

architecture SYN_BEHAVIORAL of PG_block_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_42 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_42;

architecture SYN_BEHAVIORAL of PG_block_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_38 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_38;

architecture SYN_BEHAVIORAL of PG_block_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_37 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_37;

architecture SYN_BEHAVIORAL of PG_block_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_36 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_36;

architecture SYN_BEHAVIORAL of PG_block_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_35 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_35;

architecture SYN_BEHAVIORAL of PG_block_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_34 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_34;

architecture SYN_BEHAVIORAL of PG_block_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_33 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_33;

architecture SYN_BEHAVIORAL of PG_block_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_31 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_31;

architecture SYN_BEHAVIORAL of PG_block_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_26 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_26;

architecture SYN_BEHAVIORAL of PG_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_25 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_25;

architecture SYN_BEHAVIORAL of PG_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_24 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_24;

architecture SYN_BEHAVIORAL of PG_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_23 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_23;

architecture SYN_BEHAVIORAL of PG_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_22 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_22;

architecture SYN_BEHAVIORAL of PG_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_21 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_21;

architecture SYN_BEHAVIORAL of PG_block_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_20 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_20;

architecture SYN_BEHAVIORAL of PG_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_19 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_19;

architecture SYN_BEHAVIORAL of PG_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_16 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_16;

architecture SYN_BEHAVIORAL of PG_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_15 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_15;

architecture SYN_BEHAVIORAL of PG_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_11 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_11;

architecture SYN_BEHAVIORAL of PG_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_10 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_10;

architecture SYN_BEHAVIORAL of PG_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_9 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_9;

architecture SYN_BEHAVIORAL of PG_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_8 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_8;

architecture SYN_BEHAVIORAL of PG_block_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_7 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_7;

architecture SYN_BEHAVIORAL of PG_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_6 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_6;

architecture SYN_BEHAVIORAL of PG_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_112 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_112;

architecture SYN_BEHAVIORAL of PG_block_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_72 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_72;

architecture SYN_BEHAVIORAL of PG_block_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_58 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_58;

architecture SYN_BEHAVIORAL of PG_block_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_4 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_4;

architecture SYN_BEHAVIORAL of PG_block_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_194 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_194;

architecture SYN_BEHAVIORAL of PG_block_194 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_190 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_190;

architecture SYN_BEHAVIORAL of PG_block_190 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_183 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_183;

architecture SYN_BEHAVIORAL of PG_block_183 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_180 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_180;

architecture SYN_BEHAVIORAL of PG_block_180 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_179 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_179;

architecture SYN_BEHAVIORAL of PG_block_179 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_176 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_176;

architecture SYN_BEHAVIORAL of PG_block_176 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_175 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_175;

architecture SYN_BEHAVIORAL of PG_block_175 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_165 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_165;

architecture SYN_BEHAVIORAL of PG_block_165 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_162 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_162;

architecture SYN_BEHAVIORAL of PG_block_162 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_149 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_149;

architecture SYN_BEHAVIORAL of PG_block_149 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_148 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_148;

architecture SYN_BEHAVIORAL of PG_block_148 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_147 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_147;

architecture SYN_BEHAVIORAL of PG_block_147 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_140 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_140;

architecture SYN_BEHAVIORAL of PG_block_140 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_138 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_138;

architecture SYN_BEHAVIORAL of PG_block_138 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_137 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_137;

architecture SYN_BEHAVIORAL of PG_block_137 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_135 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_135;

architecture SYN_BEHAVIORAL of PG_block_135 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_122 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_122;

architecture SYN_BEHAVIORAL of PG_block_122 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_121 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_121;

architecture SYN_BEHAVIORAL of PG_block_121 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_120 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_120;

architecture SYN_BEHAVIORAL of PG_block_120 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_113 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_113;

architecture SYN_BEHAVIORAL of PG_block_113 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_111 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_111;

architecture SYN_BEHAVIORAL of PG_block_111 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_110 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_110;

architecture SYN_BEHAVIORAL of PG_block_110 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_108 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_108;

architecture SYN_BEHAVIORAL of PG_block_108 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_95 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_95;

architecture SYN_BEHAVIORAL of PG_block_95 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_94 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_94;

architecture SYN_BEHAVIORAL of PG_block_94 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_93 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_93;

architecture SYN_BEHAVIORAL of PG_block_93 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_86 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_86;

architecture SYN_BEHAVIORAL of PG_block_86 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_84 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_84;

architecture SYN_BEHAVIORAL of PG_block_84 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_83 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_83;

architecture SYN_BEHAVIORAL of PG_block_83 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_81 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_81;

architecture SYN_BEHAVIORAL of PG_block_81 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_71 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_71;

architecture SYN_BEHAVIORAL of PG_block_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_68 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_68;

architecture SYN_BEHAVIORAL of PG_block_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_67 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_67;

architecture SYN_BEHAVIORAL of PG_block_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_66 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_66;

architecture SYN_BEHAVIORAL of PG_block_66 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_59 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_59;

architecture SYN_BEHAVIORAL of PG_block_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_57 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_57;

architecture SYN_BEHAVIORAL of PG_block_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_56 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_56;

architecture SYN_BEHAVIORAL of PG_block_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_41 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_41;

architecture SYN_BEHAVIORAL of PG_block_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_40 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_40;

architecture SYN_BEHAVIORAL of PG_block_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_39 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_39;

architecture SYN_BEHAVIORAL of PG_block_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_32 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_32;

architecture SYN_BEHAVIORAL of PG_block_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_30 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_30;

architecture SYN_BEHAVIORAL of PG_block_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_29 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_29;

architecture SYN_BEHAVIORAL of PG_block_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_27 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_27;

architecture SYN_BEHAVIORAL of PG_block_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_14 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_14;

architecture SYN_BEHAVIORAL of PG_block_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_13 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_13;

architecture SYN_BEHAVIORAL of PG_block_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_12 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_12;

architecture SYN_BEHAVIORAL of PG_block_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_5 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_5;

architecture SYN_BEHAVIORAL of PG_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_3 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_3;

architecture SYN_BEHAVIORAL of PG_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_54 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_54;

architecture SYN_BEHAVIORAL of PG_block_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_2 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_2;

architecture SYN_BEHAVIORAL of PG_block_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_210 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_210;

architecture SYN_BEHAVIORAL of PG_block_210 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n5, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_163 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_163;

architecture SYN_BEHAVIORAL of PG_block_163 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_136 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_136;

architecture SYN_BEHAVIORAL of PG_block_136 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_109 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_109;

architecture SYN_BEHAVIORAL of PG_block_109 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_82 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_82;

architecture SYN_BEHAVIORAL of PG_block_82 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_55 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_55;

architecture SYN_BEHAVIORAL of PG_block_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_28 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_28;

architecture SYN_BEHAVIORAL of PG_block_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_1 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_1;

architecture SYN_BEHAVIORAL of PG_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_32 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_32;

architecture SYN_BEHAVIORAL of G_block_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_2 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_2;

architecture SYN_BEHAVIORAL of G_block_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_70 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_70;

architecture SYN_BEHAVIORAL of G_block_70 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_69 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_69;

architecture SYN_BEHAVIORAL of G_block_69 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_68 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_68;

architecture SYN_BEHAVIORAL of G_block_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_67 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_67;

architecture SYN_BEHAVIORAL of G_block_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_66 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_66;

architecture SYN_BEHAVIORAL of G_block_66 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_65 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_65;

architecture SYN_BEHAVIORAL of G_block_65 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_64 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_64;

architecture SYN_BEHAVIORAL of G_block_64 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_63 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_63;

architecture SYN_BEHAVIORAL of G_block_63 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_62 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_62;

architecture SYN_BEHAVIORAL of G_block_62 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_61 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_61;

architecture SYN_BEHAVIORAL of G_block_61 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_60 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_60;

architecture SYN_BEHAVIORAL of G_block_60 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_59 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_59;

architecture SYN_BEHAVIORAL of G_block_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_58 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_58;

architecture SYN_BEHAVIORAL of G_block_58 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_57 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_57;

architecture SYN_BEHAVIORAL of G_block_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_56 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_56;

architecture SYN_BEHAVIORAL of G_block_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_55 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_55;

architecture SYN_BEHAVIORAL of G_block_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_54 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_54;

architecture SYN_BEHAVIORAL of G_block_54 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_53 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_53;

architecture SYN_BEHAVIORAL of G_block_53 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_51 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_51;

architecture SYN_BEHAVIORAL of G_block_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_49 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_49;

architecture SYN_BEHAVIORAL of G_block_49 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_48 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_48;

architecture SYN_BEHAVIORAL of G_block_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_47 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_47;

architecture SYN_BEHAVIORAL of G_block_47 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_46 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_46;

architecture SYN_BEHAVIORAL of G_block_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_45 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_45;

architecture SYN_BEHAVIORAL of G_block_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_44 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_44;

architecture SYN_BEHAVIORAL of G_block_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_43 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_43;

architecture SYN_BEHAVIORAL of G_block_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_42 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_42;

architecture SYN_BEHAVIORAL of G_block_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_41 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_41;

architecture SYN_BEHAVIORAL of G_block_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_40 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_40;

architecture SYN_BEHAVIORAL of G_block_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_39 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_39;

architecture SYN_BEHAVIORAL of G_block_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_37 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_37;

architecture SYN_BEHAVIORAL of G_block_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_36 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_36;

architecture SYN_BEHAVIORAL of G_block_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_35 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_35;

architecture SYN_BEHAVIORAL of G_block_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_34 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_34;

architecture SYN_BEHAVIORAL of G_block_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_33 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_33;

architecture SYN_BEHAVIORAL of G_block_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_31 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_31;

architecture SYN_BEHAVIORAL of G_block_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_30 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_30;

architecture SYN_BEHAVIORAL of G_block_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_29 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_29;

architecture SYN_BEHAVIORAL of G_block_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_28 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_28;

architecture SYN_BEHAVIORAL of G_block_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_27 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_27;

architecture SYN_BEHAVIORAL of G_block_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_26 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_26;

architecture SYN_BEHAVIORAL of G_block_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_25 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_25;

architecture SYN_BEHAVIORAL of G_block_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_24 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_24;

architecture SYN_BEHAVIORAL of G_block_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_23 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_23;

architecture SYN_BEHAVIORAL of G_block_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_22 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_22;

architecture SYN_BEHAVIORAL of G_block_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_21 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_21;

architecture SYN_BEHAVIORAL of G_block_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_20 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_20;

architecture SYN_BEHAVIORAL of G_block_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_19 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_19;

architecture SYN_BEHAVIORAL of G_block_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_18 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_18;

architecture SYN_BEHAVIORAL of G_block_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_17 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_17;

architecture SYN_BEHAVIORAL of G_block_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_16 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_16;

architecture SYN_BEHAVIORAL of G_block_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_15 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_15;

architecture SYN_BEHAVIORAL of G_block_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_14 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_14;

architecture SYN_BEHAVIORAL of G_block_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_13 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_13;

architecture SYN_BEHAVIORAL of G_block_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_12 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_12;

architecture SYN_BEHAVIORAL of G_block_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_11 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_11;

architecture SYN_BEHAVIORAL of G_block_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_10 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_10;

architecture SYN_BEHAVIORAL of G_block_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_9 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_9;

architecture SYN_BEHAVIORAL of G_block_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_8 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_8;

architecture SYN_BEHAVIORAL of G_block_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_7 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_7;

architecture SYN_BEHAVIORAL of G_block_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_6 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_6;

architecture SYN_BEHAVIORAL of G_block_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_5 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_5;

architecture SYN_BEHAVIORAL of G_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_4 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_4;

architecture SYN_BEHAVIORAL of G_block_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_3 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_3;

architecture SYN_BEHAVIORAL of G_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_1 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_1;

architecture SYN_BEHAVIORAL of G_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_6 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_6;

architecture SYN_BEHAVIORAL of ENCODER_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n10, A2 => n9, B1 => INPUT(2), B2 => n11, ZN 
                           => OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n10, B2 => n11, A => INPUT(2), ZN => OUTPUT(0)
                           );
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n10);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n11, A3 => n10, ZN => OUTPUT(2)
                           );
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_5 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_5;

architecture SYN_BEHAVIORAL of ENCODER_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n10, A2 => n9, B1 => INPUT(2), B2 => n11, ZN 
                           => OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n10, B2 => n11, A => INPUT(2), ZN => OUTPUT(0)
                           );
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n10);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n11, A3 => n10, ZN => OUTPUT(2)
                           );
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_4 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_4;

architecture SYN_BEHAVIORAL of ENCODER_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n10, A2 => n9, B1 => INPUT(2), B2 => n11, ZN 
                           => OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n10, B2 => n11, A => INPUT(2), ZN => OUTPUT(0)
                           );
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n10);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n11, A3 => n10, ZN => OUTPUT(2)
                           );
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_3 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_3;

architecture SYN_BEHAVIORAL of ENCODER_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n10, A2 => n9, B1 => INPUT(2), B2 => n11, ZN 
                           => OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n10, B2 => n11, A => INPUT(2), ZN => OUTPUT(0)
                           );
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n10);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n11, A3 => n10, ZN => OUTPUT(2)
                           );
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_2 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_2;

architecture SYN_BEHAVIORAL of ENCODER_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n10, A2 => n9, B1 => INPUT(2), B2 => n11, ZN 
                           => OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n10, B2 => n11, A => INPUT(2), ZN => OUTPUT(0)
                           );
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n10);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n11, A3 => n10, ZN => OUTPUT(2)
                           );
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_1 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_1;

architecture SYN_BEHAVIORAL of ENCODER_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n10, A2 => n9, B1 => INPUT(2), B2 => n11, ZN 
                           => OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n10, B2 => n11, A => INPUT(2), ZN => OUTPUT(0)
                           );
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n10);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n11, A3 => n10, ZN => OUTPUT(2)
                           );
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_31 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_31;

architecture SYN_ARCH1 of ND4_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_30 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_30;

architecture SYN_ARCH1 of ND4_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_29 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_29;

architecture SYN_ARCH1 of ND4_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_28 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_28;

architecture SYN_ARCH1 of ND4_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_27 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_27;

architecture SYN_ARCH1 of ND4_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_26 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_26;

architecture SYN_ARCH1 of ND4_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_25 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_25;

architecture SYN_ARCH1 of ND4_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_24 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_24;

architecture SYN_ARCH1 of ND4_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_23 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_23;

architecture SYN_ARCH1 of ND4_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_22 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_22;

architecture SYN_ARCH1 of ND4_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_21 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_21;

architecture SYN_ARCH1 of ND4_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_20 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_20;

architecture SYN_ARCH1 of ND4_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_19 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_19;

architecture SYN_ARCH1 of ND4_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_18 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_18;

architecture SYN_ARCH1 of ND4_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_17 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_17;

architecture SYN_ARCH1 of ND4_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_16 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_16;

architecture SYN_ARCH1 of ND4_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_15 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_15;

architecture SYN_ARCH1 of ND4_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_14 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_14;

architecture SYN_ARCH1 of ND4_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_13 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_13;

architecture SYN_ARCH1 of ND4_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_12 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_12;

architecture SYN_ARCH1 of ND4_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_11 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_11;

architecture SYN_ARCH1 of ND4_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_10 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_10;

architecture SYN_ARCH1 of ND4_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_9 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_9;

architecture SYN_ARCH1 of ND4_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_8 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_8;

architecture SYN_ARCH1 of ND4_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_7 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_7;

architecture SYN_ARCH1 of ND4_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_6 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_6;

architecture SYN_ARCH1 of ND4_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_5 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_5;

architecture SYN_ARCH1 of ND4_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_4 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_4;

architecture SYN_ARCH1 of ND4_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_3 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_3;

architecture SYN_ARCH1 of ND4_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_2 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_2;

architecture SYN_ARCH1 of ND4_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_1 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_1;

architecture SYN_ARCH1 of ND4_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_127 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_127;

architecture SYN_ARCH1 of ND3_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_126 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_126;

architecture SYN_ARCH1 of ND3_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_125 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_125;

architecture SYN_ARCH1 of ND3_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_124 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_124;

architecture SYN_ARCH1 of ND3_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_123 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_123;

architecture SYN_ARCH1 of ND3_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_122 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_122;

architecture SYN_ARCH1 of ND3_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_121 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_121;

architecture SYN_ARCH1 of ND3_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_120 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_120;

architecture SYN_ARCH1 of ND3_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_119 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_119;

architecture SYN_ARCH1 of ND3_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_118 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_118;

architecture SYN_ARCH1 of ND3_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_117 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_117;

architecture SYN_ARCH1 of ND3_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_116 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_116;

architecture SYN_ARCH1 of ND3_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_115 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_115;

architecture SYN_ARCH1 of ND3_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_114 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_114;

architecture SYN_ARCH1 of ND3_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_113 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_113;

architecture SYN_ARCH1 of ND3_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_112 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_112;

architecture SYN_ARCH1 of ND3_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_111 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_111;

architecture SYN_ARCH1 of ND3_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_110 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_110;

architecture SYN_ARCH1 of ND3_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_109 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_109;

architecture SYN_ARCH1 of ND3_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_108 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_108;

architecture SYN_ARCH1 of ND3_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_107 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_107;

architecture SYN_ARCH1 of ND3_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_106 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_106;

architecture SYN_ARCH1 of ND3_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_105 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_105;

architecture SYN_ARCH1 of ND3_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_104 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_104;

architecture SYN_ARCH1 of ND3_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_103 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_103;

architecture SYN_ARCH1 of ND3_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_102 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_102;

architecture SYN_ARCH1 of ND3_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_101 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_101;

architecture SYN_ARCH1 of ND3_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_100 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_100;

architecture SYN_ARCH1 of ND3_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_99 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_99;

architecture SYN_ARCH1 of ND3_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_98 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_98;

architecture SYN_ARCH1 of ND3_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_97 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_97;

architecture SYN_ARCH1 of ND3_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_96 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_96;

architecture SYN_ARCH1 of ND3_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_95 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_95;

architecture SYN_ARCH1 of ND3_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_94 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_94;

architecture SYN_ARCH1 of ND3_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_93 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_93;

architecture SYN_ARCH1 of ND3_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_92 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_92;

architecture SYN_ARCH1 of ND3_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_91 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_91;

architecture SYN_ARCH1 of ND3_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_90 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_90;

architecture SYN_ARCH1 of ND3_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_89 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_89;

architecture SYN_ARCH1 of ND3_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_88 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_88;

architecture SYN_ARCH1 of ND3_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_87 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_87;

architecture SYN_ARCH1 of ND3_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_86 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_86;

architecture SYN_ARCH1 of ND3_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_85 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_85;

architecture SYN_ARCH1 of ND3_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_84 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_84;

architecture SYN_ARCH1 of ND3_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_83 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_83;

architecture SYN_ARCH1 of ND3_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_82 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_82;

architecture SYN_ARCH1 of ND3_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_81 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_81;

architecture SYN_ARCH1 of ND3_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_80 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_80;

architecture SYN_ARCH1 of ND3_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_79 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_79;

architecture SYN_ARCH1 of ND3_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_78 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_78;

architecture SYN_ARCH1 of ND3_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_77 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_77;

architecture SYN_ARCH1 of ND3_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_76 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_76;

architecture SYN_ARCH1 of ND3_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_75 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_75;

architecture SYN_ARCH1 of ND3_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_74 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_74;

architecture SYN_ARCH1 of ND3_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_73 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_73;

architecture SYN_ARCH1 of ND3_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_72 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_72;

architecture SYN_ARCH1 of ND3_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_71 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_71;

architecture SYN_ARCH1 of ND3_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_70 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_70;

architecture SYN_ARCH1 of ND3_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_69 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_69;

architecture SYN_ARCH1 of ND3_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_68 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_68;

architecture SYN_ARCH1 of ND3_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_67 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_67;

architecture SYN_ARCH1 of ND3_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_66 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_66;

architecture SYN_ARCH1 of ND3_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_65 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_65;

architecture SYN_ARCH1 of ND3_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_64 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_64;

architecture SYN_ARCH1 of ND3_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_63 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_63;

architecture SYN_ARCH1 of ND3_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_62 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_62;

architecture SYN_ARCH1 of ND3_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_61 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_61;

architecture SYN_ARCH1 of ND3_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_60 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_60;

architecture SYN_ARCH1 of ND3_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_59 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_59;

architecture SYN_ARCH1 of ND3_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_58 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_58;

architecture SYN_ARCH1 of ND3_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_57 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_57;

architecture SYN_ARCH1 of ND3_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_56 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_56;

architecture SYN_ARCH1 of ND3_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_55 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_55;

architecture SYN_ARCH1 of ND3_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_54 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_54;

architecture SYN_ARCH1 of ND3_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_53 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_53;

architecture SYN_ARCH1 of ND3_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_52 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_52;

architecture SYN_ARCH1 of ND3_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_51 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_51;

architecture SYN_ARCH1 of ND3_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_50 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_50;

architecture SYN_ARCH1 of ND3_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_49 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_49;

architecture SYN_ARCH1 of ND3_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_48 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_48;

architecture SYN_ARCH1 of ND3_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_47 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_47;

architecture SYN_ARCH1 of ND3_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_46 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_46;

architecture SYN_ARCH1 of ND3_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_45 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_45;

architecture SYN_ARCH1 of ND3_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_44 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_44;

architecture SYN_ARCH1 of ND3_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_43 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_43;

architecture SYN_ARCH1 of ND3_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_42 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_42;

architecture SYN_ARCH1 of ND3_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_41 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_41;

architecture SYN_ARCH1 of ND3_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_40 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_40;

architecture SYN_ARCH1 of ND3_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_39 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_39;

architecture SYN_ARCH1 of ND3_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_38 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_38;

architecture SYN_ARCH1 of ND3_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_37 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_37;

architecture SYN_ARCH1 of ND3_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_36 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_36;

architecture SYN_ARCH1 of ND3_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_35 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_35;

architecture SYN_ARCH1 of ND3_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_34 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_34;

architecture SYN_ARCH1 of ND3_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_33 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_33;

architecture SYN_ARCH1 of ND3_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_32 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_32;

architecture SYN_ARCH1 of ND3_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_31 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_31;

architecture SYN_ARCH1 of ND3_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_30 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_30;

architecture SYN_ARCH1 of ND3_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_29 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_29;

architecture SYN_ARCH1 of ND3_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_28 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_28;

architecture SYN_ARCH1 of ND3_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_27 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_27;

architecture SYN_ARCH1 of ND3_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_26 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_26;

architecture SYN_ARCH1 of ND3_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_25 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_25;

architecture SYN_ARCH1 of ND3_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_24 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_24;

architecture SYN_ARCH1 of ND3_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_23 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_23;

architecture SYN_ARCH1 of ND3_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_22 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_22;

architecture SYN_ARCH1 of ND3_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_21 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_21;

architecture SYN_ARCH1 of ND3_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_20 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_20;

architecture SYN_ARCH1 of ND3_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_19 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_19;

architecture SYN_ARCH1 of ND3_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_18 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_18;

architecture SYN_ARCH1 of ND3_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_17 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_17;

architecture SYN_ARCH1 of ND3_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_16 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_16;

architecture SYN_ARCH1 of ND3_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_15 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_15;

architecture SYN_ARCH1 of ND3_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_14 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_14;

architecture SYN_ARCH1 of ND3_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_13 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_13;

architecture SYN_ARCH1 of ND3_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_12 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_12;

architecture SYN_ARCH1 of ND3_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_11 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_11;

architecture SYN_ARCH1 of ND3_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_10 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_10;

architecture SYN_ARCH1 of ND3_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_9 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_9;

architecture SYN_ARCH1 of ND3_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_8 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_8;

architecture SYN_ARCH1 of ND3_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_7 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_7;

architecture SYN_ARCH1 of ND3_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_6 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_6;

architecture SYN_ARCH1 of ND3_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_5 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_5;

architecture SYN_ARCH1 of ND3_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_4 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_4;

architecture SYN_ARCH1 of ND3_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_3 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_3;

architecture SYN_ARCH1 of ND3_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_2 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_2;

architecture SYN_ARCH1 of ND3_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_1 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_1;

architecture SYN_ARCH1 of ND3_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_228;

architecture SYN_Behavioral of AND2_228 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_227;

architecture SYN_Behavioral of AND2_227 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_226;

architecture SYN_Behavioral of AND2_226 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_225;

architecture SYN_Behavioral of AND2_225 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_224;

architecture SYN_Behavioral of AND2_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_223;

architecture SYN_Behavioral of AND2_223 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_222;

architecture SYN_Behavioral of AND2_222 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_221;

architecture SYN_Behavioral of AND2_221 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_220;

architecture SYN_Behavioral of AND2_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_219;

architecture SYN_Behavioral of AND2_219 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_218;

architecture SYN_Behavioral of AND2_218 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_217;

architecture SYN_Behavioral of AND2_217 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_216;

architecture SYN_Behavioral of AND2_216 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_215;

architecture SYN_Behavioral of AND2_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_214;

architecture SYN_Behavioral of AND2_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_213;

architecture SYN_Behavioral of AND2_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_212;

architecture SYN_Behavioral of AND2_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_211;

architecture SYN_Behavioral of AND2_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_210;

architecture SYN_Behavioral of AND2_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_209;

architecture SYN_Behavioral of AND2_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_208;

architecture SYN_Behavioral of AND2_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_207;

architecture SYN_Behavioral of AND2_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_206;

architecture SYN_Behavioral of AND2_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_205;

architecture SYN_Behavioral of AND2_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_204;

architecture SYN_Behavioral of AND2_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_203;

architecture SYN_Behavioral of AND2_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_202;

architecture SYN_Behavioral of AND2_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_201;

architecture SYN_Behavioral of AND2_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_200;

architecture SYN_Behavioral of AND2_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_199;

architecture SYN_Behavioral of AND2_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_198;

architecture SYN_Behavioral of AND2_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_197;

architecture SYN_Behavioral of AND2_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_196;

architecture SYN_Behavioral of AND2_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_195;

architecture SYN_Behavioral of AND2_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_194;

architecture SYN_Behavioral of AND2_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_193;

architecture SYN_Behavioral of AND2_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_192;

architecture SYN_Behavioral of AND2_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_191;

architecture SYN_Behavioral of AND2_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_190;

architecture SYN_Behavioral of AND2_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_189;

architecture SYN_Behavioral of AND2_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_188;

architecture SYN_Behavioral of AND2_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_187;

architecture SYN_Behavioral of AND2_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_186;

architecture SYN_Behavioral of AND2_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_185;

architecture SYN_Behavioral of AND2_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_184;

architecture SYN_Behavioral of AND2_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_183;

architecture SYN_Behavioral of AND2_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_182;

architecture SYN_Behavioral of AND2_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_181;

architecture SYN_Behavioral of AND2_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_180;

architecture SYN_Behavioral of AND2_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_179;

architecture SYN_Behavioral of AND2_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_178;

architecture SYN_Behavioral of AND2_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_177;

architecture SYN_Behavioral of AND2_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_176;

architecture SYN_Behavioral of AND2_176 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_175;

architecture SYN_Behavioral of AND2_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_174;

architecture SYN_Behavioral of AND2_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_173;

architecture SYN_Behavioral of AND2_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_172;

architecture SYN_Behavioral of AND2_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_171;

architecture SYN_Behavioral of AND2_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_170;

architecture SYN_Behavioral of AND2_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_169;

architecture SYN_Behavioral of AND2_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_168;

architecture SYN_Behavioral of AND2_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_167;

architecture SYN_Behavioral of AND2_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_166;

architecture SYN_Behavioral of AND2_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_165;

architecture SYN_Behavioral of AND2_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_164;

architecture SYN_Behavioral of AND2_164 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_163;

architecture SYN_Behavioral of AND2_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_162;

architecture SYN_Behavioral of AND2_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_161;

architecture SYN_Behavioral of AND2_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_160;

architecture SYN_Behavioral of AND2_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_159;

architecture SYN_Behavioral of AND2_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_158;

architecture SYN_Behavioral of AND2_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_157;

architecture SYN_Behavioral of AND2_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_156;

architecture SYN_Behavioral of AND2_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_155;

architecture SYN_Behavioral of AND2_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_154;

architecture SYN_Behavioral of AND2_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_153;

architecture SYN_Behavioral of AND2_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_152;

architecture SYN_Behavioral of AND2_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_151;

architecture SYN_Behavioral of AND2_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_150;

architecture SYN_Behavioral of AND2_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_149;

architecture SYN_Behavioral of AND2_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_148;

architecture SYN_Behavioral of AND2_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_147;

architecture SYN_Behavioral of AND2_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_146;

architecture SYN_Behavioral of AND2_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_145;

architecture SYN_Behavioral of AND2_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_144;

architecture SYN_Behavioral of AND2_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_143;

architecture SYN_Behavioral of AND2_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_142;

architecture SYN_Behavioral of AND2_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_141;

architecture SYN_Behavioral of AND2_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_140;

architecture SYN_Behavioral of AND2_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_139;

architecture SYN_Behavioral of AND2_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_138;

architecture SYN_Behavioral of AND2_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_137;

architecture SYN_Behavioral of AND2_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_136;

architecture SYN_Behavioral of AND2_136 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_135;

architecture SYN_Behavioral of AND2_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_134;

architecture SYN_Behavioral of AND2_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_133;

architecture SYN_Behavioral of AND2_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_132;

architecture SYN_Behavioral of AND2_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_131;

architecture SYN_Behavioral of AND2_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_130;

architecture SYN_Behavioral of AND2_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_129;

architecture SYN_Behavioral of AND2_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_128;

architecture SYN_Behavioral of AND2_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_127;

architecture SYN_Behavioral of AND2_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_126;

architecture SYN_Behavioral of AND2_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_125;

architecture SYN_Behavioral of AND2_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_124;

architecture SYN_Behavioral of AND2_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_123;

architecture SYN_Behavioral of AND2_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_122;

architecture SYN_Behavioral of AND2_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_121;

architecture SYN_Behavioral of AND2_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_120;

architecture SYN_Behavioral of AND2_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_119;

architecture SYN_Behavioral of AND2_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_118;

architecture SYN_Behavioral of AND2_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_117;

architecture SYN_Behavioral of AND2_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_116;

architecture SYN_Behavioral of AND2_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_115;

architecture SYN_Behavioral of AND2_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_114;

architecture SYN_Behavioral of AND2_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_113;

architecture SYN_Behavioral of AND2_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_112;

architecture SYN_Behavioral of AND2_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_111;

architecture SYN_Behavioral of AND2_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_110;

architecture SYN_Behavioral of AND2_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_109;

architecture SYN_Behavioral of AND2_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_108;

architecture SYN_Behavioral of AND2_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_107;

architecture SYN_Behavioral of AND2_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_106;

architecture SYN_Behavioral of AND2_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_105;

architecture SYN_Behavioral of AND2_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_104;

architecture SYN_Behavioral of AND2_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_103;

architecture SYN_Behavioral of AND2_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_102;

architecture SYN_Behavioral of AND2_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_101;

architecture SYN_Behavioral of AND2_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_100;

architecture SYN_Behavioral of AND2_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_99;

architecture SYN_Behavioral of AND2_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_98;

architecture SYN_Behavioral of AND2_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_97;

architecture SYN_Behavioral of AND2_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_96;

architecture SYN_Behavioral of AND2_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_95;

architecture SYN_Behavioral of AND2_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_94;

architecture SYN_Behavioral of AND2_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_93;

architecture SYN_Behavioral of AND2_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_92;

architecture SYN_Behavioral of AND2_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_91;

architecture SYN_Behavioral of AND2_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_90;

architecture SYN_Behavioral of AND2_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_89;

architecture SYN_Behavioral of AND2_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_88;

architecture SYN_Behavioral of AND2_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_87;

architecture SYN_Behavioral of AND2_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_86;

architecture SYN_Behavioral of AND2_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_85;

architecture SYN_Behavioral of AND2_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_84;

architecture SYN_Behavioral of AND2_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_83;

architecture SYN_Behavioral of AND2_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_82;

architecture SYN_Behavioral of AND2_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_81;

architecture SYN_Behavioral of AND2_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_80;

architecture SYN_Behavioral of AND2_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_79;

architecture SYN_Behavioral of AND2_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_78;

architecture SYN_Behavioral of AND2_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_77;

architecture SYN_Behavioral of AND2_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_76;

architecture SYN_Behavioral of AND2_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_75;

architecture SYN_Behavioral of AND2_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_74;

architecture SYN_Behavioral of AND2_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_73;

architecture SYN_Behavioral of AND2_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_72;

architecture SYN_Behavioral of AND2_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_71;

architecture SYN_Behavioral of AND2_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_70;

architecture SYN_Behavioral of AND2_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_69;

architecture SYN_Behavioral of AND2_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_68;

architecture SYN_Behavioral of AND2_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_67;

architecture SYN_Behavioral of AND2_67 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_66;

architecture SYN_Behavioral of AND2_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_65;

architecture SYN_Behavioral of AND2_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_64;

architecture SYN_Behavioral of AND2_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_63;

architecture SYN_Behavioral of AND2_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_62;

architecture SYN_Behavioral of AND2_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_61;

architecture SYN_Behavioral of AND2_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_60;

architecture SYN_Behavioral of AND2_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_59;

architecture SYN_Behavioral of AND2_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_58;

architecture SYN_Behavioral of AND2_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_57;

architecture SYN_Behavioral of AND2_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_56;

architecture SYN_Behavioral of AND2_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_55;

architecture SYN_Behavioral of AND2_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_54;

architecture SYN_Behavioral of AND2_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_53;

architecture SYN_Behavioral of AND2_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_52;

architecture SYN_Behavioral of AND2_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_51;

architecture SYN_Behavioral of AND2_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_50;

architecture SYN_Behavioral of AND2_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_49;

architecture SYN_Behavioral of AND2_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_48;

architecture SYN_Behavioral of AND2_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_47;

architecture SYN_Behavioral of AND2_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_46;

architecture SYN_Behavioral of AND2_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_45;

architecture SYN_Behavioral of AND2_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_44;

architecture SYN_Behavioral of AND2_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_43;

architecture SYN_Behavioral of AND2_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_42;

architecture SYN_Behavioral of AND2_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_40;

architecture SYN_Behavioral of AND2_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_39;

architecture SYN_Behavioral of AND2_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_38;

architecture SYN_Behavioral of AND2_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_37;

architecture SYN_Behavioral of AND2_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_36;

architecture SYN_Behavioral of AND2_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_35;

architecture SYN_Behavioral of AND2_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_34;

architecture SYN_Behavioral of AND2_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_33;

architecture SYN_Behavioral of AND2_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_32;

architecture SYN_Behavioral of AND2_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_31;

architecture SYN_Behavioral of AND2_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_30;

architecture SYN_Behavioral of AND2_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_29;

architecture SYN_Behavioral of AND2_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_28;

architecture SYN_Behavioral of AND2_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_27;

architecture SYN_Behavioral of AND2_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_26;

architecture SYN_Behavioral of AND2_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_25;

architecture SYN_Behavioral of AND2_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_24;

architecture SYN_Behavioral of AND2_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_23;

architecture SYN_Behavioral of AND2_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_22;

architecture SYN_Behavioral of AND2_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_21;

architecture SYN_Behavioral of AND2_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_20;

architecture SYN_Behavioral of AND2_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_19;

architecture SYN_Behavioral of AND2_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_18;

architecture SYN_Behavioral of AND2_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_17;

architecture SYN_Behavioral of AND2_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_16;

architecture SYN_Behavioral of AND2_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_15;

architecture SYN_Behavioral of AND2_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_14;

architecture SYN_Behavioral of AND2_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_13;

architecture SYN_Behavioral of AND2_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_12;

architecture SYN_Behavioral of AND2_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_11;

architecture SYN_Behavioral of AND2_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_10;

architecture SYN_Behavioral of AND2_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_9;

architecture SYN_Behavioral of AND2_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_8;

architecture SYN_Behavioral of AND2_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_7;

architecture SYN_Behavioral of AND2_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_6;

architecture SYN_Behavioral of AND2_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_5;

architecture SYN_Behavioral of AND2_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_4;

architecture SYN_Behavioral of AND2_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_3;

architecture SYN_Behavioral of AND2_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_2;

architecture SYN_Behavioral of AND2_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_1;

architecture SYN_Behavioral of AND2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_2;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n105, n106, n107, n108, n109, n110, n111, n112, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n108, Z => n111);
   U2 : BUF_X1 port map( A => n108, Z => n112);
   U3 : BUF_X1 port map( A => n112, Z => n105);
   U4 : BUF_X1 port map( A => n112, Z => n106);
   U5 : INV_X1 port map( A => n111, ZN => n109);
   U6 : INV_X1 port map( A => n111, ZN => n110);
   U7 : BUF_X1 port map( A => n112, Z => n107);
   U8 : BUF_X1 port map( A => SEL, Z => n108);
   U9 : INV_X1 port map( A => n145, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n109, B1 => B(0), B2 => n105, ZN 
                           => n145);
   U11 : INV_X1 port map( A => n146, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n109, B1 => B(1), B2 => n105, ZN 
                           => n146);
   U13 : INV_X1 port map( A => n147, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => n109, B1 => B(2), B2 => n105, ZN 
                           => n147);
   U15 : INV_X1 port map( A => n148, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n109, B1 => B(3), B2 => n105, ZN 
                           => n148);
   U17 : INV_X1 port map( A => n149, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n109, B1 => B(4), B2 => n105, ZN 
                           => n149);
   U19 : INV_X1 port map( A => n150, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n109, B1 => B(5), B2 => n105, ZN 
                           => n150);
   U21 : INV_X1 port map( A => n151, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n109, B1 => B(6), B2 => n105, ZN 
                           => n151);
   U23 : INV_X1 port map( A => n152, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n109, B1 => B(7), B2 => n105, ZN 
                           => n152);
   U25 : INV_X1 port map( A => n153, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n109, B1 => B(8), B2 => n105, ZN 
                           => n153);
   U27 : INV_X1 port map( A => n154, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n109, B1 => B(9), B2 => n105, ZN 
                           => n154);
   U29 : INV_X1 port map( A => n155, ZN => Y(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n109, B1 => B(10), B2 => n105, 
                           ZN => n155);
   U31 : INV_X1 port map( A => n156, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => A(11), A2 => n109, B1 => B(11), B2 => n105, 
                           ZN => n156);
   U33 : INV_X1 port map( A => n157, ZN => Y(12));
   U34 : AOI22_X1 port map( A1 => A(12), A2 => n110, B1 => B(12), B2 => n106, 
                           ZN => n157);
   U35 : INV_X1 port map( A => n158, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n110, B1 => B(13), B2 => n106, 
                           ZN => n158);
   U37 : INV_X1 port map( A => n159, ZN => Y(14));
   U38 : AOI22_X1 port map( A1 => A(14), A2 => n110, B1 => B(14), B2 => n106, 
                           ZN => n159);
   U39 : INV_X1 port map( A => n160, ZN => Y(15));
   U40 : AOI22_X1 port map( A1 => A(15), A2 => n110, B1 => B(15), B2 => n106, 
                           ZN => n160);
   U41 : INV_X1 port map( A => n161, ZN => Y(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n110, B1 => B(16), B2 => n106, 
                           ZN => n161);
   U43 : INV_X1 port map( A => n162, ZN => Y(17));
   U44 : AOI22_X1 port map( A1 => A(17), A2 => n110, B1 => B(17), B2 => n106, 
                           ZN => n162);
   U45 : INV_X1 port map( A => n163, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n110, B1 => B(18), B2 => n106, 
                           ZN => n163);
   U47 : INV_X1 port map( A => n164, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n110, B1 => B(19), B2 => n106, 
                           ZN => n164);
   U49 : INV_X1 port map( A => n165, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n110, B1 => B(20), B2 => n106, 
                           ZN => n165);
   U51 : INV_X1 port map( A => n166, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n110, B1 => B(21), B2 => n106, 
                           ZN => n166);
   U53 : INV_X1 port map( A => n167, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n110, B1 => B(22), B2 => n106, 
                           ZN => n167);
   U55 : INV_X1 port map( A => n168, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n110, B1 => B(23), B2 => n106, 
                           ZN => n168);
   U57 : INV_X1 port map( A => n169, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A(24), A2 => n109, B1 => B(24), B2 => n107, 
                           ZN => n169);
   U59 : INV_X1 port map( A => n170, ZN => Y(25));
   U60 : AOI22_X1 port map( A1 => A(25), A2 => n110, B1 => B(25), B2 => n107, 
                           ZN => n170);
   U61 : INV_X1 port map( A => n171, ZN => Y(26));
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n109, B1 => B(26), B2 => n107, 
                           ZN => n171);
   U63 : INV_X1 port map( A => n172, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n110, B1 => B(27), B2 => n107, 
                           ZN => n172);
   U65 : INV_X1 port map( A => n173, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n109, B1 => B(28), B2 => n107, 
                           ZN => n173);
   U67 : INV_X1 port map( A => n174, ZN => Y(29));
   U68 : AOI22_X1 port map( A1 => A(29), A2 => n110, B1 => B(29), B2 => n107, 
                           ZN => n174);
   U69 : INV_X1 port map( A => n175, ZN => Y(30));
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n109, B1 => B(30), B2 => n107, 
                           ZN => n175);
   U71 : INV_X1 port map( A => n176, ZN => Y(31));
   U72 : AOI22_X1 port map( A1 => A(31), A2 => n110, B1 => n107, B2 => B(31), 
                           ZN => n176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_6 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_6;

architecture SYN_Behavioral of REG_NBIT32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n215, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n215, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n215, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n215, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n215, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n215, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n215, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n215, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n215, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n215, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n215, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n215, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n216, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n216, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n216, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n216, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n216, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n216, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n216, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n206, Z => n214);
   U3 : BUF_X1 port map( A => n206, Z => n213);
   U4 : BUF_X1 port map( A => n219, Z => n218);
   U5 : BUF_X1 port map( A => n214, Z => n208);
   U6 : BUF_X1 port map( A => n214, Z => n207);
   U7 : BUF_X1 port map( A => n214, Z => n209);
   U8 : BUF_X1 port map( A => n213, Z => n211);
   U9 : BUF_X1 port map( A => n213, Z => n210);
   U10 : BUF_X1 port map( A => n218, Z => n216);
   U11 : BUF_X1 port map( A => n218, Z => n215);
   U12 : BUF_X1 port map( A => n218, Z => n217);
   U13 : BUF_X1 port map( A => n213, Z => n212);
   U14 : INV_X1 port map( A => reset, ZN => n219);
   U15 : BUF_X1 port map( A => enable, Z => n206);
   U16 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n251, ZN => n141);
   U17 : NAND2_X1 port map( A1 => n212, A2 => data_in(0), ZN => n251);
   U18 : OAI21_X1 port map( B1 => n172, B2 => n209, A => n250, ZN => n140);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n207, ZN => n250);
   U20 : OAI21_X1 port map( B1 => n171, B2 => n209, A => n249, ZN => n139);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n207, ZN => n249);
   U22 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n248, ZN => n138);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n207, ZN => n248);
   U24 : OAI21_X1 port map( B1 => n169, B2 => n209, A => n247, ZN => n137);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n207, ZN => n247);
   U26 : OAI21_X1 port map( B1 => n168, B2 => n209, A => n246, ZN => n136);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n208, ZN => n246);
   U28 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n245, ZN => n135);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n208, ZN => n245);
   U30 : OAI21_X1 port map( B1 => n166, B2 => n209, A => n244, ZN => n134);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n208, ZN => n244);
   U32 : OAI21_X1 port map( B1 => n165, B2 => n210, A => n243, ZN => n133);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n208, ZN => n243);
   U34 : OAI21_X1 port map( B1 => n164, B2 => n210, A => n242, ZN => n132);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n209, ZN => n242);
   U36 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n241, ZN => n131);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n208, ZN => n241);
   U38 : OAI21_X1 port map( B1 => n162, B2 => n210, A => n240, ZN => n130);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n209, ZN => n240);
   U40 : OAI21_X1 port map( B1 => n161, B2 => n210, A => n239, ZN => n129);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n209, ZN => n239);
   U42 : OAI21_X1 port map( B1 => n160, B2 => n210, A => n238, ZN => n128);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n209, ZN => n238);
   U44 : OAI21_X1 port map( B1 => n159, B2 => n210, A => n237, ZN => n127);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n209, ZN => n237);
   U46 : OAI21_X1 port map( B1 => n158, B2 => n210, A => n236, ZN => n126);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n209, ZN => n236);
   U48 : OAI21_X1 port map( B1 => n157, B2 => n211, A => n235, ZN => n125);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n209, ZN => n235);
   U50 : OAI21_X1 port map( B1 => n156, B2 => n211, A => n234, ZN => n124);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n208, ZN => n234);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n211, A => n233, ZN => n123);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n208, ZN => n233);
   U54 : OAI21_X1 port map( B1 => n154, B2 => n211, A => n232, ZN => n122);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n208, ZN => n232);
   U56 : OAI21_X1 port map( B1 => n153, B2 => n211, A => n231, ZN => n121);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n208, ZN => n231);
   U58 : OAI21_X1 port map( B1 => n152, B2 => n211, A => n230, ZN => n120);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n208, ZN => n230);
   U60 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n229, ZN => n119);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n208, ZN => n229);
   U62 : OAI21_X1 port map( B1 => n150, B2 => n211, A => n228, ZN => n118);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n208, ZN => n228);
   U64 : OAI21_X1 port map( B1 => n149, B2 => n211, A => n227, ZN => n117);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n207, ZN => n227);
   U66 : OAI21_X1 port map( B1 => n148, B2 => n211, A => n226, ZN => n116);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n207, ZN => n226);
   U68 : OAI21_X1 port map( B1 => n147, B2 => n211, A => n225, ZN => n115);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n207, ZN => n225);
   U70 : OAI21_X1 port map( B1 => n146, B2 => n211, A => n224, ZN => n114);
   U71 : NAND2_X1 port map( A1 => data_in(27), A2 => n207, ZN => n224);
   U72 : OAI21_X1 port map( B1 => n145, B2 => n212, A => n223, ZN => n113);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n207, ZN => n223);
   U74 : OAI21_X1 port map( B1 => n144, B2 => n212, A => n222, ZN => n112);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n207, ZN => n222);
   U76 : OAI21_X1 port map( B1 => n143, B2 => n212, A => n221, ZN => n111);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n207, ZN => n221);
   U78 : OAI21_X1 port map( B1 => n142, B2 => n210, A => n220, ZN => n110);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n207, ZN => n220);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_1;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n6, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_2;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n6, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_3;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n6, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_6;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n6, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_7;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n6, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_8;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U3 : INV_X1 port map( A => n8, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U5 : INV_X1 port map( A => n7, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U7 : INV_X1 port map( A => n6, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U9 : INV_X1 port map( A => SEL, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_10;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n9, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U4 : INV_X1 port map( A => n8, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U6 : INV_X1 port map( A => n7, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_11;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n9, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U4 : INV_X1 port map( A => n8, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U6 : INV_X1 port map( A => n7, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_17;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n6, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n9, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U8 : INV_X1 port map( A => n8, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_27;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n9, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_33;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n6, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U4 : INV_X1 port map( A => n9, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n7, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_40;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n6, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_43;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n9, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_44;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n9, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_47;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n9, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_48;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => Y(2));
   U2 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U3 : INV_X1 port map( A => n8, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U5 : INV_X1 port map( A => n9, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U7 : INV_X1 port map( A => SEL, ZN => n18);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_54;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n9, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U4 : INV_X1 port map( A => n8, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U6 : INV_X1 port map( A => n7, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U8 : INV_X1 port map( A => n6, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_55;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n6, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U4 : INV_X1 port map( A => n9, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n7, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_56;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U4 : INV_X1 port map( A => n7, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U6 : INV_X1 port map( A => n6, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_1;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_1 is

   component MUX2to1_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1076, n_1077 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1076);
   RCA0 : RCAN_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1077);
   MUX21 : MUX2to1_NBIT4_1 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_2;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_2 is

   component MUX2to1_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1078, n_1079 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1078);
   RCA0 : RCAN_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1079);
   MUX21 : MUX2to1_NBIT4_2 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_3;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_3 is

   component MUX2to1_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1080, n_1081 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1080);
   RCA0 : RCAN_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1081);
   MUX21 : MUX2to1_NBIT4_3 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_6;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_6 is

   component MUX2to1_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1082, n_1083 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1082);
   RCA0 : RCAN_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1083);
   MUX21 : MUX2to1_NBIT4_6 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_7;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_7 is

   component MUX2to1_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1084, n_1085 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1084);
   RCA0 : RCAN_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1085);
   MUX21 : MUX2to1_NBIT4_7 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_8;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_8 is

   component MUX2to1_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1086, n_1087 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1086);
   RCA0 : RCAN_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1087);
   MUX21 : MUX2to1_NBIT4_8 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_1;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U2 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U3 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U4 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U5 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U6 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U7 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U8 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U9 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U10 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U11 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U14 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U18 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U20 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U21 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U22 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U23 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U24 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U25 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U26 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U27 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U28 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U29 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U30 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U31 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_10;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_10 is

   component MUX2to1_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1088, n_1089 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1088);
   RCA0 : RCAN_NBIT4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1089);
   MUX21 : MUX2to1_NBIT4_10 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_11;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_11 is

   component MUX2to1_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1090, n_1091 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1090);
   RCA0 : RCAN_NBIT4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1091);
   MUX21 : MUX2to1_NBIT4_11 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_2;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U2 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U3 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U4 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U5 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U6 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U7 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U8 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U9 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U10 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U11 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U14 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U18 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U20 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U21 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U22 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U23 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U24 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U25 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U26 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U27 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U28 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U29 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U30 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U31 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_17;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_17 is

   component MUX2to1_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1092, n_1093 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_34 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1092);
   RCA0 : RCAN_NBIT4_33 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1093);
   MUX21 : MUX2to1_NBIT4_17 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_3;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U2 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U3 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U4 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U5 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U6 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U7 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U8 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U9 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U10 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U11 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U12 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U13 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U14 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U18 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U19 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U20 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U21 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U22 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U23 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U24 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U25 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U26 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U27 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U28 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U29 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U30 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_27;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_27 is

   component MUX2to1_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1094, n_1095 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_54 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1094);
   RCA0 : RCAN_NBIT4_53 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1095);
   MUX21 : MUX2to1_NBIT4_27 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_4;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U3 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U4 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U5 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U6 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U7 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U8 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U9 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U10 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U11 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U12 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U13 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U14 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U15 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U16 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U17 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U18 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U19 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U20 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U21 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U22 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U23 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U24 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U25 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U26 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U27 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U28 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U29 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U30 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_33;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_33 is

   component MUX2to1_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_65
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_66
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1096, n_1097 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_66 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1096);
   RCA0 : RCAN_NBIT4_65 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1097);
   MUX21 : MUX2to1_NBIT4_33 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_40;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_40 is

   component MUX2to1_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_79
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_80
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1098, n_1099 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_80 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1098);
   RCA0 : RCAN_NBIT4_79 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1099);
   MUX21 : MUX2to1_NBIT4_40 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_38 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_38;

architecture SYN_BEHAVIORAL of G_block_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_125 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_125;

architecture SYN_BEHAVIORAL of PG_block_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_5;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U2 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U3 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U4 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U5 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U6 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U7 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U8 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U9 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U10 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U11 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U12 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U13 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U14 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U18 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U19 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U20 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U21 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U22 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U23 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U24 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U25 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U26 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U27 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U28 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U29 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U30 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_43;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_43 is

   component MUX2to1_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_85
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_86
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1100, n_1101 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_86 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1100);
   RCA0 : RCAN_NBIT4_85 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1101);
   MUX21 : MUX2to1_NBIT4_43 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_44;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_44 is

   component MUX2to1_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_87
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_88
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1102, n_1103 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_88 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1102);
   RCA0 : RCAN_NBIT4_87 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1103);
   MUX21 : MUX2to1_NBIT4_44 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_47;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_47 is

   component MUX2to1_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_93
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_94
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1104, n_1105 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_94 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1104);
   RCA0 : RCAN_NBIT4_93 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1105);
   MUX21 : MUX2to1_NBIT4_47 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_48;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_48 is

   component MUX2to1_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_95
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_96
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1106, n_1107 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_96 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1106);
   RCA0 : RCAN_NBIT4_95 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1107);
   MUX21 : MUX2to1_NBIT4_48 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_50 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_50;

architecture SYN_BEHAVIORAL of G_block_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_52 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_52;

architecture SYN_BEHAVIORAL of G_block_52 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_6;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U3 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U4 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U5 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U6 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U7 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U8 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U9 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U10 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U11 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U12 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U13 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U14 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U15 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U16 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U17 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U18 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U19 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U20 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U21 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U22 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U23 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U24 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U25 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U26 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U27 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U28 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U29 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U30 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_54;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_54 is

   component MUX2to1_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_107
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_108
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1108, n_1109 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_108 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1108);
   RCA0 : RCAN_NBIT4_107 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1109);
   MUX21 : MUX2to1_NBIT4_54 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_55;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_55 is

   component MUX2to1_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_109
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_110
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1110, n_1111 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_110 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1110);
   RCA0 : RCAN_NBIT4_109 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1111);
   MUX21 : MUX2to1_NBIT4_55 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_56;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_56 is

   component MUX2to1_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_111
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_112
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1112, n_1113 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_112 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1112);
   RCA0 : RCAN_NBIT4_111 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1113);
   MUX21 : MUX2to1_NBIT4_56 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_7;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U2 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U3 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U4 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U5 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U6 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U7 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U8 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U9 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U10 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U11 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U14 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U18 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U20 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U21 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U22 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U23 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U24 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U25 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U26 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U27 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U28 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U29 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U30 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U31 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_57;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_58;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_59;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_61;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_62;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_63;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n18 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n18);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n18, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n18, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n18, B1 => B(0), B2 => SEL, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_0;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n14 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n14);
   U2 : INV_X1 port map( A => n6, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n14, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U4 : INV_X1 port map( A => n9, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n14, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n14, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : INV_X1 port map( A => n7, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n14, B1 => B(2), B2 => SEL, ZN => 
                           n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_127 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_127;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_127 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_0;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 is

   component CARRY_SEL_N_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_1
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_2
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_3
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_4
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_1
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_2
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_5
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_6
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_3
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_4
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_5
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_7
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_6
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_7
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_8
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_9
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_10
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_11
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_12
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_8
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_13
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_14
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_15
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_16
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_17
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_18
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_19
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_20
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_21
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_22
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_23
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_24
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_25
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_26
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_27
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_9
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n5, n3, n4, n7, n8, n_1114 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_1 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1114, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_9 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B 
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_27 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_26 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_25 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_24 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_23 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_22 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_21 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_20 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_19 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_18 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_17 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_16 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_15 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_14 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_13 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_8 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B 
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_12 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_11 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_10 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_9 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_8 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_7 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_6 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_7 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B 
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_5 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_4 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_3 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_6 port map( A(1) => P_12_9_port, A(0) => G_12_9_port, 
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_5 port map( A(1) => P_16_9_port, A(0) => G_16_9_port, 
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_2 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_1 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_4 port map( A(1) => P_20_17_port, A(0) => G_20_17_port
                           , B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_3 port map( A(1) => P_24_17_port, A(0) => G_24_17_port
                           , B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_2 port map( A(1) => P_28_17_port, A(0) => G_28_17_port
                           , B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_1 port map( A(1) => P_32_17_port, A(0) => G_32_17_port
                           , B => Co_4_port, Gout => Co_8_port);
   U1 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n8, ZN => n3);
   U2 : INV_X1 port map( A => n4, ZN => n8);
   U3 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n7, A2 => n3, ZN => G_1_0_port);
   U5 : INV_X1 port map( A => n5, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 is

   component CARRY_SEL_N_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_15 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_14 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_13 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_12 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_11 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_10 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_9 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_10
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_11
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_12
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_13
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_28
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_29
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_14
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_15
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_30
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_31
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_32
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_16
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_33
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_34
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_35
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_36
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_37
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_38
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_39
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_17
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_40
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_41
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_42
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_43
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_44
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_45
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_46
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_47
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_48
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_49
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_50
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_51
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_52
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_53
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_54
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_18
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n5, n3, n4, n7, n8, n_1115 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_2 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1115, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_18 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_54 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_53 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_52 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_51 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_50 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_49 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_48 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_47 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_46 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_45 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_44 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_43 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_42 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_41 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_40 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_17 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_39 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_38 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_37 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_36 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_35 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_34 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_33 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_16 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_32 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_31 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_30 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_15 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_14 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_29 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_28 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_13 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_12 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_11 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_10 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n8, ZN => n3);
   U2 : INV_X1 port map( A => n4, ZN => n8);
   U3 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n7, A2 => n3, ZN => G_1_0_port);
   U5 : INV_X1 port map( A => n5, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 is

   component CARRY_SEL_N_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_23 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_22 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_21 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_20 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_19 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_18 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_17 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_19
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_20
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_21
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_22
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_55
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_56
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_23
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_24
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_57
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_58
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_59
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_25
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_60
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_61
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_62
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_63
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_64
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_65
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_66
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_26
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_67
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_68
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_69
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_70
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_71
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_72
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_73
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_74
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_75
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_76
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_77
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_78
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_79
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_80
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_81
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_27
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n5, n3, n4, n7, n8, n_1116 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_3 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1116, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_27 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_81 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_80 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_79 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_78 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_77 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_76 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_75 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_74 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_73 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_72 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_71 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_70 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_69 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_68 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_67 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_26 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_66 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_65 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_64 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_63 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_62 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_61 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_60 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_25 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_59 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_58 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_57 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_24 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_23 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_56 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_55 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_22 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_21 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_20 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_19 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NOR2_X1 port map( A1 => n7, A2 => n3, ZN => G_1_0_port);
   U2 : INV_X1 port map( A => n5, ZN => n7);
   U3 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n8, ZN => n3);
   U4 : INV_X1 port map( A => n4, ZN => n8);
   U5 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 is

   component CARRY_SEL_N_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_31 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_30 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_29 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_28 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_27 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_26 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_25 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_28
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_29
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_30
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_31
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_82
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_83
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_32
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_33
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_84
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_85
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_86
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_34
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_87
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_88
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_89
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_90
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_91
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_92
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_93
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_35
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_94
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_95
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_96
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_97
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_98
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_99
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_100
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_101
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_102
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_103
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_104
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_105
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_106
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_107
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_108
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_36
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, n7,
      n8, G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, G_16_9_port, 
      G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, G_12_12_port, 
      G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, G_10_9_port, 
      G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, G_6_6_port, 
      G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, G_2_2_port, 
      G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, G_32_25_port, 
      G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, G_29_29_port, 
      G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, G_27_27_port, 
      G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, G_24_23_port, 
      G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, G_22_21_port, 
      G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, G_19_19_port, 
      G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, P_32_32_port, P_32_31_port, P_32_29_port, 
      P_32_25_port, P_32_17_port, P_31_31_port, P_30_30_port, P_30_29_port, 
      P_29_29_port, P_28_28_port, P_28_27_port, P_28_25_port, P_28_17_port, 
      P_27_27_port, P_26_26_port, P_26_25_port, P_25_25_port, P_24_24_port, 
      P_24_23_port, P_24_21_port, P_24_17_port, P_23_23_port, P_22_22_port, 
      P_22_21_port, P_21_21_port, P_20_20_port, P_20_19_port, P_20_17_port, 
      P_19_19_port, P_18_18_port, P_18_17_port, P_17_17_port, n5, n3, n4, n9, 
      n10, n_1117 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, n7
      , n8, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_4 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1117, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_36 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_108 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_107 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_106 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_105 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_104 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_103 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_102 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_101 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_100 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_99 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_98 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_97 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_96 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_95 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_94 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_35 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => n8);
   pgblock1_2_2 : PG_block_93 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_92 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_91 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_90 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_89 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_88 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_87 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_34 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => n8, Gout => n7);
   pgblock1_3_2 : PG_block_86 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_85 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_84 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_33 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => n7, Gout => Co_3_port);
   gblock2_4_4 : G_block_32 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => n7, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_83 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_82 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_31 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_30 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_29 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_28 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NOR2_X1 port map( A1 => n9, A2 => n3, ZN => G_1_0_port);
   U2 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n10, ZN => n3);
   U3 : INV_X1 port map( A => n5, ZN => n9);
   U4 : INV_X1 port map( A => n4, ZN => n10);
   U5 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 is

   component CARRY_SEL_N_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_39 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_38 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_37 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_36 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_35 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_34 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_33 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_37
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_38
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_39
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_40
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_109
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_110
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_41
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_42
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_111
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_112
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_113
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_43
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_114
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_115
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_116
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_117
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_118
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_119
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_120
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_44
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_121
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_122
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_123
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_124
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_125
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_126
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_127
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_128
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_129
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_130
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_131
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_132
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_133
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_134
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_135
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_45
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n5, n3, n4, n7, n8, n_1118 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_5 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1118, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_45 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_135 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_134 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_133 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_132 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_131 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_130 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_129 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_128 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_127 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_126 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_125 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_124 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_123 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_122 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_121 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_44 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_120 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_119 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_118 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_117 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_116 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_115 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_114 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_43 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_113 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_112 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_111 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_42 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_41 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_110 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_109 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_40 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_39 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_38 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_37 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NOR2_X1 port map( A1 => n7, A2 => n3, ZN => G_1_0_port);
   U2 : INV_X1 port map( A => n5, ZN => n7);
   U3 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n8, ZN => n3);
   U4 : INV_X1 port map( A => n4, ZN => n8);
   U5 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 is

   component CARRY_SEL_N_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_47 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_46 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_45 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_44 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_43 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_42 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_41 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_46
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_47
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_48
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_49
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_136
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_137
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_50
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_51
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_138
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_139
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_140
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_52
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_141
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_142
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_143
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_144
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_145
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_146
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_147
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_53
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_148
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_149
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_150
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_151
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_152
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_153
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_154
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_155
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_156
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_157
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_158
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_159
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_160
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_161
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_162
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_54
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n3, n4, n5, n6, n7, n_1119 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_6 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1119, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n3);
   gblock1_1_1 : G_block_54 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_162 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_161 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_160 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_159 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_158 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_157 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_156 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_155 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_154 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_153 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_152 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_151 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_150 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_149 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_148 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_53 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_147 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_146 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_145 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_144 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_143 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_142 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_141 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_52 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_140 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_139 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_138 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_51 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_50 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_137 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_136 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_49 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_48 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_47 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_46 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NOR2_X1 port map( A1 => n6, A2 => n4, ZN => G_1_0_port);
   U2 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n7, ZN => n4);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : INV_X1 port map( A => n5, ZN => n7);
   U5 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n5);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 is

   component CARRY_SEL_N_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_55 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_54 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_53 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_52 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_51 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_50 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_49 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_55
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_56
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_57
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_58
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_163
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_164
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_59
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_60
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_165
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_166
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_167
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_61
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_168
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_169
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_170
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_171
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_172
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_173
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_174
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_62
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_175
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_176
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_177
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_178
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_179
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_180
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_181
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_182
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_183
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_184
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_185
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_186
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_187
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_188
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_189
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_63
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n5, n3, n4, n7, n8, n_1120 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_7 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1120, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_63 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_189 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_188 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_187 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_186 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_185 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_184 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_183 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_182 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_181 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_180 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_179 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_178 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_177 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_176 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_175 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_62 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_174 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_173 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_172 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_171 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_170 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_169 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_168 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_61 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_167 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_166 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_165 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_60 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_59 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_164 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_163 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_58 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_57 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_56 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_55 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n8, ZN => n3);
   U2 : INV_X1 port map( A => n4, ZN => n8);
   U3 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n7, A2 => n3, ZN => G_1_0_port);
   U5 : INV_X1 port map( A => n5, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_57;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_57 is

   component MUX2to1_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_113
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_114
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1121, n_1122 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_114 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1121);
   RCA0 : RCAN_NBIT4_113 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1122);
   MUX21 : MUX2to1_NBIT4_57 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_58;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_58 is

   component MUX2to1_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_115
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_116
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1123, n_1124 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_116 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1123);
   RCA0 : RCAN_NBIT4_115 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1124);
   MUX21 : MUX2to1_NBIT4_58 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_59;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_59 is

   component MUX2to1_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_117
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_118
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1125, n_1126 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_118 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1125);
   RCA0 : RCAN_NBIT4_117 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1126);
   MUX21 : MUX2to1_NBIT4_59 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_61;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_61 is

   component MUX2to1_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_121
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_122
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1127, n_1128 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_122 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1127);
   RCA0 : RCAN_NBIT4_121 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1128);
   MUX21 : MUX2to1_NBIT4_61 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_62;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_62 is

   component MUX2to1_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_123
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_124
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1129, n_1130 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_124 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1129);
   RCA0 : RCAN_NBIT4_123 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1130);
   MUX21 : MUX2to1_NBIT4_62 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_63;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_63 is

   component MUX2to1_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_125
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_126
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1131, n_1132 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_126 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1131);
   RCA0 : RCAN_NBIT4_125 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1132);
   MUX21 : MUX2to1_NBIT4_63 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_0;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_0 is

   component MUX2to1_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_127
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1133, n_1134 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1133);
   RCA0 : RCAN_NBIT4_127 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1134);
   MUX21 : MUX2to1_NBIT4_0 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_191 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_191;

architecture SYN_BEHAVIORAL of PG_block_191 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_193 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_193;

architecture SYN_BEHAVIORAL of PG_block_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_201 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_201;

architecture SYN_BEHAVIORAL of PG_block_201 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_71 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_71;

architecture SYN_BEHAVIORAL of G_block_71 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_212 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_212;

architecture SYN_BEHAVIORAL of PG_block_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_214 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_214;

architecture SYN_BEHAVIORAL of PG_block_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_215 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_215;

architecture SYN_BEHAVIORAL of PG_block_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_0 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_0;

architecture SYN_BEHAVIORAL of PG_block_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_0 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_0;

architecture SYN_BEHAVIORAL of G_block_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_0;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U2 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U3 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U4 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U5 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U6 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U7 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U8 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U9 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U10 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U11 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U12 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U13 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U14 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U15 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U16 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U17 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U18 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U19 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U20 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U21 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U22 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U23 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U24 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U25 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U26 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U27 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U28 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U29 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U30 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U31 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_1 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_1;

architecture SYN_Behavioral of REG_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n199, n200, n201, n202 : std_logic;

begin
   
   reg_reg_27_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n200, Q => 
                           data_out(27), QN => n139);
   reg_reg_26_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n201, Q => 
                           data_out(26), QN => n140);
   reg_reg_25_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n200, Q => 
                           data_out(25), QN => n141);
   reg_reg_24_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n200, Q => 
                           data_out(24), QN => n142);
   reg_reg_23_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n201, Q => 
                           data_out(23), QN => n143);
   reg_reg_22_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n201, Q => 
                           data_out(22), QN => n144);
   reg_reg_21_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n201, Q => 
                           data_out(21), QN => n145);
   reg_reg_20_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n200, Q => 
                           data_out(20), QN => n146);
   reg_reg_19_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n199, Q => 
                           data_out(19), QN => n147);
   reg_reg_18_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n199, Q => 
                           data_out(18), QN => n148);
   reg_reg_17_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n199, Q => 
                           data_out(17), QN => n149);
   reg_reg_16_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n199, Q => 
                           data_out(16), QN => n150);
   reg_reg_15_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n199, Q => 
                           data_out(15), QN => n151);
   reg_reg_14_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n199, Q => 
                           data_out(14), QN => n152);
   reg_reg_13_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n199, Q => 
                           data_out(13), QN => n153);
   reg_reg_12_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n199, Q => 
                           data_out(12), QN => n154);
   reg_reg_11_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n199, Q => 
                           data_out(11), QN => n155);
   reg_reg_10_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n199, Q => 
                           data_out(10), QN => n156);
   reg_reg_9_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n199, Q => 
                           data_out(9), QN => n157);
   reg_reg_8_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n199, Q => 
                           data_out(8), QN => n158);
   reg_reg_7_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n200, Q => 
                           data_out(7), QN => n159);
   reg_reg_6_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n200, Q => 
                           data_out(6), QN => n160);
   reg_reg_5_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n200, Q => 
                           data_out(5), QN => n161);
   reg_reg_4_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n200, Q => 
                           data_out(4), QN => n162);
   reg_reg_3_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n200, Q => 
                           data_out(3), QN => n163);
   reg_reg_2_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n200, Q => 
                           data_out(2), QN => n164);
   reg_reg_1_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n200, Q => 
                           data_out(1), QN => n165);
   reg_reg_0_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n200, Q => 
                           data_out(0), QN => n166);
   reg_reg_31_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n201, Q => 
                           data_out(31), QN => n135);
   reg_reg_29_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n201, Q => 
                           data_out(29), QN => n137);
   reg_reg_28_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n201, Q => 
                           data_out(28), QN => n138);
   reg_reg_30_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n201, Q => 
                           data_out(30), QN => n136);
   U2 : BUF_X1 port map( A => n202, Z => n199);
   U3 : BUF_X1 port map( A => n202, Z => n200);
   U4 : BUF_X1 port map( A => n202, Z => n201);
   U5 : OAI21_X1 port map( B1 => n135, B2 => enable, A => n33, ZN => n103);
   U6 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n33);
   U7 : OAI21_X1 port map( B1 => n136, B2 => enable, A => n32, ZN => n104);
   U8 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n138, B2 => enable, A => n30, ZN => n106);
   U10 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n30);
   U11 : OAI21_X1 port map( B1 => n137, B2 => enable, A => n31, ZN => n105);
   U12 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n31);
   U13 : OAI21_X1 port map( B1 => n139, B2 => enable, A => n29, ZN => n107);
   U14 : NAND2_X1 port map( A1 => data_in(27), A2 => enable, ZN => n29);
   U15 : OAI21_X1 port map( B1 => n142, B2 => enable, A => n26, ZN => n110);
   U16 : NAND2_X1 port map( A1 => data_in(24), A2 => enable, ZN => n26);
   U17 : OAI21_X1 port map( B1 => n141, B2 => enable, A => n27, ZN => n109);
   U18 : NAND2_X1 port map( A1 => data_in(25), A2 => enable, ZN => n27);
   U19 : OAI21_X1 port map( B1 => n140, B2 => enable, A => n28, ZN => n108);
   U20 : NAND2_X1 port map( A1 => data_in(26), A2 => enable, ZN => n28);
   U21 : OAI21_X1 port map( B1 => n143, B2 => enable, A => n25, ZN => n111);
   U22 : NAND2_X1 port map( A1 => data_in(23), A2 => enable, ZN => n25);
   U23 : OAI21_X1 port map( B1 => n146, B2 => enable, A => n22, ZN => n114);
   U24 : NAND2_X1 port map( A1 => data_in(20), A2 => enable, ZN => n22);
   U25 : OAI21_X1 port map( B1 => n145, B2 => enable, A => n23, ZN => n113);
   U26 : NAND2_X1 port map( A1 => data_in(21), A2 => enable, ZN => n23);
   U27 : OAI21_X1 port map( B1 => n144, B2 => enable, A => n24, ZN => n112);
   U28 : NAND2_X1 port map( A1 => data_in(22), A2 => enable, ZN => n24);
   U29 : OAI21_X1 port map( B1 => n147, B2 => enable, A => n21, ZN => n115);
   U30 : NAND2_X1 port map( A1 => data_in(19), A2 => enable, ZN => n21);
   U31 : OAI21_X1 port map( B1 => n150, B2 => enable, A => n18, ZN => n118);
   U32 : NAND2_X1 port map( A1 => data_in(16), A2 => enable, ZN => n18);
   U33 : OAI21_X1 port map( B1 => n149, B2 => enable, A => n19, ZN => n117);
   U34 : NAND2_X1 port map( A1 => data_in(17), A2 => enable, ZN => n19);
   U35 : OAI21_X1 port map( B1 => n148, B2 => enable, A => n20, ZN => n116);
   U36 : NAND2_X1 port map( A1 => data_in(18), A2 => enable, ZN => n20);
   U37 : OAI21_X1 port map( B1 => n151, B2 => enable, A => n17, ZN => n119);
   U38 : NAND2_X1 port map( A1 => data_in(15), A2 => enable, ZN => n17);
   U39 : OAI21_X1 port map( B1 => n154, B2 => enable, A => n14, ZN => n122);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => enable, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n153, B2 => enable, A => n15, ZN => n121);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => enable, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n152, B2 => enable, A => n16, ZN => n120);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => enable, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n155, B2 => enable, A => n13, ZN => n123);
   U46 : NAND2_X1 port map( A1 => data_in(11), A2 => enable, ZN => n13);
   U47 : OAI21_X1 port map( B1 => n156, B2 => enable, A => n12, ZN => n124);
   U48 : NAND2_X1 port map( A1 => data_in(10), A2 => enable, ZN => n12);
   U49 : OAI21_X1 port map( B1 => n158, B2 => enable, A => n10, ZN => n126);
   U50 : NAND2_X1 port map( A1 => data_in(8), A2 => enable, ZN => n10);
   U51 : OAI21_X1 port map( B1 => n157, B2 => enable, A => n11, ZN => n125);
   U52 : NAND2_X1 port map( A1 => data_in(9), A2 => enable, ZN => n11);
   U53 : OAI21_X1 port map( B1 => n159, B2 => enable, A => n9, ZN => n127);
   U54 : NAND2_X1 port map( A1 => data_in(7), A2 => enable, ZN => n9);
   U55 : OAI21_X1 port map( B1 => n160, B2 => enable, A => n8, ZN => n128);
   U56 : NAND2_X1 port map( A1 => data_in(6), A2 => enable, ZN => n8);
   U57 : OAI21_X1 port map( B1 => n162, B2 => enable, A => n6, ZN => n130);
   U58 : NAND2_X1 port map( A1 => data_in(4), A2 => enable, ZN => n6);
   U59 : OAI21_X1 port map( B1 => n161, B2 => enable, A => n7, ZN => n129);
   U60 : NAND2_X1 port map( A1 => data_in(5), A2 => enable, ZN => n7);
   U61 : OAI21_X1 port map( B1 => n163, B2 => enable, A => n5, ZN => n131);
   U62 : NAND2_X1 port map( A1 => data_in(3), A2 => enable, ZN => n5);
   U63 : OAI21_X1 port map( B1 => n164, B2 => enable, A => n4, ZN => n132);
   U64 : NAND2_X1 port map( A1 => data_in(2), A2 => enable, ZN => n4);
   U65 : OAI21_X1 port map( B1 => n165, B2 => enable, A => n3, ZN => n133);
   U66 : NAND2_X1 port map( A1 => data_in(1), A2 => enable, ZN => n3);
   U67 : OAI21_X1 port map( B1 => n166, B2 => enable, A => n2, ZN => n134);
   U68 : NAND2_X1 port map( A1 => enable, A2 => data_in(0), ZN => n2);
   U69 : INV_X1 port map( A => reset, ZN => n202);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_4 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_4;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_2 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_2;

architecture SYN_Behavioral of REG_NBIT32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n197, n198, n199, n200 : std_logic;

begin
   
   reg_reg_19_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n197, Q => 
                           data_out(19), QN => n145);
   reg_reg_18_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n197, Q => 
                           data_out(18), QN => n146);
   reg_reg_17_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n197, Q => 
                           data_out(17), QN => n147);
   reg_reg_16_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n197, Q => 
                           data_out(16), QN => n148);
   reg_reg_15_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n197, Q => 
                           data_out(15), QN => n149);
   reg_reg_14_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n197, Q => 
                           data_out(14), QN => n150);
   reg_reg_13_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n197, Q => 
                           data_out(13), QN => n151);
   reg_reg_12_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n197, Q => 
                           data_out(12), QN => n152);
   reg_reg_11_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n197, Q => 
                           data_out(11), QN => n153);
   reg_reg_10_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n197, Q => 
                           data_out(10), QN => n154);
   reg_reg_9_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n197, Q => 
                           data_out(9), QN => n155);
   reg_reg_8_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n197, Q => 
                           data_out(8), QN => n156);
   reg_reg_7_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n198, Q => 
                           data_out(7), QN => n157);
   reg_reg_6_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n198, Q => 
                           data_out(6), QN => n158);
   reg_reg_5_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n198, Q => 
                           data_out(5), QN => n159);
   reg_reg_4_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n198, Q => 
                           data_out(4), QN => n160);
   reg_reg_3_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n198, Q => 
                           data_out(3), QN => n161);
   reg_reg_2_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n198, Q => 
                           data_out(2), QN => n162);
   reg_reg_1_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n198, Q => 
                           data_out(1), QN => n163);
   reg_reg_0_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n198, Q => 
                           data_out(0), QN => n164);
   reg_reg_22_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n198, Q => 
                           data_out(22), QN => n142);
   reg_reg_21_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n198, Q => 
                           data_out(21), QN => n143);
   reg_reg_20_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n198, Q => 
                           data_out(20), QN => n144);
   reg_reg_26_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n198, Q => 
                           data_out(26), QN => n138);
   reg_reg_25_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n199, Q => 
                           data_out(25), QN => n139);
   reg_reg_24_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n199, Q => 
                           data_out(24), QN => n140);
   reg_reg_23_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n199, Q => 
                           data_out(23), QN => n141);
   reg_reg_27_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n199, Q => 
                           data_out(27), QN => n137);
   reg_reg_30_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n199, Q => 
                           data_out(30), QN => n134);
   reg_reg_29_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n199, Q => 
                           data_out(29), QN => n135);
   reg_reg_28_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n199, Q => 
                           data_out(28), QN => n136);
   reg_reg_31_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n199, Q => 
                           data_out(31), QN => n133);
   U2 : BUF_X1 port map( A => n200, Z => n198);
   U3 : BUF_X1 port map( A => n200, Z => n197);
   U4 : BUF_X1 port map( A => n200, Z => n199);
   U5 : OAI21_X1 port map( B1 => n133, B2 => enable, A => n33, ZN => n101);
   U6 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n33);
   U7 : OAI21_X1 port map( B1 => n136, B2 => enable, A => n30, ZN => n104);
   U8 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n30);
   U9 : OAI21_X1 port map( B1 => n135, B2 => enable, A => n31, ZN => n103);
   U10 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n31);
   U11 : OAI21_X1 port map( B1 => n134, B2 => enable, A => n32, ZN => n102);
   U12 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n32);
   U13 : OAI21_X1 port map( B1 => n137, B2 => enable, A => n29, ZN => n105);
   U14 : NAND2_X1 port map( A1 => data_in(27), A2 => enable, ZN => n29);
   U15 : OAI21_X1 port map( B1 => n140, B2 => enable, A => n26, ZN => n108);
   U16 : NAND2_X1 port map( A1 => data_in(24), A2 => enable, ZN => n26);
   U17 : OAI21_X1 port map( B1 => n139, B2 => enable, A => n27, ZN => n107);
   U18 : NAND2_X1 port map( A1 => data_in(25), A2 => enable, ZN => n27);
   U19 : OAI21_X1 port map( B1 => n138, B2 => enable, A => n28, ZN => n106);
   U20 : NAND2_X1 port map( A1 => data_in(26), A2 => enable, ZN => n28);
   U21 : OAI21_X1 port map( B1 => n141, B2 => enable, A => n25, ZN => n109);
   U22 : NAND2_X1 port map( A1 => data_in(23), A2 => enable, ZN => n25);
   U23 : OAI21_X1 port map( B1 => n144, B2 => enable, A => n22, ZN => n112);
   U24 : NAND2_X1 port map( A1 => data_in(20), A2 => enable, ZN => n22);
   U25 : OAI21_X1 port map( B1 => n143, B2 => enable, A => n23, ZN => n111);
   U26 : NAND2_X1 port map( A1 => data_in(21), A2 => enable, ZN => n23);
   U27 : OAI21_X1 port map( B1 => n142, B2 => enable, A => n24, ZN => n110);
   U28 : NAND2_X1 port map( A1 => data_in(22), A2 => enable, ZN => n24);
   U29 : OAI21_X1 port map( B1 => n145, B2 => enable, A => n21, ZN => n113);
   U30 : NAND2_X1 port map( A1 => data_in(19), A2 => enable, ZN => n21);
   U31 : OAI21_X1 port map( B1 => n148, B2 => enable, A => n18, ZN => n116);
   U32 : NAND2_X1 port map( A1 => data_in(16), A2 => enable, ZN => n18);
   U33 : OAI21_X1 port map( B1 => n147, B2 => enable, A => n19, ZN => n115);
   U34 : NAND2_X1 port map( A1 => data_in(17), A2 => enable, ZN => n19);
   U35 : OAI21_X1 port map( B1 => n146, B2 => enable, A => n20, ZN => n114);
   U36 : NAND2_X1 port map( A1 => data_in(18), A2 => enable, ZN => n20);
   U37 : OAI21_X1 port map( B1 => n149, B2 => enable, A => n17, ZN => n117);
   U38 : NAND2_X1 port map( A1 => data_in(15), A2 => enable, ZN => n17);
   U39 : OAI21_X1 port map( B1 => n152, B2 => enable, A => n14, ZN => n120);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => enable, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n151, B2 => enable, A => n15, ZN => n119);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => enable, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n150, B2 => enable, A => n16, ZN => n118);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => enable, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n153, B2 => enable, A => n13, ZN => n121);
   U46 : NAND2_X1 port map( A1 => data_in(11), A2 => enable, ZN => n13);
   U47 : OAI21_X1 port map( B1 => n154, B2 => enable, A => n12, ZN => n122);
   U48 : NAND2_X1 port map( A1 => data_in(10), A2 => enable, ZN => n12);
   U49 : OAI21_X1 port map( B1 => n156, B2 => enable, A => n10, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(8), A2 => enable, ZN => n10);
   U51 : OAI21_X1 port map( B1 => n155, B2 => enable, A => n11, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(9), A2 => enable, ZN => n11);
   U53 : OAI21_X1 port map( B1 => n157, B2 => enable, A => n9, ZN => n125);
   U54 : NAND2_X1 port map( A1 => data_in(7), A2 => enable, ZN => n9);
   U55 : OAI21_X1 port map( B1 => n158, B2 => enable, A => n8, ZN => n126);
   U56 : NAND2_X1 port map( A1 => data_in(6), A2 => enable, ZN => n8);
   U57 : OAI21_X1 port map( B1 => n160, B2 => enable, A => n6, ZN => n128);
   U58 : NAND2_X1 port map( A1 => data_in(4), A2 => enable, ZN => n6);
   U59 : OAI21_X1 port map( B1 => n159, B2 => enable, A => n7, ZN => n127);
   U60 : NAND2_X1 port map( A1 => data_in(5), A2 => enable, ZN => n7);
   U61 : OAI21_X1 port map( B1 => n161, B2 => enable, A => n5, ZN => n129);
   U62 : NAND2_X1 port map( A1 => data_in(3), A2 => enable, ZN => n5);
   U63 : OAI21_X1 port map( B1 => n162, B2 => enable, A => n4, ZN => n130);
   U64 : NAND2_X1 port map( A1 => data_in(2), A2 => enable, ZN => n4);
   U65 : OAI21_X1 port map( B1 => n163, B2 => enable, A => n3, ZN => n131);
   U66 : NAND2_X1 port map( A1 => data_in(1), A2 => enable, ZN => n3);
   U67 : OAI21_X1 port map( B1 => n164, B2 => enable, A => n2, ZN => n132);
   U68 : NAND2_X1 port map( A1 => enable, A2 => data_in(0), ZN => n2);
   U69 : INV_X1 port map( A => reset, ZN => n200);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_5 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_5;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_5 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_6 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_6;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_6 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_3 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_3;

architecture SYN_Behavioral of REG_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n197, n198, n199, n200 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n198, Q => 
                           data_out(31), QN => n133);
   reg_reg_30_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n198, Q => 
                           data_out(30), QN => n134);
   reg_reg_29_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n198, Q => 
                           data_out(29), QN => n135);
   reg_reg_28_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n198, Q => 
                           data_out(28), QN => n136);
   reg_reg_27_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n198, Q => 
                           data_out(27), QN => n137);
   reg_reg_26_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n198, Q => 
                           data_out(26), QN => n138);
   reg_reg_25_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n198, Q => 
                           data_out(25), QN => n139);
   reg_reg_24_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n198, Q => 
                           data_out(24), QN => n140);
   reg_reg_23_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n198, Q => 
                           data_out(23), QN => n141);
   reg_reg_22_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n198, Q => 
                           data_out(22), QN => n142);
   reg_reg_21_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n198, Q => 
                           data_out(21), QN => n143);
   reg_reg_20_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n198, Q => 
                           data_out(20), QN => n144);
   reg_reg_19_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n197, Q => 
                           data_out(19), QN => n145);
   reg_reg_18_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n197, Q => 
                           data_out(18), QN => n146);
   reg_reg_17_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n197, Q => 
                           data_out(17), QN => n147);
   reg_reg_16_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n197, Q => 
                           data_out(16), QN => n148);
   reg_reg_15_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n197, Q => 
                           data_out(15), QN => n149);
   reg_reg_14_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n197, Q => 
                           data_out(14), QN => n150);
   reg_reg_13_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n197, Q => 
                           data_out(13), QN => n151);
   reg_reg_12_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n197, Q => 
                           data_out(12), QN => n152);
   reg_reg_11_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n197, Q => 
                           data_out(11), QN => n153);
   reg_reg_10_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n197, Q => 
                           data_out(10), QN => n154);
   reg_reg_9_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n197, Q => 
                           data_out(9), QN => n155);
   reg_reg_8_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n197, Q => 
                           data_out(8), QN => n156);
   reg_reg_7_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n199, Q => 
                           data_out(7), QN => n157);
   reg_reg_6_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n199, Q => 
                           data_out(6), QN => n158);
   reg_reg_5_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n199, Q => 
                           data_out(5), QN => n159);
   reg_reg_4_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n199, Q => 
                           data_out(4), QN => n160);
   reg_reg_3_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n199, Q => 
                           data_out(3), QN => n161);
   reg_reg_2_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n199, Q => 
                           data_out(2), QN => n162);
   reg_reg_1_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n199, Q => 
                           data_out(1), QN => n163);
   reg_reg_0_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n199, Q => 
                           data_out(0), QN => n164);
   U2 : BUF_X1 port map( A => n200, Z => n197);
   U3 : BUF_X1 port map( A => n200, Z => n198);
   U4 : BUF_X1 port map( A => n200, Z => n199);
   U5 : OAI21_X1 port map( B1 => n145, B2 => enable, A => n21, ZN => n113);
   U6 : NAND2_X1 port map( A1 => data_in(19), A2 => enable, ZN => n21);
   U7 : OAI21_X1 port map( B1 => n157, B2 => enable, A => n9, ZN => n125);
   U8 : NAND2_X1 port map( A1 => data_in(7), A2 => enable, ZN => n9);
   U9 : OAI21_X1 port map( B1 => n156, B2 => enable, A => n10, ZN => n124);
   U10 : NAND2_X1 port map( A1 => data_in(8), A2 => enable, ZN => n10);
   U11 : OAI21_X1 port map( B1 => n155, B2 => enable, A => n11, ZN => n123);
   U12 : NAND2_X1 port map( A1 => data_in(9), A2 => enable, ZN => n11);
   U13 : OAI21_X1 port map( B1 => n154, B2 => enable, A => n12, ZN => n122);
   U14 : NAND2_X1 port map( A1 => data_in(10), A2 => enable, ZN => n12);
   U15 : OAI21_X1 port map( B1 => n153, B2 => enable, A => n13, ZN => n121);
   U16 : NAND2_X1 port map( A1 => data_in(11), A2 => enable, ZN => n13);
   U17 : OAI21_X1 port map( B1 => n149, B2 => enable, A => n17, ZN => n117);
   U18 : NAND2_X1 port map( A1 => data_in(15), A2 => enable, ZN => n17);
   U19 : OAI21_X1 port map( B1 => n148, B2 => enable, A => n18, ZN => n116);
   U20 : NAND2_X1 port map( A1 => data_in(16), A2 => enable, ZN => n18);
   U21 : OAI21_X1 port map( B1 => n147, B2 => enable, A => n19, ZN => n115);
   U22 : NAND2_X1 port map( A1 => data_in(17), A2 => enable, ZN => n19);
   U23 : OAI21_X1 port map( B1 => n146, B2 => enable, A => n20, ZN => n114);
   U24 : NAND2_X1 port map( A1 => data_in(18), A2 => enable, ZN => n20);
   U25 : OAI21_X1 port map( B1 => n141, B2 => enable, A => n25, ZN => n109);
   U26 : NAND2_X1 port map( A1 => data_in(23), A2 => enable, ZN => n25);
   U27 : OAI21_X1 port map( B1 => n137, B2 => enable, A => n29, ZN => n105);
   U28 : NAND2_X1 port map( A1 => data_in(27), A2 => enable, ZN => n29);
   U29 : OAI21_X1 port map( B1 => n133, B2 => enable, A => n33, ZN => n101);
   U30 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n33);
   U31 : OAI21_X1 port map( B1 => n160, B2 => enable, A => n6, ZN => n128);
   U32 : NAND2_X1 port map( A1 => data_in(4), A2 => enable, ZN => n6);
   U33 : OAI21_X1 port map( B1 => n159, B2 => enable, A => n7, ZN => n127);
   U34 : NAND2_X1 port map( A1 => data_in(5), A2 => enable, ZN => n7);
   U35 : OAI21_X1 port map( B1 => n158, B2 => enable, A => n8, ZN => n126);
   U36 : NAND2_X1 port map( A1 => data_in(6), A2 => enable, ZN => n8);
   U37 : OAI21_X1 port map( B1 => n152, B2 => enable, A => n14, ZN => n120);
   U38 : NAND2_X1 port map( A1 => data_in(12), A2 => enable, ZN => n14);
   U39 : OAI21_X1 port map( B1 => n151, B2 => enable, A => n15, ZN => n119);
   U40 : NAND2_X1 port map( A1 => data_in(13), A2 => enable, ZN => n15);
   U41 : OAI21_X1 port map( B1 => n150, B2 => enable, A => n16, ZN => n118);
   U42 : NAND2_X1 port map( A1 => data_in(14), A2 => enable, ZN => n16);
   U43 : OAI21_X1 port map( B1 => n144, B2 => enable, A => n22, ZN => n112);
   U44 : NAND2_X1 port map( A1 => data_in(20), A2 => enable, ZN => n22);
   U45 : OAI21_X1 port map( B1 => n143, B2 => enable, A => n23, ZN => n111);
   U46 : NAND2_X1 port map( A1 => data_in(21), A2 => enable, ZN => n23);
   U47 : OAI21_X1 port map( B1 => n142, B2 => enable, A => n24, ZN => n110);
   U48 : NAND2_X1 port map( A1 => data_in(22), A2 => enable, ZN => n24);
   U49 : OAI21_X1 port map( B1 => n140, B2 => enable, A => n26, ZN => n108);
   U50 : NAND2_X1 port map( A1 => data_in(24), A2 => enable, ZN => n26);
   U51 : OAI21_X1 port map( B1 => n139, B2 => enable, A => n27, ZN => n107);
   U52 : NAND2_X1 port map( A1 => data_in(25), A2 => enable, ZN => n27);
   U53 : OAI21_X1 port map( B1 => n138, B2 => enable, A => n28, ZN => n106);
   U54 : NAND2_X1 port map( A1 => data_in(26), A2 => enable, ZN => n28);
   U55 : OAI21_X1 port map( B1 => n136, B2 => enable, A => n30, ZN => n104);
   U56 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n30);
   U57 : OAI21_X1 port map( B1 => n135, B2 => enable, A => n31, ZN => n103);
   U58 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n31);
   U59 : OAI21_X1 port map( B1 => n134, B2 => enable, A => n32, ZN => n102);
   U60 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n32);
   U61 : OAI21_X1 port map( B1 => n163, B2 => enable, A => n3, ZN => n131);
   U62 : NAND2_X1 port map( A1 => data_in(1), A2 => enable, ZN => n3);
   U63 : OAI21_X1 port map( B1 => n162, B2 => enable, A => n4, ZN => n130);
   U64 : NAND2_X1 port map( A1 => data_in(2), A2 => enable, ZN => n4);
   U65 : OAI21_X1 port map( B1 => n161, B2 => enable, A => n5, ZN => n129);
   U66 : NAND2_X1 port map( A1 => data_in(3), A2 => enable, ZN => n5);
   U67 : OAI21_X1 port map( B1 => n164, B2 => enable, A => n2, ZN => n132);
   U68 : NAND2_X1 port map( A1 => enable, A2 => data_in(0), ZN => n2);
   U69 : INV_X1 port map( A => reset, ZN => n200);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_7 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_7;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_1 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_1;

architecture SYN_Behavioral of MUX5to1_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n188, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n187, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n188, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n189, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n188, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n187);
   U10 : BUF_X1 port map( A => n190, Z => n188);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U37 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U38 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U39 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U40 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U41 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U42 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U43 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U44 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U45 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U46 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U47 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U48 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U49 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U50 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U51 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U52 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U53 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U54 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U55 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U56 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U57 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U58 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U59 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179, 
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U60 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U61 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U62 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179, 
                           C1 => B(25), C2 => n175, ZN => n21);
   U63 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U64 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U65 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179, 
                           C1 => B(26), C2 => n175, ZN => n19);
   U66 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U67 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U68 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179, 
                           C1 => B(27), C2 => n175, ZN => n17);
   U69 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U70 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U71 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179, 
                           C1 => B(28), C2 => n175, ZN => n15);
   U72 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U73 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U74 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U75 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U76 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179, 
                           C1 => B(24), C2 => n175, ZN => n23);
   U77 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U78 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U79 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179, 
                           C1 => B(29), C2 => n175, ZN => n13);
   U80 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U81 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U82 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U83 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179, 
                           C1 => B(30), C2 => n175, ZN => n11);
   U84 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U85 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U86 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U87 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U88 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U89 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179, 
                           C1 => B(31), C2 => n175, ZN => n4);
   U90 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U91 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN 
                           => n70);
   U92 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, C1
                           => B(0), C2 => n177, ZN => n71);
   U93 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U94 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN 
                           => n68);
   U95 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, C1
                           => B(1), C2 => n177, ZN => n69);
   U96 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U97 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN 
                           => n66);
   U98 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, C1
                           => B(2), C2 => n177, ZN => n67);
   U99 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U100 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN
                           => n64);
   U101 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, 
                           C1 => B(3), C2 => n177, ZN => n65);
   U102 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U103 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN
                           => n62);
   U104 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, 
                           C1 => B(4), C2 => n177, ZN => n63);
   U105 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U106 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN
                           => n60);
   U107 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, 
                           C1 => B(5), C2 => n177, ZN => n61);
   U108 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U109 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN
                           => n58);
   U110 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, 
                           C1 => B(6), C2 => n177, ZN => n59);
   U111 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U112 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN
                           => n56_port);
   U113 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, 
                           C1 => B(7), C2 => n177, ZN => n57_port);
   U114 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U115 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN
                           => n54_port);
   U116 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, 
                           C1 => B(8), C2 => n176, ZN => n55_port);
   U117 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U118 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN
                           => n52_port);
   U119 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, 
                           C1 => B(9), C2 => n176, ZN => n53_port);
   U120 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U121 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U122 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180,
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U123 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U124 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U125 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180,
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U126 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U127 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U128 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180,
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U129 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U130 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U131 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180,
                           C1 => B(13), C2 => n176, ZN => n45_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_2 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_2;

architecture SYN_Behavioral of MUX5to1_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n188, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n187, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n188, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n188, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n187);
   U10 : BUF_X1 port map( A => n190, Z => n188);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U37 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U38 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U39 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U40 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U41 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U42 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U43 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U44 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U45 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U46 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U47 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U48 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U49 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U50 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U51 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U52 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U53 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U54 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U55 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U56 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U57 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U58 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U59 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U60 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U61 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U62 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179, 
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U63 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U64 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U65 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179, 
                           C1 => B(24), C2 => n175, ZN => n23);
   U66 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U67 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U68 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179, 
                           C1 => B(25), C2 => n175, ZN => n21);
   U69 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U70 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U71 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179, 
                           C1 => B(26), C2 => n175, ZN => n19);
   U72 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U73 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U74 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U75 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U76 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U77 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U78 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U79 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179, 
                           C1 => B(27), C2 => n175, ZN => n17);
   U80 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U81 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U82 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U83 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179, 
                           C1 => B(28), C2 => n175, ZN => n15);
   U84 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U85 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U86 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U87 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U88 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U89 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179, 
                           C1 => B(29), C2 => n175, ZN => n13);
   U90 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U91 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U92 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179, 
                           C1 => B(30), C2 => n175, ZN => n11);
   U93 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U94 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U95 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179, 
                           C1 => B(31), C2 => n175, ZN => n4);
   U96 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U97 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN 
                           => n70);
   U98 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, C1
                           => B(0), C2 => n177, ZN => n71);
   U99 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U100 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN
                           => n68);
   U101 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, 
                           C1 => B(1), C2 => n177, ZN => n69);
   U102 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U103 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN
                           => n66);
   U104 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, 
                           C1 => B(2), C2 => n177, ZN => n67);
   U105 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U106 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN
                           => n64);
   U107 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, 
                           C1 => B(3), C2 => n177, ZN => n65);
   U108 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U109 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN
                           => n62);
   U110 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, 
                           C1 => B(4), C2 => n177, ZN => n63);
   U111 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U112 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN
                           => n60);
   U113 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, 
                           C1 => B(5), C2 => n177, ZN => n61);
   U114 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U115 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN
                           => n58);
   U116 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, 
                           C1 => B(6), C2 => n177, ZN => n59);
   U117 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U118 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN
                           => n56_port);
   U119 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, 
                           C1 => B(7), C2 => n177, ZN => n57_port);
   U120 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U121 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN
                           => n54_port);
   U122 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, 
                           C1 => B(8), C2 => n176, ZN => n55_port);
   U123 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U124 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN
                           => n52_port);
   U125 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, 
                           C1 => B(9), C2 => n176, ZN => n53_port);
   U126 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U127 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U128 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180,
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U129 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U130 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U131 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180,
                           C1 => B(11), C2 => n176, ZN => n49_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_3 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_3;

architecture SYN_Behavioral of MUX5to1_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n187, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n188, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n189, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n188, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n188);
   U10 : BUF_X1 port map( A => n190, Z => n187);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U37 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U38 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180, 
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U39 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U40 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U41 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U42 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U43 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U44 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U45 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U46 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U47 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U48 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U49 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U50 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U51 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U52 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U53 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U54 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U55 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U56 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U57 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U58 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U59 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U60 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U61 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U62 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U63 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U64 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U65 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U66 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U67 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U68 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179, 
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U69 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U70 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U71 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179, 
                           C1 => B(24), C2 => n175, ZN => n23);
   U72 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U73 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U74 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U75 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U76 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U77 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U78 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U79 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179, 
                           C1 => B(25), C2 => n175, ZN => n21);
   U80 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U81 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U82 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U83 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179, 
                           C1 => B(26), C2 => n175, ZN => n19);
   U84 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U85 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U86 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180, 
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U87 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U88 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U89 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179, 
                           C1 => B(27), C2 => n175, ZN => n17);
   U90 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U91 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U92 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179, 
                           C1 => B(28), C2 => n175, ZN => n15);
   U93 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U94 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U95 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179, 
                           C1 => B(29), C2 => n175, ZN => n13);
   U96 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U97 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U98 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179, 
                           C1 => B(30), C2 => n175, ZN => n11);
   U99 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U100 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U101 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179,
                           C1 => B(31), C2 => n175, ZN => n4);
   U102 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U103 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN
                           => n70);
   U104 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, 
                           C1 => B(0), C2 => n177, ZN => n71);
   U105 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U106 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN
                           => n68);
   U107 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, 
                           C1 => B(1), C2 => n177, ZN => n69);
   U108 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U109 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN
                           => n66);
   U110 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, 
                           C1 => B(2), C2 => n177, ZN => n67);
   U111 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U112 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN
                           => n64);
   U113 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, 
                           C1 => B(3), C2 => n177, ZN => n65);
   U114 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U115 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN
                           => n62);
   U116 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, 
                           C1 => B(4), C2 => n177, ZN => n63);
   U117 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U118 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN
                           => n60);
   U119 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, 
                           C1 => B(5), C2 => n177, ZN => n61);
   U120 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U121 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN
                           => n58);
   U122 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, 
                           C1 => B(6), C2 => n177, ZN => n59);
   U123 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U124 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN
                           => n56_port);
   U125 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, 
                           C1 => B(7), C2 => n177, ZN => n57_port);
   U126 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U127 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN
                           => n54_port);
   U128 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, 
                           C1 => B(8), C2 => n176, ZN => n55_port);
   U129 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U130 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN
                           => n52_port);
   U131 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, 
                           C1 => B(9), C2 => n176, ZN => n53_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_4 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_4;

architecture SYN_Behavioral of MUX5to1_NBIT32_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n188, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n187, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n188, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n187);
   U10 : BUF_X1 port map( A => n190, Z => n188);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U37 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN 
                           => n52_port);
   U38 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, C1
                           => B(9), C2 => n176, ZN => n53_port);
   U39 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U40 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U41 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180, 
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U42 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U43 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U44 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180, 
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U45 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U46 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U47 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U48 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U49 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U50 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U51 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U52 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U53 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U54 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U55 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U56 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U57 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U58 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U59 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U60 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U61 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U62 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U63 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U64 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U65 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U66 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U67 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U68 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U69 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U70 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U71 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U72 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U73 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U74 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U75 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U76 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U77 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U78 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U79 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179, 
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U80 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U81 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U82 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U83 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179, 
                           C1 => B(24), C2 => n175, ZN => n23);
   U84 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U85 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN 
                           => n54_port);
   U86 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, C1
                           => B(8), C2 => n176, ZN => n55_port);
   U87 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U88 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U89 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179, 
                           C1 => B(25), C2 => n175, ZN => n21);
   U90 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U91 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U92 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179, 
                           C1 => B(26), C2 => n175, ZN => n19);
   U93 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U94 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U95 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179, 
                           C1 => B(27), C2 => n175, ZN => n17);
   U96 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U97 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U98 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179, 
                           C1 => B(28), C2 => n175, ZN => n15);
   U99 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U100 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U101 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179,
                           C1 => B(29), C2 => n175, ZN => n13);
   U102 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U103 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U104 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179,
                           C1 => B(30), C2 => n175, ZN => n11);
   U105 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U106 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U107 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179,
                           C1 => B(31), C2 => n175, ZN => n4);
   U108 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U109 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN
                           => n70);
   U110 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, 
                           C1 => B(0), C2 => n177, ZN => n71);
   U111 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U112 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN
                           => n68);
   U113 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, 
                           C1 => B(1), C2 => n177, ZN => n69);
   U114 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U115 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN
                           => n66);
   U116 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, 
                           C1 => B(2), C2 => n177, ZN => n67);
   U117 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U118 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN
                           => n64);
   U119 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, 
                           C1 => B(3), C2 => n177, ZN => n65);
   U120 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U121 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN
                           => n62);
   U122 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, 
                           C1 => B(4), C2 => n177, ZN => n63);
   U123 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U124 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN
                           => n60);
   U125 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, 
                           C1 => B(5), C2 => n177, ZN => n61);
   U126 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U127 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN
                           => n58);
   U128 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, 
                           C1 => B(6), C2 => n177, ZN => n59);
   U129 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U130 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN
                           => n56_port);
   U131 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, 
                           C1 => B(7), C2 => n177, ZN => n57_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_5 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_5;

architecture SYN_Behavioral of MUX5to1_NBIT32_5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n188, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n187, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n189, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n188, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n187);
   U10 : BUF_X1 port map( A => n190, Z => n188);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U37 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN 
                           => n56_port);
   U38 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, C1
                           => B(7), C2 => n177, ZN => n57_port);
   U39 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U40 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN 
                           => n54_port);
   U41 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, C1
                           => B(8), C2 => n176, ZN => n55_port);
   U42 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U43 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN 
                           => n52_port);
   U44 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, C1
                           => B(9), C2 => n176, ZN => n53_port);
   U45 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U46 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U47 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180, 
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U48 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U49 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U50 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U51 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U52 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U53 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U54 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U55 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U56 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U57 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U58 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U59 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U60 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U61 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U62 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U63 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U64 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U65 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U66 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U67 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U68 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U69 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U70 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U71 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U72 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U73 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180, 
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U74 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U75 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U76 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U77 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U78 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U79 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U80 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U81 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U82 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U83 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U84 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U85 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN 
                           => n58);
   U86 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, C1
                           => B(6), C2 => n177, ZN => n59);
   U87 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U88 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U89 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179, 
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U90 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U91 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U92 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179, 
                           C1 => B(24), C2 => n175, ZN => n23);
   U93 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U94 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U95 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179, 
                           C1 => B(25), C2 => n175, ZN => n21);
   U96 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U97 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U98 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179, 
                           C1 => B(26), C2 => n175, ZN => n19);
   U99 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U100 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U101 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179,
                           C1 => B(27), C2 => n175, ZN => n17);
   U102 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U103 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U104 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179,
                           C1 => B(28), C2 => n175, ZN => n15);
   U105 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U106 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U107 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179,
                           C1 => B(29), C2 => n175, ZN => n13);
   U108 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U109 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U110 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179,
                           C1 => B(30), C2 => n175, ZN => n11);
   U111 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U112 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U113 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179,
                           C1 => B(31), C2 => n175, ZN => n4);
   U114 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U115 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN
                           => n70);
   U116 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, 
                           C1 => B(0), C2 => n177, ZN => n71);
   U117 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U118 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN
                           => n68);
   U119 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, 
                           C1 => B(1), C2 => n177, ZN => n69);
   U120 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U121 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN
                           => n66);
   U122 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, 
                           C1 => B(2), C2 => n177, ZN => n67);
   U123 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U124 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN
                           => n64);
   U125 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, 
                           C1 => B(3), C2 => n177, ZN => n65);
   U126 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U127 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN
                           => n62);
   U128 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, 
                           C1 => B(4), C2 => n177, ZN => n63);
   U129 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U130 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN
                           => n60);
   U131 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, 
                           C1 => B(5), C2 => n177, ZN => n61);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_6 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_6;

architecture SYN_Behavioral of MUX5to1_NBIT32_6 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n187, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n188, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n189, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n188, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n188);
   U10 : BUF_X1 port map( A => n190, Z => n187);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U37 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN 
                           => n60);
   U38 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, C1
                           => B(5), C2 => n177, ZN => n61);
   U39 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U40 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN 
                           => n58);
   U41 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, C1
                           => B(6), C2 => n177, ZN => n59);
   U42 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U43 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN 
                           => n56_port);
   U44 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, C1
                           => B(7), C2 => n177, ZN => n57_port);
   U45 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U46 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN 
                           => n54_port);
   U47 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, C1
                           => B(8), C2 => n176, ZN => n55_port);
   U48 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U49 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U50 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180, 
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U51 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U52 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U53 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180, 
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U54 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U55 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U56 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U57 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U58 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U59 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U60 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U61 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U62 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U63 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U64 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U65 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U66 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U67 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U68 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U69 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U70 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U71 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U72 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U73 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, C1
                           => B(9), C2 => n176, ZN => n53_port);
   U74 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN 
                           => n52_port);
   U75 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U76 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U77 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U78 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U79 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U80 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U81 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U82 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U83 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U84 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U85 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN 
                           => n62);
   U86 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, C1
                           => B(4), C2 => n177, ZN => n63);
   U87 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U88 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U89 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U90 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U91 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U92 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U93 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U94 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U95 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179, 
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U96 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U97 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U98 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179, 
                           C1 => B(24), C2 => n175, ZN => n23);
   U99 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U100 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U101 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179,
                           C1 => B(25), C2 => n175, ZN => n21);
   U102 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U103 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U104 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179,
                           C1 => B(26), C2 => n175, ZN => n19);
   U105 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U106 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U107 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179,
                           C1 => B(27), C2 => n175, ZN => n17);
   U108 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U109 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U110 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179,
                           C1 => B(28), C2 => n175, ZN => n15);
   U111 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U112 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U113 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179,
                           C1 => B(29), C2 => n175, ZN => n13);
   U114 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U115 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U116 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179,
                           C1 => B(30), C2 => n175, ZN => n11);
   U117 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U118 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U119 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179,
                           C1 => B(31), C2 => n175, ZN => n4);
   U120 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U121 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN
                           => n70);
   U122 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, 
                           C1 => B(0), C2 => n177, ZN => n71);
   U123 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U124 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN
                           => n68);
   U125 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, 
                           C1 => B(1), C2 => n177, ZN => n69);
   U126 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U127 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN
                           => n66);
   U128 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, 
                           C1 => B(2), C2 => n177, ZN => n67);
   U129 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U130 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN
                           => n64);
   U131 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, 
                           C1 => B(3), C2 => n177, ZN => n65);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_7 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_7;

architecture SYN_Behavioral of MUX5to1_NBIT32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n187, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n188, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n189, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n188, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n189, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n188);
   U10 : BUF_X1 port map( A => n190, Z => n187);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n191);
   U30 : INV_X1 port map( A => SEL(0), ZN => n192);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n191, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n192, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n191, A2 => SEL(2), A3 => n192, ZN => n8);
   U35 : AND3_X1 port map( A1 => n192, A2 => n191, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U37 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN 
                           => n64);
   U38 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, C1
                           => B(3), C2 => n177, ZN => n65);
   U39 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U40 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN 
                           => n62);
   U41 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, C1
                           => B(4), C2 => n177, ZN => n63);
   U42 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U43 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN 
                           => n60);
   U44 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, C1
                           => B(5), C2 => n177, ZN => n61);
   U45 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U46 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN 
                           => n58);
   U47 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, C1
                           => B(6), C2 => n177, ZN => n59);
   U48 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U49 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN 
                           => n54_port);
   U50 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, C1
                           => B(8), C2 => n176, ZN => n55_port);
   U51 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U52 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN 
                           => n52_port);
   U53 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, C1
                           => B(9), C2 => n176, ZN => n53_port);
   U54 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U55 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U56 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180, 
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U57 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U58 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U59 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180, 
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U60 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U61 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U62 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U63 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U64 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U65 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U66 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U67 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U68 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U69 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U70 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U71 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U72 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U73 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, C1
                           => B(7), C2 => n177, ZN => n57_port);
   U74 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN 
                           => n56_port);
   U75 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U76 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U77 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U78 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U79 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U80 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U81 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U82 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U83 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U84 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U85 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN 
                           => n66);
   U86 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, C1
                           => B(2), C2 => n177, ZN => n67);
   U87 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U88 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U89 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U90 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U91 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U92 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U93 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U94 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U95 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179, 
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U96 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U97 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U98 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179, 
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U99 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U100 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U101 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179,
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U102 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U103 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U104 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179,
                           C1 => B(24), C2 => n175, ZN => n23);
   U105 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U106 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U107 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179,
                           C1 => B(25), C2 => n175, ZN => n21);
   U108 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U109 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U110 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179,
                           C1 => B(26), C2 => n175, ZN => n19);
   U111 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U112 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U113 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179,
                           C1 => B(27), C2 => n175, ZN => n17);
   U114 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U115 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U116 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179,
                           C1 => B(28), C2 => n175, ZN => n15);
   U117 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U118 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U119 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179,
                           C1 => B(29), C2 => n175, ZN => n13);
   U120 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U121 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U122 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179,
                           C1 => B(30), C2 => n175, ZN => n11);
   U123 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U124 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U125 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179,
                           C1 => B(31), C2 => n175, ZN => n4);
   U126 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U127 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN
                           => n70);
   U128 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, 
                           C1 => B(0), C2 => n177, ZN => n71);
   U129 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U130 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN
                           => n68);
   U131 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, 
                           C1 => B(1), C2 => n177, ZN => n69);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_8 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_8;

architecture SYN_Behavioral of MUX5to1_NBIT32_8 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n167, n168, n169, n170, n171, n172, n173,
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n187, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n188, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n188, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n188, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n188, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n188, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n188, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n188, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n188, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n188, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n188, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n189, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n189, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n189, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n189, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n189, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n189, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n189, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n189, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n188, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n189, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n189, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n187, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n187, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n187, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n187, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n187, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n187, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n187, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n187, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n187, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n187, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n190);
   U4 : BUF_X1 port map( A => n6, Z => n182);
   U5 : BUF_X1 port map( A => n7, Z => n178);
   U6 : BUF_X1 port map( A => n5, Z => n186);
   U7 : BUF_X1 port map( A => n8, Z => n174);
   U8 : BUF_X1 port map( A => n9, Z => n167);
   U9 : BUF_X1 port map( A => n190, Z => n188);
   U10 : BUF_X1 port map( A => n190, Z => n187);
   U11 : BUF_X1 port map( A => n190, Z => n189);
   U12 : OR4_X1 port map( A1 => n173, A2 => n170, A3 => n185, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n177, A2 => n181, ZN => n72);
   U14 : BUF_X1 port map( A => n174, Z => n172);
   U15 : BUF_X1 port map( A => n174, Z => n171);
   U16 : BUF_X1 port map( A => n182, Z => n180);
   U17 : BUF_X1 port map( A => n182, Z => n179);
   U18 : BUF_X1 port map( A => n167, Z => n169);
   U19 : BUF_X1 port map( A => n167, Z => n168);
   U20 : BUF_X1 port map( A => n178, Z => n176);
   U21 : BUF_X1 port map( A => n178, Z => n175);
   U22 : BUF_X1 port map( A => n186, Z => n184);
   U23 : BUF_X1 port map( A => n186, Z => n183);
   U24 : BUF_X1 port map( A => n174, Z => n173);
   U25 : BUF_X1 port map( A => n182, Z => n181);
   U26 : BUF_X1 port map( A => n167, Z => n170);
   U27 : BUF_X1 port map( A => n178, Z => n177);
   U28 : BUF_X1 port map( A => n186, Z => n185);
   U29 : INV_X1 port map( A => SEL(1), ZN => n192);
   U30 : INV_X1 port map( A => SEL(0), ZN => n191);
   U31 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n192, ZN => n6);
   U32 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n191, ZN => n7);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U34 : NOR3_X1 port map( A1 => n192, A2 => SEL(2), A3 => n191, ZN => n8);
   U35 : AND3_X1 port map( A1 => n191, A2 => n192, A3 => SEL(2), ZN => n9);
   U36 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U37 : AOI22_X1 port map( A1 => D(1), A2 => n173, B1 => E(1), B2 => n170, ZN 
                           => n68);
   U38 : AOI222_X1 port map( A1 => A(1), A2 => n185, B1 => C(1), B2 => n181, C1
                           => B(1), C2 => n177, ZN => n69);
   U39 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U40 : AOI22_X1 port map( A1 => D(2), A2 => n173, B1 => E(2), B2 => n170, ZN 
                           => n66);
   U41 : AOI222_X1 port map( A1 => A(2), A2 => n185, B1 => C(2), B2 => n181, C1
                           => B(2), C2 => n177, ZN => n67);
   U42 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U43 : AOI22_X1 port map( A1 => D(3), A2 => n173, B1 => E(3), B2 => n170, ZN 
                           => n64);
   U44 : AOI222_X1 port map( A1 => A(3), A2 => n185, B1 => C(3), B2 => n181, C1
                           => B(3), C2 => n177, ZN => n65);
   U45 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U46 : AOI22_X1 port map( A1 => D(4), A2 => n173, B1 => E(4), B2 => n170, ZN 
                           => n62);
   U47 : AOI222_X1 port map( A1 => A(4), A2 => n185, B1 => C(4), B2 => n181, C1
                           => B(4), C2 => n177, ZN => n63);
   U48 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U49 : AOI22_X1 port map( A1 => D(6), A2 => n173, B1 => E(6), B2 => n170, ZN 
                           => n58);
   U50 : AOI222_X1 port map( A1 => A(6), A2 => n185, B1 => C(6), B2 => n181, C1
                           => B(6), C2 => n177, ZN => n59);
   U51 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U52 : AOI22_X1 port map( A1 => D(7), A2 => n173, B1 => E(7), B2 => n170, ZN 
                           => n56_port);
   U53 : AOI222_X1 port map( A1 => A(7), A2 => n185, B1 => C(7), B2 => n181, C1
                           => B(7), C2 => n177, ZN => n57_port);
   U54 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U55 : AOI22_X1 port map( A1 => D(8), A2 => n172, B1 => E(8), B2 => n169, ZN 
                           => n54_port);
   U56 : AOI222_X1 port map( A1 => A(8), A2 => n184, B1 => C(8), B2 => n180, C1
                           => B(8), C2 => n176, ZN => n55_port);
   U57 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U58 : AOI22_X1 port map( A1 => D(9), A2 => n172, B1 => E(9), B2 => n169, ZN 
                           => n52_port);
   U59 : AOI222_X1 port map( A1 => A(9), A2 => n184, B1 => C(9), B2 => n180, C1
                           => B(9), C2 => n176, ZN => n53_port);
   U60 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U61 : AOI22_X1 port map( A1 => D(11), A2 => n172, B1 => E(11), B2 => n169, 
                           ZN => n48_port);
   U62 : AOI222_X1 port map( A1 => A(11), A2 => n184, B1 => C(11), B2 => n180, 
                           C1 => B(11), C2 => n176, ZN => n49_port);
   U63 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U64 : AOI22_X1 port map( A1 => D(12), A2 => n172, B1 => E(12), B2 => n169, 
                           ZN => n46_port);
   U65 : AOI222_X1 port map( A1 => A(12), A2 => n184, B1 => C(12), B2 => n180, 
                           C1 => B(12), C2 => n176, ZN => n47_port);
   U66 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U67 : AOI22_X1 port map( A1 => D(13), A2 => n172, B1 => E(13), B2 => n169, 
                           ZN => n44_port);
   U68 : AOI222_X1 port map( A1 => A(13), A2 => n184, B1 => C(13), B2 => n180, 
                           C1 => B(13), C2 => n176, ZN => n45_port);
   U69 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U70 : AOI22_X1 port map( A1 => D(14), A2 => n172, B1 => E(14), B2 => n169, 
                           ZN => n42_port);
   U71 : AOI222_X1 port map( A1 => A(14), A2 => n184, B1 => C(14), B2 => n180, 
                           C1 => B(14), C2 => n176, ZN => n43_port);
   U72 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U73 : AOI222_X1 port map( A1 => A(5), A2 => n185, B1 => C(5), B2 => n181, C1
                           => B(5), C2 => n177, ZN => n61);
   U74 : AOI22_X1 port map( A1 => D(5), A2 => n173, B1 => E(5), B2 => n170, ZN 
                           => n60);
   U75 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U76 : AOI222_X1 port map( A1 => A(10), A2 => n184, B1 => C(10), B2 => n180, 
                           C1 => B(10), C2 => n176, ZN => n51_port);
   U77 : AOI22_X1 port map( A1 => D(10), A2 => n172, B1 => E(10), B2 => n169, 
                           ZN => n50_port);
   U78 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U79 : AOI222_X1 port map( A1 => A(15), A2 => n184, B1 => C(15), B2 => n180, 
                           C1 => B(15), C2 => n176, ZN => n41_port);
   U80 : AOI22_X1 port map( A1 => D(15), A2 => n172, B1 => E(15), B2 => n169, 
                           ZN => n40_port);
   U81 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U82 : AOI22_X1 port map( A1 => D(16), A2 => n172, B1 => E(16), B2 => n169, 
                           ZN => n38_port);
   U83 : AOI222_X1 port map( A1 => A(16), A2 => n184, B1 => C(16), B2 => n180, 
                           C1 => B(16), C2 => n176, ZN => n39_port);
   U84 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U85 : AOI22_X1 port map( A1 => D(0), A2 => n173, B1 => E(0), B2 => n170, ZN 
                           => n70);
   U86 : AOI222_X1 port map( A1 => A(0), A2 => n185, B1 => C(0), B2 => n181, C1
                           => B(0), C2 => n177, ZN => n71);
   U87 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U88 : AOI22_X1 port map( A1 => D(17), A2 => n172, B1 => E(17), B2 => n169, 
                           ZN => n36_port);
   U89 : AOI222_X1 port map( A1 => A(17), A2 => n184, B1 => C(17), B2 => n180, 
                           C1 => B(17), C2 => n176, ZN => n37_port);
   U90 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U91 : AOI22_X1 port map( A1 => D(18), A2 => n172, B1 => E(18), B2 => n169, 
                           ZN => n34_port);
   U92 : AOI222_X1 port map( A1 => A(18), A2 => n184, B1 => C(18), B2 => n180, 
                           C1 => B(18), C2 => n176, ZN => n35_port);
   U93 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U94 : AOI22_X1 port map( A1 => D(19), A2 => n172, B1 => E(19), B2 => n169, 
                           ZN => n32_port);
   U95 : AOI222_X1 port map( A1 => A(19), A2 => n184, B1 => C(19), B2 => n180, 
                           C1 => B(19), C2 => n176, ZN => n33_port);
   U96 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U97 : AOI22_X1 port map( A1 => D(20), A2 => n171, B1 => E(20), B2 => n168, 
                           ZN => n30_port);
   U98 : AOI222_X1 port map( A1 => A(20), A2 => n183, B1 => C(20), B2 => n179, 
                           C1 => B(20), C2 => n175, ZN => n31_port);
   U99 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U100 : AOI22_X1 port map( A1 => D(21), A2 => n171, B1 => E(21), B2 => n168, 
                           ZN => n28_port);
   U101 : AOI222_X1 port map( A1 => A(21), A2 => n183, B1 => C(21), B2 => n179,
                           C1 => B(21), C2 => n175, ZN => n29_port);
   U102 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U103 : AOI22_X1 port map( A1 => D(22), A2 => n171, B1 => E(22), B2 => n168, 
                           ZN => n26_port);
   U104 : AOI222_X1 port map( A1 => A(22), A2 => n183, B1 => C(22), B2 => n179,
                           C1 => B(22), C2 => n175, ZN => n27_port);
   U105 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U106 : AOI22_X1 port map( A1 => D(23), A2 => n171, B1 => E(23), B2 => n168, 
                           ZN => n24);
   U107 : AOI222_X1 port map( A1 => A(23), A2 => n183, B1 => C(23), B2 => n179,
                           C1 => B(23), C2 => n175, ZN => n25_port);
   U108 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U109 : AOI22_X1 port map( A1 => D(24), A2 => n171, B1 => E(24), B2 => n168, 
                           ZN => n22);
   U110 : AOI222_X1 port map( A1 => A(24), A2 => n183, B1 => C(24), B2 => n179,
                           C1 => B(24), C2 => n175, ZN => n23);
   U111 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U112 : AOI22_X1 port map( A1 => D(25), A2 => n171, B1 => E(25), B2 => n168, 
                           ZN => n20);
   U113 : AOI222_X1 port map( A1 => A(25), A2 => n183, B1 => C(25), B2 => n179,
                           C1 => B(25), C2 => n175, ZN => n21);
   U114 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U115 : AOI22_X1 port map( A1 => D(26), A2 => n171, B1 => E(26), B2 => n168, 
                           ZN => n18);
   U116 : AOI222_X1 port map( A1 => A(26), A2 => n183, B1 => C(26), B2 => n179,
                           C1 => B(26), C2 => n175, ZN => n19);
   U117 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U118 : AOI22_X1 port map( A1 => D(27), A2 => n171, B1 => E(27), B2 => n168, 
                           ZN => n16);
   U119 : AOI222_X1 port map( A1 => A(27), A2 => n183, B1 => C(27), B2 => n179,
                           C1 => B(27), C2 => n175, ZN => n17);
   U120 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U121 : AOI22_X1 port map( A1 => D(28), A2 => n171, B1 => E(28), B2 => n168, 
                           ZN => n14);
   U122 : AOI222_X1 port map( A1 => A(28), A2 => n183, B1 => C(28), B2 => n179,
                           C1 => B(28), C2 => n175, ZN => n15);
   U123 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U124 : AOI22_X1 port map( A1 => D(29), A2 => n171, B1 => E(29), B2 => n168, 
                           ZN => n12);
   U125 : AOI222_X1 port map( A1 => A(29), A2 => n183, B1 => C(29), B2 => n179,
                           C1 => B(29), C2 => n175, ZN => n13);
   U126 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U127 : AOI22_X1 port map( A1 => D(30), A2 => n171, B1 => E(30), B2 => n168, 
                           ZN => n10);
   U128 : AOI222_X1 port map( A1 => A(30), A2 => n183, B1 => C(30), B2 => n179,
                           C1 => B(30), C2 => n175, ZN => n11);
   U129 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U130 : AOI22_X1 port map( A1 => D(31), A2 => n171, B1 => E(31), B2 => n168, 
                           ZN => n3);
   U131 : AOI222_X1 port map( A1 => A(31), A2 => n183, B1 => C(31), B2 => n179,
                           C1 => B(31), C2 => n175, ZN => n4);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_7 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_7;

architecture SYN_BEHAVIORAL of ENCODER_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n9 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n3, A2 => n9, B1 => INPUT(2), B2 => n2, ZN => 
                           OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n9);
   U3 : AOI21_X1 port map( B1 => n3, B2 => n2, A => INPUT(2), ZN => OUTPUT(0));
   U4 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n3);
   U5 : AND3_X1 port map( A1 => INPUT(2), A2 => n2, A3 => n3, ZN => OUTPUT(2));
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_0 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_0;

architecture SYN_BEHAVIORAL of ENCODER_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => INPUT(2), B2 => n2, ZN => 
                           OUTPUT(1));
   U2 : INV_X1 port map( A => INPUT(2), ZN => n4);
   U3 : AOI21_X1 port map( B1 => n3, B2 => n2, A => INPUT(2), ZN => OUTPUT(0));
   U4 : AND3_X1 port map( A1 => INPUT(2), A2 => n2, A3 => n3, ZN => OUTPUT(2));
   U5 : XNOR2_X1 port map( A => INPUT(0), B => INPUT(1), ZN => n3);
   U6 : NAND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_0 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_0;

architecture SYN_ARCH1 of ND4_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_0 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_0;

architecture SYN_ARCH1 of ND3_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 is

   component CARRY_SEL_N_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_63 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_62 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_61 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_60 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_59 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_58 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_57 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_64
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_65
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_66
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_67
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_190
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_191
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_68
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_69
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_192
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_193
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_194
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_70
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_195
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_196
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_197
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_198
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_199
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_200
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_201
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_71
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_202
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_203
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_204
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_205
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_206
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_207
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_208
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_209
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_210
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_211
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_212
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_213
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_214
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_215
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_0
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_0
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n3, n4, n5, n6, n7, n_1135 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_0 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1135, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n3);
   gblock1_1_1 : G_block_0 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B 
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_0 port map( A(1) => P_4_4_port, A(0) => G_4_4_port, 
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_215 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_214 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_213 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_212 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_211 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_210 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_209 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_208 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_207 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_206 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_205 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_204 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_203 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_202 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_71 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_201 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_200 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_199 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_198 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_197 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_196 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_195 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_70 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_194 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_193 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_192 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_69 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_68 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_191 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_190 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_67 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_66 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_65 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_64 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NOR2_X1 port map( A1 => n6, A2 => n4, ZN => G_1_0_port);
   U2 : INV_X1 port map( A => n3, ZN => n6);
   U3 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n7, ZN => n4);
   U4 : INV_X1 port map( A => n5, ZN => n7);
   U5 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n5);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1;

architecture SYN_rpl of HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n6, n7, n9, n11, n12, n15, n16, n17, n18, n20, n21, n22, n23,
      n25, n26, n27, n28, n30, n32, n33, n34, n35, n73, n74, n75, n76, n77, n78
      , n79, n80, n82, n83, n84, n85, n86, n87, n89, n91, n92, n94, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n111, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n86, ZN => n127);
   U2 : INV_X1 port map( A => n7, ZN => n124);
   U3 : INV_X1 port map( A => n4, ZN => n122);
   U4 : INV_X1 port map( A => n2, ZN => n119);
   U5 : INV_X1 port map( A => n9, ZN => n117);
   U6 : NAND2_X1 port map( A1 => n96, A2 => n146, ZN => n9);
   U7 : NAND2_X1 port map( A1 => n94, A2 => n144, ZN => n2);
   U8 : NAND2_X1 port map( A1 => n91, A2 => n141, ZN => n4);
   U9 : NAND2_X1 port map( A1 => n89, A2 => n139, ZN => n7);
   U10 : NAND2_X1 port map( A1 => n84, A2 => n135, ZN => n82);
   U11 : AND2_X1 port map( A1 => n87, A2 => n137, ZN => n86);
   U12 : AND2_X1 port map( A1 => n92, A2 => n142, ZN => n91);
   U13 : INV_X1 port map( A => n98, ZN => n128);
   U14 : INV_X1 port map( A => n80, ZN => n130);
   U15 : INV_X1 port map( A => n79, ZN => n129);
   U16 : AND2_X1 port map( A1 => n153, A2 => n28, ZN => n26);
   U17 : AND2_X1 port map( A1 => n151, A2 => n23, ZN => n21);
   U18 : INV_X1 port map( A => n87, ZN => n125);
   U19 : INV_X1 port map( A => n89, ZN => n123);
   U20 : INV_X1 port map( A => n92, ZN => n120);
   U21 : INV_X1 port map( A => n94, ZN => n118);
   U22 : INV_X1 port map( A => n96, ZN => n116);
   U23 : INV_X1 port map( A => n78, ZN => n115);
   U24 : INV_X1 port map( A => n105, ZN => n111);
   U25 : AND2_X1 port map( A1 => n17, A2 => n18, ZN => n99);
   U26 : AND2_X1 port map( A1 => n78, A2 => n157, ZN => n17);
   U27 : INV_X1 port map( A => n35, ZN => n109);
   U28 : INV_X1 port map( A => n34, ZN => n108);
   U29 : OAI21_X1 port map( B1 => n117, B2 => n145, A => n118, ZN => SUM(18));
   U30 : INV_X1 port map( A => A(18), ZN => n145);
   U31 : OAI21_X1 port map( B1 => n91, B2 => n141, A => n4, ZN => SUM(22));
   U32 : INV_X1 port map( A => n73, ZN => SUM(9));
   U33 : AOI21_X1 port map( B1 => n74, B2 => A(9), A => n75, ZN => n73);
   U34 : INV_X1 port map( A => n100, ZN => SUM(13));
   U35 : AOI21_X1 port map( B1 => n101, B2 => A(13), A => n99, ZN => n100);
   U36 : OAI21_X1 port map( B1 => n96, B2 => n146, A => n9, ZN => SUM(17));
   U37 : OAI21_X1 port map( B1 => n84, B2 => n135, A => n82, ZN => SUM(29));
   U38 : OAI21_X1 port map( B1 => n76, B2 => n155, A => n74, ZN => SUM(8));
   U39 : INV_X1 port map( A => A(8), ZN => n155);
   U40 : OAI21_X1 port map( B1 => n102, B2 => n151, A => n101, ZN => SUM(12));
   U41 : OAI21_X1 port map( B1 => n97, B2 => n147, A => n116, ZN => SUM(16));
   U42 : INV_X1 port map( A => A(16), ZN => n147);
   U43 : INV_X1 port map( A => n85, ZN => SUM(28));
   U44 : AOI21_X1 port map( B1 => n33, B2 => A(28), A => n84, ZN => n85);
   U45 : OAI21_X1 port map( B1 => n94, B2 => n144, A => n2, ZN => SUM(19));
   U46 : OAI21_X1 port map( B1 => n122, B2 => n140, A => n123, ZN => SUM(23));
   U47 : INV_X1 port map( A => A(23), ZN => n140);
   U48 : INV_X1 port map( A => n77, ZN => SUM(7));
   U49 : AOI21_X1 port map( B1 => n111, B2 => A(7), A => n76, ZN => n77);
   U50 : INV_X1 port map( A => n103, ZN => SUM(11));
   U51 : AOI21_X1 port map( B1 => n104, B2 => A(11), A => n102, ZN => n103);
   U52 : OAI21_X1 port map( B1 => n98, B2 => n148, A => n11, ZN => SUM(15));
   U53 : INV_X1 port map( A => A(15), ZN => n148);
   U54 : OAI21_X1 port map( B1 => n86, B2 => n136, A => n33, ZN => SUM(27));
   U55 : OAI21_X1 port map( B1 => n75, B2 => n153, A => n104, ZN => SUM(10));
   U56 : OAI21_X1 port map( B1 => n99, B2 => n149, A => n128, ZN => SUM(14));
   U57 : INV_X1 port map( A => A(14), ZN => n149);
   U58 : OAI21_X1 port map( B1 => n119, B2 => n143, A => n120, ZN => SUM(20));
   U59 : INV_X1 port map( A => A(20), ZN => n143);
   U60 : OAI21_X1 port map( B1 => n92, B2 => n142, A => n121, ZN => SUM(21));
   U61 : INV_X1 port map( A => n91, ZN => n121);
   U62 : OAI21_X1 port map( B1 => n89, B2 => n139, A => n7, ZN => SUM(24));
   U63 : OAI21_X1 port map( B1 => n124, B2 => n138, A => n125, ZN => SUM(25));
   U64 : INV_X1 port map( A => A(25), ZN => n138);
   U65 : OAI21_X1 port map( B1 => n87, B2 => n137, A => n127, ZN => SUM(26));
   U66 : XNOR2_X1 port map( A => A(30), B => n82, ZN => SUM(30));
   U67 : OAI21_X1 port map( B1 => n79, B2 => n131, A => n115, ZN => SUM(5));
   U68 : INV_X1 port map( A => A(5), ZN => n131);
   U69 : OAI21_X1 port map( B1 => n80, B2 => n132, A => n129, ZN => SUM(4));
   U70 : INV_X1 port map( A => A(4), ZN => n132);
   U71 : OAI21_X1 port map( B1 => n109, B2 => n133, A => n130, ZN => SUM(3));
   U72 : INV_X1 port map( A => A(3), ZN => n133);
   U73 : OAI21_X1 port map( B1 => n78, B2 => n157, A => n111, ZN => SUM(6));
   U74 : OAI21_X1 port map( B1 => n34, B2 => n134, A => n35, ZN => SUM(2));
   U75 : NOR2_X1 port map( A1 => n129, A2 => A(5), ZN => n78);
   U76 : NOR2_X1 port map( A1 => n11, A2 => A(16), ZN => n96);
   U77 : NOR2_X1 port map( A1 => n9, A2 => A(18), ZN => n94);
   U78 : NOR2_X1 port map( A1 => n4, A2 => A(23), ZN => n89);
   U79 : NOR2_X1 port map( A1 => n32, A2 => A(28), ZN => n84);
   U80 : NAND2_X1 port map( A1 => n86, A2 => n136, ZN => n32);
   U81 : NOR2_X1 port map( A1 => n7, A2 => A(25), ZN => n87);
   U82 : NOR2_X1 port map( A1 => n2, A2 => A(20), ZN => n92);
   U83 : XNOR2_X1 port map( A => A(31), B => n12, ZN => SUM(31));
   U84 : OR2_X1 port map( A1 => A(30), A2 => n82, ZN => n12);
   U85 : NOR2_X1 port map( A1 => n16, A2 => A(14), ZN => n98);
   U86 : NAND2_X1 port map( A1 => n15, A2 => n78, ZN => n16);
   U87 : AND2_X1 port map( A1 => n18, A2 => n157, ZN => n15);
   U88 : NOR2_X1 port map( A1 => n35, A2 => A(3), ZN => n80);
   U89 : NOR2_X1 port map( A1 => n130, A2 => A(4), ZN => n79);
   U90 : NAND2_X1 port map( A1 => n83, A2 => n134, ZN => n35);
   U91 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n83);
   U92 : OR2_X1 port map( A1 => n128, A2 => A(15), ZN => n11);
   U93 : INV_X1 port map( A => A(2), ZN => n134);
   U94 : NOR2_X1 port map( A1 => A(9), A2 => n106, ZN => n28);
   U95 : OR2_X1 port map( A1 => A(8), A2 => A(7), ZN => n106);
   U96 : AND2_X1 port map( A1 => n152, A2 => n26, ZN => n23);
   U97 : INV_X1 port map( A => A(11), ZN => n152);
   U98 : AND2_X1 port map( A1 => n150, A2 => n21, ZN => n18);
   U99 : INV_X1 port map( A => A(13), ZN => n150);
   U100 : INV_X1 port map( A => A(10), ZN => n153);
   U101 : OR2_X1 port map( A1 => n127, A2 => A(27), ZN => n33);
   U102 : INV_X1 port map( A => A(12), ZN => n151);
   U103 : INV_X1 port map( A => A(6), ZN => n157);
   U104 : OAI21_X1 port map( B1 => n154, B2 => n107, A => n108, ZN => SUM(1));
   U105 : INV_X1 port map( A => A(0), ZN => n154);
   U106 : INV_X1 port map( A => A(17), ZN => n146);
   U107 : INV_X1 port map( A => A(19), ZN => n144);
   U108 : INV_X1 port map( A => A(21), ZN => n142);
   U109 : INV_X1 port map( A => A(22), ZN => n141);
   U110 : NOR2_X1 port map( A1 => n115, A2 => A(6), ZN => n105);
   U111 : AND2_X1 port map( A1 => n105, A2 => n156, ZN => n76);
   U112 : INV_X1 port map( A => A(7), ZN => n156);
   U113 : NAND2_X1 port map( A1 => n30, A2 => n6, ZN => n74);
   U114 : NOR2_X1 port map( A1 => A(8), A2 => A(7), ZN => n6);
   U115 : NOR2_X1 port map( A1 => n115, A2 => A(6), ZN => n30);
   U116 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n104);
   U117 : NOR2_X1 port map( A1 => n115, A2 => A(6), ZN => n25);
   U118 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n101);
   U119 : NOR2_X1 port map( A1 => n115, A2 => A(6), ZN => n20);
   U120 : AND2_X1 port map( A1 => n27, A2 => n28, ZN => n75);
   U121 : NOR2_X1 port map( A1 => n115, A2 => A(6), ZN => n27);
   U122 : AND2_X1 port map( A1 => n22, A2 => n23, ZN => n102);
   U123 : NOR2_X1 port map( A1 => n115, A2 => A(6), ZN => n22);
   U124 : NOR2_X1 port map( A1 => n128, A2 => A(15), ZN => n97);
   U125 : INV_X1 port map( A => A(24), ZN => n139);
   U126 : INV_X1 port map( A => A(26), ZN => n137);
   U127 : INV_X1 port map( A => A(27), ZN => n136);
   U128 : INV_X1 port map( A => A(29), ZN => n135);
   U129 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n34);
   U130 : INV_X1 port map( A => A(1), ZN => n107);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX4to1_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX4to1_NBIT32_1;

architecture SYN_Behavioral of MUX4to1_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n157);
   U2 : BUF_X1 port map( A => n7, Z => n153);
   U3 : BUF_X1 port map( A => n4, Z => n162);
   U4 : BUF_X1 port map( A => n5, Z => n158);
   U5 : BUF_X1 port map( A => n157, Z => n154);
   U6 : BUF_X1 port map( A => n157, Z => n155);
   U7 : BUF_X1 port map( A => n162, Z => n163);
   U8 : BUF_X1 port map( A => n162, Z => n164);
   U9 : BUF_X1 port map( A => n153, Z => n150);
   U10 : BUF_X1 port map( A => n153, Z => n151);
   U11 : BUF_X1 port map( A => n158, Z => n159);
   U12 : BUF_X1 port map( A => n158, Z => n160);
   U13 : BUF_X1 port map( A => n157, Z => n156);
   U14 : BUF_X1 port map( A => n162, Z => n165);
   U15 : BUF_X1 port map( A => n153, Z => n152);
   U16 : BUF_X1 port map( A => n158, Z => n161);
   U17 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n6);
   U18 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n7);
   U19 : INV_X1 port map( A => SEL(0), ZN => n166);
   U20 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n4);
   U21 : AND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n5);
   U22 : AOI22_X1 port map( A1 => C(5), A2 => n165, B1 => D(5), B2 => n161, ZN 
                           => n15);
   U23 : AOI22_X1 port map( A1 => C(6), A2 => n165, B1 => D(6), B2 => n161, ZN 
                           => n13);
   U24 : AOI22_X1 port map( A1 => C(7), A2 => n165, B1 => D(7), B2 => n161, ZN 
                           => n11);
   U25 : AOI22_X1 port map( A1 => C(9), A2 => n165, B1 => D(9), B2 => n161, ZN 
                           => n3);
   U26 : AOI22_X1 port map( A1 => C(10), A2 => n163, B1 => D(10), B2 => n159, 
                           ZN => n67);
   U27 : AOI22_X1 port map( A1 => C(11), A2 => n163, B1 => D(11), B2 => n159, 
                           ZN => n65);
   U28 : AOI22_X1 port map( A1 => C(13), A2 => n163, B1 => D(13), B2 => n159, 
                           ZN => n61);
   U29 : AOI22_X1 port map( A1 => C(14), A2 => n163, B1 => D(14), B2 => n159, 
                           ZN => n59);
   U30 : AOI22_X1 port map( A1 => C(15), A2 => n163, B1 => D(15), B2 => n159, 
                           ZN => n57);
   U31 : AOI22_X1 port map( A1 => C(17), A2 => n163, B1 => D(17), B2 => n159, 
                           ZN => n53);
   U32 : AOI22_X1 port map( A1 => C(18), A2 => n163, B1 => D(18), B2 => n159, 
                           ZN => n51);
   U33 : AOI22_X1 port map( A1 => C(19), A2 => n163, B1 => D(19), B2 => n159, 
                           ZN => n49);
   U34 : AOI22_X1 port map( A1 => C(21), A2 => n164, B1 => D(21), B2 => n160, 
                           ZN => n43);
   U35 : AOI22_X1 port map( A1 => C(22), A2 => n164, B1 => D(22), B2 => n160, 
                           ZN => n41);
   U36 : AOI22_X1 port map( A1 => C(23), A2 => n164, B1 => D(23), B2 => n160, 
                           ZN => n39);
   U37 : AOI22_X1 port map( A1 => C(25), A2 => n164, B1 => D(25), B2 => n160, 
                           ZN => n35);
   U38 : AOI22_X1 port map( A1 => C(26), A2 => n164, B1 => D(26), B2 => n160, 
                           ZN => n33);
   U39 : AOI22_X1 port map( A1 => C(27), A2 => n164, B1 => D(27), B2 => n160, 
                           ZN => n31);
   U40 : AOI22_X1 port map( A1 => C(29), A2 => n164, B1 => D(29), B2 => n160, 
                           ZN => n27);
   U41 : AOI22_X1 port map( A1 => C(30), A2 => n164, B1 => D(30), B2 => n160, 
                           ZN => n23);
   U42 : AOI22_X1 port map( A1 => C(31), A2 => n165, B1 => D(31), B2 => n161, 
                           ZN => n21);
   U43 : AOI22_X1 port map( A1 => C(16), A2 => n163, B1 => D(16), B2 => n159, 
                           ZN => n55);
   U44 : AOI22_X1 port map( A1 => C(0), A2 => n163, B1 => D(0), B2 => n159, ZN 
                           => n69);
   U45 : AOI22_X1 port map( A1 => C(1), A2 => n163, B1 => D(1), B2 => n159, ZN 
                           => n47);
   U46 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => D(2), B2 => n160, ZN 
                           => n25);
   U47 : AOI22_X1 port map( A1 => C(3), A2 => n165, B1 => D(3), B2 => n161, ZN 
                           => n19);
   U48 : AOI22_X1 port map( A1 => C(4), A2 => n165, B1 => D(4), B2 => n161, ZN 
                           => n17);
   U49 : AOI22_X1 port map( A1 => C(8), A2 => n165, B1 => D(8), B2 => n161, ZN 
                           => n9);
   U50 : AOI22_X1 port map( A1 => C(12), A2 => n163, B1 => D(12), B2 => n159, 
                           ZN => n63);
   U51 : AOI22_X1 port map( A1 => C(20), A2 => n164, B1 => D(20), B2 => n160, 
                           ZN => n45);
   U52 : AOI22_X1 port map( A1 => C(24), A2 => n164, B1 => D(24), B2 => n160, 
                           ZN => n37);
   U53 : AOI22_X1 port map( A1 => C(28), A2 => n164, B1 => D(28), B2 => n160, 
                           ZN => n29);
   U54 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(16));
   U55 : AOI22_X1 port map( A1 => A(16), A2 => n154, B1 => B(16), B2 => n150, 
                           ZN => n54);
   U56 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(0));
   U57 : AOI22_X1 port map( A1 => A(0), A2 => n154, B1 => B(0), B2 => n150, ZN 
                           => n68);
   U58 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(1));
   U59 : AOI22_X1 port map( A1 => A(1), A2 => n154, B1 => B(1), B2 => n150, ZN 
                           => n46);
   U60 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(2));
   U61 : AOI22_X1 port map( A1 => A(2), A2 => n155, B1 => B(2), B2 => n151, ZN 
                           => n24);
   U62 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(3));
   U63 : AOI22_X1 port map( A1 => A(3), A2 => n156, B1 => B(3), B2 => n152, ZN 
                           => n18);
   U64 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(4));
   U65 : AOI22_X1 port map( A1 => A(4), A2 => n156, B1 => B(4), B2 => n152, ZN 
                           => n16);
   U66 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(5));
   U67 : AOI22_X1 port map( A1 => A(5), A2 => n156, B1 => B(5), B2 => n152, ZN 
                           => n14);
   U68 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(6));
   U69 : AOI22_X1 port map( A1 => A(6), A2 => n156, B1 => B(6), B2 => n152, ZN 
                           => n12);
   U70 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(7));
   U71 : AOI22_X1 port map( A1 => A(7), A2 => n156, B1 => B(7), B2 => n152, ZN 
                           => n10);
   U72 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(8));
   U73 : AOI22_X1 port map( A1 => A(8), A2 => n156, B1 => B(8), B2 => n152, ZN 
                           => n8);
   U74 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(9));
   U75 : AOI22_X1 port map( A1 => A(9), A2 => n156, B1 => B(9), B2 => n152, ZN 
                           => n2);
   U76 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(10));
   U77 : AOI22_X1 port map( A1 => A(10), A2 => n154, B1 => B(10), B2 => n150, 
                           ZN => n66);
   U78 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(11));
   U79 : AOI22_X1 port map( A1 => A(11), A2 => n154, B1 => B(11), B2 => n150, 
                           ZN => n64);
   U80 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(12));
   U81 : AOI22_X1 port map( A1 => A(12), A2 => n154, B1 => B(12), B2 => n150, 
                           ZN => n62);
   U82 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(13));
   U83 : AOI22_X1 port map( A1 => A(13), A2 => n154, B1 => B(13), B2 => n150, 
                           ZN => n60);
   U84 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(14));
   U85 : AOI22_X1 port map( A1 => A(14), A2 => n154, B1 => B(14), B2 => n150, 
                           ZN => n58);
   U86 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(15));
   U87 : AOI22_X1 port map( A1 => A(15), A2 => n154, B1 => B(15), B2 => n150, 
                           ZN => n56);
   U88 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(17));
   U89 : AOI22_X1 port map( A1 => A(17), A2 => n154, B1 => B(17), B2 => n150, 
                           ZN => n52);
   U90 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(18));
   U91 : AOI22_X1 port map( A1 => A(18), A2 => n154, B1 => B(18), B2 => n150, 
                           ZN => n50);
   U92 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(19));
   U93 : AOI22_X1 port map( A1 => A(19), A2 => n154, B1 => B(19), B2 => n150, 
                           ZN => n48);
   U94 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(20));
   U95 : AOI22_X1 port map( A1 => A(20), A2 => n155, B1 => B(20), B2 => n151, 
                           ZN => n44);
   U96 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(21));
   U97 : AOI22_X1 port map( A1 => A(21), A2 => n155, B1 => B(21), B2 => n151, 
                           ZN => n42);
   U98 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(22));
   U99 : AOI22_X1 port map( A1 => A(22), A2 => n155, B1 => B(22), B2 => n151, 
                           ZN => n40);
   U100 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(23));
   U101 : AOI22_X1 port map( A1 => A(23), A2 => n155, B1 => B(23), B2 => n151, 
                           ZN => n38);
   U102 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(24));
   U103 : AOI22_X1 port map( A1 => A(24), A2 => n155, B1 => B(24), B2 => n151, 
                           ZN => n36);
   U104 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(25));
   U105 : AOI22_X1 port map( A1 => A(25), A2 => n155, B1 => B(25), B2 => n151, 
                           ZN => n34);
   U106 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(26));
   U107 : AOI22_X1 port map( A1 => A(26), A2 => n155, B1 => B(26), B2 => n151, 
                           ZN => n32);
   U108 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(27));
   U109 : AOI22_X1 port map( A1 => A(27), A2 => n155, B1 => B(27), B2 => n151, 
                           ZN => n30);
   U110 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(28));
   U111 : AOI22_X1 port map( A1 => A(28), A2 => n155, B1 => B(28), B2 => n151, 
                           ZN => n28);
   U112 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(29));
   U113 : AOI22_X1 port map( A1 => A(29), A2 => n155, B1 => B(29), B2 => n151, 
                           ZN => n26);
   U114 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(30));
   U115 : AOI22_X1 port map( A1 => A(30), A2 => n155, B1 => B(30), B2 => n151, 
                           ZN => n22);
   U116 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(31));
   U117 : AOI22_X1 port map( A1 => A(31), A2 => n156, B1 => B(31), B2 => n152, 
                           ZN => n20);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUL is

   port( CLOCK : in std_logic;  A, B : in std_logic_vector (15 downto 0);  Y : 
         out std_logic_vector (31 downto 0));

end MUL;

architecture SYN_BEHAVIORAL of MUL is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_1
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_4
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_2
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_5
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_6
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_3
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_7
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component MUX5to1_NBIT32_1
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_2
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_3
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_4
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_5
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_6
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_7
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_8
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component ENCODER_1
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_2
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_3
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_4
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_5
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_6
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_7
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_0
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, A_neg_9_24_port, A_neg_9_23_port, 
      A_neg_9_22_port, A_neg_9_21_port, A_neg_9_20_port, A_neg_9_19_port, 
      A_neg_9_18_port, A_neg_9_17_port, A_neg_9_16_port, A_neg_9_15_port, 
      A_neg_9_14_port, A_neg_9_13_port, A_neg_9_12_port, A_neg_9_11_port, 
      A_neg_9_10_port, mux_out_7_31_port, mux_out_7_30_port, mux_out_7_29_port,
      mux_out_7_28_port, mux_out_7_27_port, mux_out_7_26_port, 
      mux_out_7_25_port, mux_out_7_24_port, mux_out_7_23_port, 
      mux_out_7_22_port, mux_out_7_21_port, mux_out_7_20_port, 
      mux_out_7_19_port, mux_out_7_18_port, mux_out_7_17_port, 
      mux_out_7_16_port, mux_out_7_15_port, mux_out_7_14_port, 
      mux_out_7_13_port, mux_out_7_12_port, mux_out_7_11_port, 
      mux_out_7_10_port, mux_out_7_9_port, mux_out_7_8_port, mux_out_7_7_port, 
      mux_out_7_6_port, mux_out_7_5_port, mux_out_7_4_port, mux_out_7_3_port, 
      mux_out_7_2_port, mux_out_7_1_port, mux_out_7_0_port, mux_out_6_31_port, 
      mux_out_6_30_port, mux_out_6_29_port, mux_out_6_28_port, 
      mux_out_6_27_port, mux_out_6_26_port, mux_out_6_25_port, 
      mux_out_6_24_port, mux_out_6_23_port, mux_out_6_22_port, 
      mux_out_6_21_port, mux_out_6_20_port, mux_out_6_19_port, 
      mux_out_6_18_port, mux_out_6_17_port, mux_out_6_16_port, 
      mux_out_6_15_port, mux_out_6_14_port, mux_out_6_13_port, 
      mux_out_6_12_port, mux_out_6_11_port, mux_out_6_10_port, mux_out_6_9_port
      , mux_out_6_8_port, mux_out_6_7_port, mux_out_6_6_port, mux_out_6_5_port,
      mux_out_6_4_port, mux_out_6_3_port, mux_out_6_2_port, mux_out_6_1_port, 
      mux_out_6_0_port, mux_out_5_31_port, mux_out_5_30_port, mux_out_5_29_port
      , mux_out_5_28_port, mux_out_5_27_port, mux_out_5_26_port, 
      mux_out_5_25_port, mux_out_5_24_port, mux_out_5_23_port, 
      mux_out_5_22_port, mux_out_5_21_port, mux_out_5_20_port, 
      mux_out_5_19_port, mux_out_5_18_port, mux_out_5_17_port, 
      mux_out_5_16_port, mux_out_5_15_port, mux_out_5_14_port, 
      mux_out_5_13_port, mux_out_5_12_port, mux_out_5_11_port, 
      mux_out_5_10_port, mux_out_5_9_port, mux_out_5_8_port, mux_out_5_7_port, 
      mux_out_5_6_port, mux_out_5_5_port, mux_out_5_4_port, mux_out_5_3_port, 
      mux_out_5_2_port, mux_out_5_1_port, mux_out_5_0_port, mux_out_4_31_port, 
      mux_out_4_30_port, mux_out_4_29_port, mux_out_4_28_port, 
      mux_out_4_27_port, mux_out_4_26_port, mux_out_4_25_port, 
      mux_out_4_24_port, mux_out_4_23_port, mux_out_4_22_port, 
      mux_out_4_21_port, mux_out_4_20_port, mux_out_4_19_port, 
      mux_out_4_18_port, mux_out_4_17_port, mux_out_4_16_port, 
      mux_out_4_15_port, mux_out_4_14_port, mux_out_4_13_port, 
      mux_out_4_12_port, mux_out_4_11_port, mux_out_4_10_port, mux_out_4_9_port
      , mux_out_4_8_port, mux_out_4_7_port, mux_out_4_6_port, mux_out_4_5_port,
      mux_out_4_4_port, mux_out_4_3_port, mux_out_4_2_port, mux_out_4_1_port, 
      mux_out_4_0_port, mux_out_3_31_port, mux_out_3_30_port, mux_out_3_29_port
      , mux_out_3_28_port, mux_out_3_27_port, mux_out_3_26_port, 
      mux_out_3_25_port, mux_out_3_24_port, mux_out_3_23_port, 
      mux_out_3_22_port, mux_out_3_21_port, mux_out_3_20_port, 
      mux_out_3_19_port, mux_out_3_18_port, mux_out_3_17_port, 
      mux_out_3_16_port, mux_out_3_15_port, mux_out_3_14_port, 
      mux_out_3_13_port, mux_out_3_12_port, mux_out_3_11_port, 
      mux_out_3_10_port, mux_out_3_9_port, mux_out_3_8_port, mux_out_3_7_port, 
      mux_out_3_6_port, mux_out_3_5_port, mux_out_3_4_port, mux_out_3_3_port, 
      mux_out_3_2_port, mux_out_3_1_port, mux_out_3_0_port, mux_out_2_31_port, 
      mux_out_2_30_port, mux_out_2_29_port, mux_out_2_28_port, 
      mux_out_2_27_port, mux_out_2_26_port, mux_out_2_25_port, 
      mux_out_2_24_port, mux_out_2_23_port, mux_out_2_22_port, 
      mux_out_2_21_port, mux_out_2_20_port, mux_out_2_19_port, 
      mux_out_2_18_port, mux_out_2_17_port, mux_out_2_16_port, 
      mux_out_2_15_port, mux_out_2_14_port, mux_out_2_13_port, 
      mux_out_2_12_port, mux_out_2_11_port, mux_out_2_10_port, mux_out_2_9_port
      , mux_out_2_8_port, mux_out_2_7_port, mux_out_2_6_port, mux_out_2_5_port,
      mux_out_2_4_port, mux_out_2_3_port, mux_out_2_2_port, mux_out_2_1_port, 
      mux_out_2_0_port, addends_7_31_port, addends_7_30_port, addends_7_29_port
      , addends_7_28_port, addends_7_27_port, addends_7_26_port, 
      addends_7_25_port, addends_7_24_port, addends_7_23_port, 
      addends_7_22_port, addends_7_21_port, addends_7_20_port, 
      addends_7_19_port, addends_7_18_port, addends_7_17_port, 
      addends_7_16_port, addends_7_15_port, addends_7_14_port, 
      addends_7_13_port, addends_7_12_port, addends_7_11_port, 
      addends_7_10_port, addends_7_9_port, addends_7_8_port, addends_7_7_port, 
      addends_7_6_port, addends_7_5_port, addends_7_4_port, addends_7_3_port, 
      addends_7_2_port, addends_7_1_port, addends_7_0_port, addends_6_31_port, 
      addends_6_30_port, addends_6_29_port, addends_6_28_port, 
      addends_6_27_port, addends_6_26_port, addends_6_25_port, 
      addends_6_24_port, addends_6_23_port, addends_6_22_port, 
      addends_6_21_port, addends_6_20_port, addends_6_19_port, 
      addends_6_18_port, addends_6_17_port, addends_6_16_port, 
      addends_6_15_port, addends_6_14_port, addends_6_13_port, 
      addends_6_12_port, addends_6_11_port, addends_6_10_port, addends_6_9_port
      , addends_6_8_port, addends_6_7_port, addends_6_6_port, addends_6_5_port,
      addends_6_4_port, addends_6_3_port, addends_6_2_port, addends_6_1_port, 
      addends_6_0_port, addends_5_31_port, addends_5_30_port, addends_5_29_port
      , addends_5_28_port, addends_5_27_port, addends_5_26_port, 
      addends_5_25_port, addends_5_24_port, addends_5_23_port, 
      addends_5_22_port, addends_5_21_port, addends_5_20_port, 
      addends_5_19_port, addends_5_18_port, addends_5_17_port, 
      addends_5_16_port, addends_5_15_port, addends_5_14_port, 
      addends_5_13_port, addends_5_12_port, addends_5_11_port, 
      addends_5_10_port, addends_5_9_port, addends_5_8_port, addends_5_7_port, 
      addends_5_6_port, addends_5_5_port, addends_5_4_port, addends_5_3_port, 
      addends_5_2_port, addends_5_1_port, addends_5_0_port, addends_4_31_port, 
      addends_4_30_port, addends_4_29_port, addends_4_28_port, 
      addends_4_27_port, addends_4_26_port, addends_4_25_port, 
      addends_4_24_port, addends_4_23_port, addends_4_22_port, 
      addends_4_21_port, addends_4_20_port, addends_4_19_port, 
      addends_4_18_port, addends_4_17_port, addends_4_16_port, 
      addends_4_15_port, addends_4_14_port, addends_4_13_port, 
      addends_4_12_port, addends_4_11_port, addends_4_10_port, addends_4_9_port
      , addends_4_8_port, addends_4_7_port, addends_4_6_port, addends_4_5_port,
      addends_4_4_port, addends_4_3_port, addends_4_2_port, addends_4_1_port, 
      addends_4_0_port, addends_3_31_port, addends_3_30_port, addends_3_29_port
      , addends_3_28_port, addends_3_27_port, addends_3_26_port, 
      addends_3_25_port, addends_3_24_port, addends_3_23_port, 
      addends_3_22_port, addends_3_21_port, addends_3_20_port, 
      addends_3_19_port, addends_3_18_port, addends_3_17_port, 
      addends_3_16_port, addends_3_15_port, addends_3_14_port, 
      addends_3_13_port, addends_3_12_port, addends_3_11_port, 
      addends_3_10_port, addends_3_9_port, addends_3_8_port, addends_3_7_port, 
      addends_3_6_port, addends_3_5_port, addends_3_4_port, addends_3_3_port, 
      addends_3_2_port, addends_3_1_port, addends_3_0_port, addends_2_31_port, 
      addends_2_30_port, addends_2_29_port, addends_2_28_port, 
      addends_2_27_port, addends_2_26_port, addends_2_25_port, 
      addends_2_24_port, addends_2_23_port, addends_2_22_port, 
      addends_2_21_port, addends_2_20_port, addends_2_19_port, 
      addends_2_18_port, addends_2_17_port, addends_2_16_port, 
      addends_2_15_port, addends_2_14_port, addends_2_13_port, 
      addends_2_12_port, addends_2_11_port, addends_2_10_port, addends_2_9_port
      , addends_2_8_port, addends_2_7_port, addends_2_6_port, addends_2_5_port,
      addends_2_4_port, addends_2_3_port, addends_2_2_port, addends_2_1_port, 
      addends_2_0_port, addends_1_31_port, addends_1_30_port, addends_1_29_port
      , addends_1_28_port, addends_1_27_port, addends_1_26_port, 
      addends_1_25_port, addends_1_24_port, addends_1_23_port, 
      addends_1_22_port, addends_1_21_port, addends_1_20_port, 
      addends_1_19_port, addends_1_18_port, addends_1_17_port, 
      addends_1_16_port, addends_1_15_port, addends_1_14_port, 
      addends_1_13_port, addends_1_12_port, addends_1_11_port, 
      addends_1_10_port, addends_1_9_port, addends_1_8_port, addends_1_7_port, 
      addends_1_6_port, addends_1_5_port, addends_1_4_port, addends_1_3_port, 
      addends_1_2_port, addends_1_1_port, addends_1_0_port, addends_0_31_port, 
      addends_0_30_port, addends_0_29_port, addends_0_28_port, 
      addends_0_27_port, addends_0_26_port, addends_0_25_port, 
      addends_0_24_port, addends_0_23_port, addends_0_22_port, 
      addends_0_21_port, addends_0_20_port, addends_0_19_port, 
      addends_0_18_port, addends_0_17_port, addends_0_16_port, 
      addends_0_15_port, addends_0_14_port, addends_0_13_port, 
      addends_0_12_port, addends_0_11_port, addends_0_10_port, addends_0_9_port
      , addends_0_8_port, addends_0_7_port, addends_0_6_port, addends_0_5_port,
      addends_0_4_port, addends_0_3_port, addends_0_2_port, addends_0_1_port, 
      addends_0_0_port, pipe1_3_31_port, pipe1_3_30_port, pipe1_3_29_port, 
      pipe1_3_28_port, pipe1_3_27_port, pipe1_3_26_port, pipe1_3_25_port, 
      pipe1_3_24_port, pipe1_3_23_port, pipe1_3_22_port, pipe1_3_21_port, 
      pipe1_3_20_port, pipe1_3_19_port, pipe1_3_18_port, pipe1_3_17_port, 
      pipe1_3_16_port, pipe1_3_15_port, pipe1_3_14_port, pipe1_3_13_port, 
      pipe1_3_12_port, pipe1_3_11_port, pipe1_3_10_port, pipe1_3_9_port, 
      pipe1_3_8_port, pipe1_3_7_port, pipe1_3_6_port, pipe1_3_5_port, 
      pipe1_3_4_port, pipe1_3_3_port, pipe1_3_2_port, pipe1_3_1_port, 
      pipe1_3_0_port, pipe1_2_31_port, pipe1_2_30_port, pipe1_2_29_port, 
      pipe1_2_28_port, pipe1_2_27_port, pipe1_2_26_port, pipe1_2_25_port, 
      pipe1_2_24_port, pipe1_2_23_port, pipe1_2_22_port, pipe1_2_21_port, 
      pipe1_2_20_port, pipe1_2_19_port, pipe1_2_18_port, pipe1_2_17_port, 
      pipe1_2_16_port, pipe1_2_15_port, pipe1_2_14_port, pipe1_2_13_port, 
      pipe1_2_12_port, pipe1_2_11_port, pipe1_2_10_port, pipe1_2_9_port, 
      pipe1_2_8_port, pipe1_2_7_port, pipe1_2_6_port, pipe1_2_5_port, 
      pipe1_2_4_port, pipe1_2_3_port, pipe1_2_2_port, pipe1_2_1_port, 
      pipe1_2_0_port, pipe1_1_31_port, pipe1_1_30_port, pipe1_1_29_port, 
      pipe1_1_28_port, pipe1_1_27_port, pipe1_1_26_port, pipe1_1_25_port, 
      pipe1_1_24_port, pipe1_1_23_port, pipe1_1_22_port, pipe1_1_21_port, 
      pipe1_1_20_port, pipe1_1_19_port, pipe1_1_18_port, pipe1_1_17_port, 
      pipe1_1_16_port, pipe1_1_15_port, pipe1_1_14_port, pipe1_1_13_port, 
      pipe1_1_12_port, pipe1_1_11_port, pipe1_1_10_port, pipe1_1_9_port, 
      pipe1_1_8_port, pipe1_1_7_port, pipe1_1_6_port, pipe1_1_5_port, 
      pipe1_1_4_port, pipe1_1_3_port, pipe1_1_2_port, pipe1_1_1_port, 
      pipe1_1_0_port, pipe1_0_31_port, pipe1_0_30_port, pipe1_0_29_port, 
      pipe1_0_28_port, pipe1_0_27_port, pipe1_0_26_port, pipe1_0_25_port, 
      pipe1_0_24_port, pipe1_0_23_port, pipe1_0_22_port, pipe1_0_21_port, 
      pipe1_0_20_port, pipe1_0_19_port, pipe1_0_18_port, pipe1_0_17_port, 
      pipe1_0_16_port, pipe1_0_15_port, pipe1_0_14_port, pipe1_0_13_port, 
      pipe1_0_12_port, pipe1_0_11_port, pipe1_0_10_port, pipe1_0_9_port, 
      pipe1_0_8_port, pipe1_0_7_port, pipe1_0_6_port, pipe1_0_5_port, 
      pipe1_0_4_port, pipe1_0_3_port, pipe1_0_2_port, pipe1_0_1_port, 
      pipe1_0_0_port, pipe2_1_31_port, pipe2_1_30_port, pipe2_1_29_port, 
      pipe2_1_28_port, pipe2_1_27_port, pipe2_1_26_port, pipe2_1_25_port, 
      pipe2_1_24_port, pipe2_1_23_port, pipe2_1_22_port, pipe2_1_21_port, 
      pipe2_1_20_port, pipe2_1_19_port, pipe2_1_18_port, pipe2_1_17_port, 
      pipe2_1_16_port, pipe2_1_15_port, pipe2_1_14_port, pipe2_1_13_port, 
      pipe2_1_12_port, pipe2_1_11_port, pipe2_1_10_port, pipe2_1_9_port, 
      pipe2_1_8_port, pipe2_1_7_port, pipe2_1_6_port, pipe2_1_5_port, 
      pipe2_1_4_port, pipe2_1_3_port, pipe2_1_2_port, pipe2_1_1_port, 
      pipe2_1_0_port, pipe2_0_31_port, pipe2_0_30_port, pipe2_0_29_port, 
      pipe2_0_28_port, pipe2_0_27_port, pipe2_0_26_port, pipe2_0_25_port, 
      pipe2_0_24_port, pipe2_0_23_port, pipe2_0_22_port, pipe2_0_21_port, 
      pipe2_0_20_port, pipe2_0_19_port, pipe2_0_18_port, pipe2_0_17_port, 
      pipe2_0_16_port, pipe2_0_15_port, pipe2_0_14_port, pipe2_0_13_port, 
      pipe2_0_12_port, pipe2_0_11_port, pipe2_0_10_port, pipe2_0_9_port, 
      pipe2_0_8_port, pipe2_0_7_port, pipe2_0_6_port, pipe2_0_5_port, 
      pipe2_0_4_port, pipe2_0_3_port, pipe2_0_2_port, pipe2_0_1_port, 
      pipe2_0_0_port, selector_23_port, selector_22_port, selector_21_port, 
      selector_20_port, selector_19_port, selector_18_port, selector_17_port, 
      selector_16_port, selector_15_port, selector_14_port, selector_13_port, 
      selector_12_port, selector_11_port, selector_10_port, selector_9_port, 
      selector_8_port, selector_7_port, selector_6_port, selector_5_port, 
      selector_4_port, selector_3_port, selector_2_port, selector_1_port, 
      selector_0_port, reg_in_2_31_port, reg_in_2_30_port, reg_in_2_29_port, 
      reg_in_2_28_port, reg_in_2_27_port, reg_in_2_26_port, reg_in_2_25_port, 
      reg_in_2_24_port, reg_in_2_23_port, reg_in_2_22_port, reg_in_2_21_port, 
      reg_in_2_20_port, reg_in_2_19_port, reg_in_2_18_port, reg_in_2_17_port, 
      reg_in_2_16_port, reg_in_2_15_port, reg_in_2_14_port, reg_in_2_13_port, 
      reg_in_2_12_port, reg_in_2_11_port, reg_in_2_10_port, reg_in_2_9_port, 
      reg_in_2_8_port, reg_in_2_7_port, reg_in_2_6_port, reg_in_2_5_port, 
      reg_in_2_4_port, reg_in_2_3_port, reg_in_2_2_port, reg_in_2_1_port, 
      reg_in_2_0_port, reg_in_1_31_port, reg_in_1_30_port, reg_in_1_29_port, 
      reg_in_1_28_port, reg_in_1_27_port, reg_in_1_26_port, reg_in_1_25_port, 
      reg_in_1_24_port, reg_in_1_23_port, reg_in_1_22_port, reg_in_1_21_port, 
      reg_in_1_20_port, reg_in_1_19_port, reg_in_1_18_port, reg_in_1_17_port, 
      reg_in_1_16_port, reg_in_1_15_port, reg_in_1_14_port, reg_in_1_13_port, 
      reg_in_1_12_port, reg_in_1_11_port, reg_in_1_10_port, reg_in_1_9_port, 
      reg_in_1_8_port, reg_in_1_7_port, reg_in_1_6_port, reg_in_1_5_port, 
      reg_in_1_4_port, reg_in_1_3_port, reg_in_1_2_port, reg_in_1_1_port, 
      reg_in_1_0_port, reg_in_0_31_port, reg_in_0_30_port, reg_in_0_29_port, 
      reg_in_0_28_port, reg_in_0_27_port, reg_in_0_26_port, reg_in_0_25_port, 
      reg_in_0_24_port, reg_in_0_23_port, reg_in_0_22_port, reg_in_0_21_port, 
      reg_in_0_20_port, reg_in_0_19_port, reg_in_0_18_port, reg_in_0_17_port, 
      reg_in_0_16_port, reg_in_0_15_port, reg_in_0_14_port, reg_in_0_13_port, 
      reg_in_0_12_port, reg_in_0_11_port, reg_in_0_10_port, reg_in_0_9_port, 
      reg_in_0_8_port, reg_in_0_7_port, reg_in_0_6_port, reg_in_0_5_port, 
      reg_in_0_4_port, reg_in_0_3_port, reg_in_0_2_port, reg_in_0_1_port, 
      reg_in_0_0_port, reg_out_2_31_port, reg_out_2_30_port, reg_out_2_29_port,
      reg_out_2_28_port, reg_out_2_27_port, reg_out_2_26_port, 
      reg_out_2_25_port, reg_out_2_24_port, reg_out_2_23_port, 
      reg_out_2_22_port, reg_out_2_21_port, reg_out_2_20_port, 
      reg_out_2_19_port, reg_out_2_18_port, reg_out_2_17_port, 
      reg_out_2_16_port, reg_out_2_15_port, reg_out_2_14_port, 
      reg_out_2_13_port, reg_out_2_12_port, reg_out_2_11_port, 
      reg_out_2_10_port, reg_out_2_9_port, reg_out_2_8_port, reg_out_2_7_port, 
      reg_out_2_6_port, reg_out_2_5_port, reg_out_2_4_port, reg_out_2_3_port, 
      reg_out_2_2_port, reg_out_2_1_port, reg_out_2_0_port, reg_out_1_31_port, 
      reg_out_1_30_port, reg_out_1_29_port, reg_out_1_28_port, 
      reg_out_1_27_port, reg_out_1_26_port, reg_out_1_25_port, 
      reg_out_1_24_port, reg_out_1_23_port, reg_out_1_22_port, 
      reg_out_1_21_port, reg_out_1_20_port, reg_out_1_19_port, 
      reg_out_1_18_port, reg_out_1_17_port, reg_out_1_16_port, 
      reg_out_1_15_port, reg_out_1_14_port, reg_out_1_13_port, 
      reg_out_1_12_port, reg_out_1_11_port, reg_out_1_10_port, reg_out_1_9_port
      , reg_out_1_8_port, reg_out_1_7_port, reg_out_1_6_port, reg_out_1_5_port,
      reg_out_1_4_port, reg_out_1_3_port, reg_out_1_2_port, reg_out_1_1_port, 
      reg_out_1_0_port, reg_out_0_31_port, reg_out_0_30_port, reg_out_0_29_port
      , reg_out_0_28_port, reg_out_0_27_port, reg_out_0_26_port, 
      reg_out_0_25_port, reg_out_0_24_port, reg_out_0_23_port, 
      reg_out_0_22_port, reg_out_0_21_port, reg_out_0_20_port, 
      reg_out_0_19_port, reg_out_0_18_port, reg_out_0_17_port, 
      reg_out_0_16_port, reg_out_0_15_port, reg_out_0_14_port, 
      reg_out_0_13_port, reg_out_0_12_port, reg_out_0_11_port, 
      reg_out_0_10_port, reg_out_0_9_port, reg_out_0_8_port, reg_out_0_7_port, 
      reg_out_0_6_port, reg_out_0_5_port, reg_out_0_4_port, reg_out_0_3_port, 
      reg_out_0_2_port, reg_out_0_1_port, reg_out_0_0_port, add_out_2_31_port, 
      add_out_2_30_port, add_out_2_29_port, add_out_2_28_port, 
      add_out_2_27_port, add_out_2_26_port, add_out_2_25_port, 
      add_out_2_24_port, add_out_2_23_port, add_out_2_22_port, 
      add_out_2_21_port, add_out_2_20_port, add_out_2_19_port, 
      add_out_2_18_port, add_out_2_17_port, add_out_2_16_port, 
      add_out_2_15_port, add_out_2_14_port, add_out_2_13_port, 
      add_out_2_12_port, add_out_2_11_port, add_out_2_10_port, add_out_2_9_port
      , add_out_2_8_port, add_out_2_7_port, add_out_2_6_port, add_out_2_5_port,
      add_out_2_4_port, add_out_2_3_port, add_out_2_2_port, add_out_2_1_port, 
      add_out_2_0_port, add_out_1_31_port, add_out_1_30_port, add_out_1_29_port
      , add_out_1_28_port, add_out_1_27_port, add_out_1_26_port, 
      add_out_1_25_port, add_out_1_24_port, add_out_1_23_port, 
      add_out_1_22_port, add_out_1_21_port, add_out_1_20_port, 
      add_out_1_19_port, add_out_1_18_port, add_out_1_17_port, 
      add_out_1_16_port, add_out_1_15_port, add_out_1_14_port, 
      add_out_1_13_port, add_out_1_12_port, add_out_1_11_port, 
      add_out_1_10_port, add_out_1_9_port, add_out_1_8_port, add_out_1_7_port, 
      add_out_1_6_port, add_out_1_5_port, add_out_1_4_port, add_out_1_3_port, 
      add_out_1_2_port, add_out_1_1_port, add_out_1_0_port, add_out_0_31_port, 
      add_out_0_30_port, add_out_0_29_port, add_out_0_28_port, 
      add_out_0_27_port, add_out_0_26_port, add_out_0_25_port, 
      add_out_0_24_port, add_out_0_23_port, add_out_0_22_port, 
      add_out_0_21_port, add_out_0_20_port, add_out_0_19_port, 
      add_out_0_18_port, add_out_0_17_port, add_out_0_16_port, 
      add_out_0_15_port, add_out_0_14_port, add_out_0_13_port, 
      add_out_0_12_port, add_out_0_11_port, add_out_0_10_port, add_out_0_9_port
      , add_out_0_8_port, add_out_0_7_port, add_out_0_6_port, add_out_0_5_port,
      add_out_0_4_port, add_out_0_3_port, add_out_0_2_port, add_out_0_1_port, 
      add_out_0_0_port, n9, n69, n4, n5, n7, n8, n10, n12, n14, n16, n18, n19, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144
      , n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153,
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526, n_1527 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   addends_reg_3_31_inst : DFF_X1 port map( D => mux_out_3_31_port, CK => CLOCK
                           , Q => addends_3_31_port, QN => n_1137);
   addends_reg_3_30_inst : DFF_X1 port map( D => mux_out_3_30_port, CK => CLOCK
                           , Q => addends_3_30_port, QN => n_1138);
   addends_reg_3_29_inst : DFF_X1 port map( D => mux_out_3_29_port, CK => CLOCK
                           , Q => addends_3_29_port, QN => n_1139);
   addends_reg_3_28_inst : DFF_X1 port map( D => mux_out_3_28_port, CK => CLOCK
                           , Q => addends_3_28_port, QN => n_1140);
   addends_reg_3_27_inst : DFF_X1 port map( D => mux_out_3_27_port, CK => CLOCK
                           , Q => addends_3_27_port, QN => n_1141);
   addends_reg_3_26_inst : DFF_X1 port map( D => mux_out_3_26_port, CK => CLOCK
                           , Q => addends_3_26_port, QN => n_1142);
   addends_reg_3_25_inst : DFF_X1 port map( D => mux_out_3_25_port, CK => CLOCK
                           , Q => addends_3_25_port, QN => n_1143);
   addends_reg_3_24_inst : DFF_X1 port map( D => mux_out_3_24_port, CK => CLOCK
                           , Q => addends_3_24_port, QN => n_1144);
   addends_reg_3_23_inst : DFF_X1 port map( D => mux_out_3_23_port, CK => CLOCK
                           , Q => addends_3_23_port, QN => n_1145);
   addends_reg_3_22_inst : DFF_X1 port map( D => mux_out_3_22_port, CK => CLOCK
                           , Q => addends_3_22_port, QN => n_1146);
   addends_reg_3_21_inst : DFF_X1 port map( D => mux_out_3_21_port, CK => CLOCK
                           , Q => addends_3_21_port, QN => n_1147);
   addends_reg_3_20_inst : DFF_X1 port map( D => mux_out_3_20_port, CK => CLOCK
                           , Q => addends_3_20_port, QN => n_1148);
   addends_reg_3_19_inst : DFF_X1 port map( D => mux_out_3_19_port, CK => CLOCK
                           , Q => addends_3_19_port, QN => n_1149);
   addends_reg_3_18_inst : DFF_X1 port map( D => mux_out_3_18_port, CK => CLOCK
                           , Q => addends_3_18_port, QN => n_1150);
   addends_reg_3_17_inst : DFF_X1 port map( D => mux_out_3_17_port, CK => CLOCK
                           , Q => addends_3_17_port, QN => n_1151);
   addends_reg_3_16_inst : DFF_X1 port map( D => mux_out_3_16_port, CK => CLOCK
                           , Q => addends_3_16_port, QN => n_1152);
   addends_reg_3_15_inst : DFF_X1 port map( D => mux_out_3_15_port, CK => CLOCK
                           , Q => addends_3_15_port, QN => n_1153);
   addends_reg_3_14_inst : DFF_X1 port map( D => mux_out_3_14_port, CK => CLOCK
                           , Q => addends_3_14_port, QN => n_1154);
   addends_reg_3_13_inst : DFF_X1 port map( D => mux_out_3_13_port, CK => CLOCK
                           , Q => addends_3_13_port, QN => n_1155);
   addends_reg_3_12_inst : DFF_X1 port map( D => mux_out_3_12_port, CK => CLOCK
                           , Q => addends_3_12_port, QN => n_1156);
   addends_reg_3_11_inst : DFF_X1 port map( D => mux_out_3_11_port, CK => CLOCK
                           , Q => addends_3_11_port, QN => n_1157);
   addends_reg_3_10_inst : DFF_X1 port map( D => mux_out_3_10_port, CK => CLOCK
                           , Q => addends_3_10_port, QN => n_1158);
   addends_reg_3_9_inst : DFF_X1 port map( D => mux_out_3_9_port, CK => CLOCK, 
                           Q => addends_3_9_port, QN => n_1159);
   addends_reg_3_8_inst : DFF_X1 port map( D => mux_out_3_8_port, CK => CLOCK, 
                           Q => addends_3_8_port, QN => n_1160);
   addends_reg_3_7_inst : DFF_X1 port map( D => mux_out_3_7_port, CK => CLOCK, 
                           Q => addends_3_7_port, QN => n_1161);
   addends_reg_3_6_inst : DFF_X1 port map( D => mux_out_3_6_port, CK => CLOCK, 
                           Q => addends_3_6_port, QN => n_1162);
   addends_reg_3_5_inst : DFF_X1 port map( D => mux_out_3_5_port, CK => CLOCK, 
                           Q => addends_3_5_port, QN => n_1163);
   addends_reg_3_4_inst : DFF_X1 port map( D => mux_out_3_4_port, CK => CLOCK, 
                           Q => addends_3_4_port, QN => n_1164);
   addends_reg_3_3_inst : DFF_X1 port map( D => mux_out_3_3_port, CK => CLOCK, 
                           Q => addends_3_3_port, QN => n_1165);
   addends_reg_3_2_inst : DFF_X1 port map( D => mux_out_3_2_port, CK => CLOCK, 
                           Q => addends_3_2_port, QN => n_1166);
   addends_reg_3_1_inst : DFF_X1 port map( D => mux_out_3_1_port, CK => CLOCK, 
                           Q => addends_3_1_port, QN => n_1167);
   addends_reg_3_0_inst : DFF_X1 port map( D => mux_out_3_0_port, CK => CLOCK, 
                           Q => addends_3_0_port, QN => n_1168);
   addends_reg_2_31_inst : DFF_X1 port map( D => mux_out_2_31_port, CK => CLOCK
                           , Q => addends_2_31_port, QN => n_1169);
   addends_reg_2_30_inst : DFF_X1 port map( D => mux_out_2_30_port, CK => CLOCK
                           , Q => addends_2_30_port, QN => n_1170);
   addends_reg_2_29_inst : DFF_X1 port map( D => mux_out_2_29_port, CK => CLOCK
                           , Q => addends_2_29_port, QN => n_1171);
   addends_reg_2_28_inst : DFF_X1 port map( D => mux_out_2_28_port, CK => CLOCK
                           , Q => addends_2_28_port, QN => n_1172);
   addends_reg_2_27_inst : DFF_X1 port map( D => mux_out_2_27_port, CK => CLOCK
                           , Q => addends_2_27_port, QN => n_1173);
   addends_reg_2_26_inst : DFF_X1 port map( D => mux_out_2_26_port, CK => CLOCK
                           , Q => addends_2_26_port, QN => n_1174);
   addends_reg_2_25_inst : DFF_X1 port map( D => mux_out_2_25_port, CK => CLOCK
                           , Q => addends_2_25_port, QN => n_1175);
   addends_reg_2_24_inst : DFF_X1 port map( D => mux_out_2_24_port, CK => CLOCK
                           , Q => addends_2_24_port, QN => n_1176);
   addends_reg_2_23_inst : DFF_X1 port map( D => mux_out_2_23_port, CK => CLOCK
                           , Q => addends_2_23_port, QN => n_1177);
   addends_reg_2_22_inst : DFF_X1 port map( D => mux_out_2_22_port, CK => CLOCK
                           , Q => addends_2_22_port, QN => n_1178);
   addends_reg_2_21_inst : DFF_X1 port map( D => mux_out_2_21_port, CK => CLOCK
                           , Q => addends_2_21_port, QN => n_1179);
   addends_reg_2_20_inst : DFF_X1 port map( D => mux_out_2_20_port, CK => CLOCK
                           , Q => addends_2_20_port, QN => n_1180);
   addends_reg_2_19_inst : DFF_X1 port map( D => mux_out_2_19_port, CK => CLOCK
                           , Q => addends_2_19_port, QN => n_1181);
   addends_reg_2_18_inst : DFF_X1 port map( D => mux_out_2_18_port, CK => CLOCK
                           , Q => addends_2_18_port, QN => n_1182);
   addends_reg_2_17_inst : DFF_X1 port map( D => mux_out_2_17_port, CK => CLOCK
                           , Q => addends_2_17_port, QN => n_1183);
   addends_reg_2_16_inst : DFF_X1 port map( D => mux_out_2_16_port, CK => CLOCK
                           , Q => addends_2_16_port, QN => n_1184);
   addends_reg_2_15_inst : DFF_X1 port map( D => mux_out_2_15_port, CK => CLOCK
                           , Q => addends_2_15_port, QN => n_1185);
   addends_reg_2_14_inst : DFF_X1 port map( D => mux_out_2_14_port, CK => CLOCK
                           , Q => addends_2_14_port, QN => n_1186);
   addends_reg_2_13_inst : DFF_X1 port map( D => mux_out_2_13_port, CK => CLOCK
                           , Q => addends_2_13_port, QN => n_1187);
   addends_reg_2_12_inst : DFF_X1 port map( D => mux_out_2_12_port, CK => CLOCK
                           , Q => addends_2_12_port, QN => n_1188);
   addends_reg_2_11_inst : DFF_X1 port map( D => mux_out_2_11_port, CK => CLOCK
                           , Q => addends_2_11_port, QN => n_1189);
   addends_reg_2_10_inst : DFF_X1 port map( D => mux_out_2_10_port, CK => CLOCK
                           , Q => addends_2_10_port, QN => n_1190);
   addends_reg_2_9_inst : DFF_X1 port map( D => mux_out_2_9_port, CK => CLOCK, 
                           Q => addends_2_9_port, QN => n_1191);
   addends_reg_2_8_inst : DFF_X1 port map( D => mux_out_2_8_port, CK => CLOCK, 
                           Q => addends_2_8_port, QN => n_1192);
   addends_reg_2_7_inst : DFF_X1 port map( D => mux_out_2_7_port, CK => CLOCK, 
                           Q => addends_2_7_port, QN => n_1193);
   addends_reg_2_6_inst : DFF_X1 port map( D => mux_out_2_6_port, CK => CLOCK, 
                           Q => addends_2_6_port, QN => n_1194);
   addends_reg_2_5_inst : DFF_X1 port map( D => mux_out_2_5_port, CK => CLOCK, 
                           Q => addends_2_5_port, QN => n_1195);
   addends_reg_2_4_inst : DFF_X1 port map( D => mux_out_2_4_port, CK => CLOCK, 
                           Q => addends_2_4_port, QN => n_1196);
   addends_reg_2_3_inst : DFF_X1 port map( D => mux_out_2_3_port, CK => CLOCK, 
                           Q => addends_2_3_port, QN => n_1197);
   addends_reg_2_2_inst : DFF_X1 port map( D => mux_out_2_2_port, CK => CLOCK, 
                           Q => addends_2_2_port, QN => n_1198);
   addends_reg_2_1_inst : DFF_X1 port map( D => mux_out_2_1_port, CK => CLOCK, 
                           Q => addends_2_1_port, QN => n_1199);
   addends_reg_2_0_inst : DFF_X1 port map( D => mux_out_2_0_port, CK => CLOCK, 
                           Q => addends_2_0_port, QN => n_1200);
   pipe1_reg_3_31_inst : DFF_X1 port map( D => mux_out_7_31_port, CK => CLOCK, 
                           Q => pipe1_3_31_port, QN => n_1201);
   pipe1_reg_3_30_inst : DFF_X1 port map( D => mux_out_7_30_port, CK => CLOCK, 
                           Q => pipe1_3_30_port, QN => n_1202);
   pipe1_reg_3_29_inst : DFF_X1 port map( D => mux_out_7_29_port, CK => CLOCK, 
                           Q => pipe1_3_29_port, QN => n_1203);
   pipe1_reg_3_28_inst : DFF_X1 port map( D => mux_out_7_28_port, CK => CLOCK, 
                           Q => pipe1_3_28_port, QN => n_1204);
   pipe1_reg_3_27_inst : DFF_X1 port map( D => mux_out_7_27_port, CK => CLOCK, 
                           Q => pipe1_3_27_port, QN => n_1205);
   pipe1_reg_3_26_inst : DFF_X1 port map( D => mux_out_7_26_port, CK => CLOCK, 
                           Q => pipe1_3_26_port, QN => n_1206);
   pipe1_reg_3_25_inst : DFF_X1 port map( D => mux_out_7_25_port, CK => CLOCK, 
                           Q => pipe1_3_25_port, QN => n_1207);
   pipe1_reg_3_24_inst : DFF_X1 port map( D => mux_out_7_24_port, CK => CLOCK, 
                           Q => pipe1_3_24_port, QN => n_1208);
   pipe1_reg_3_23_inst : DFF_X1 port map( D => mux_out_7_23_port, CK => CLOCK, 
                           Q => pipe1_3_23_port, QN => n_1209);
   pipe1_reg_3_22_inst : DFF_X1 port map( D => mux_out_7_22_port, CK => CLOCK, 
                           Q => pipe1_3_22_port, QN => n_1210);
   pipe1_reg_3_21_inst : DFF_X1 port map( D => mux_out_7_21_port, CK => CLOCK, 
                           Q => pipe1_3_21_port, QN => n_1211);
   pipe1_reg_3_20_inst : DFF_X1 port map( D => mux_out_7_20_port, CK => CLOCK, 
                           Q => pipe1_3_20_port, QN => n_1212);
   pipe1_reg_3_19_inst : DFF_X1 port map( D => mux_out_7_19_port, CK => CLOCK, 
                           Q => pipe1_3_19_port, QN => n_1213);
   pipe1_reg_3_18_inst : DFF_X1 port map( D => mux_out_7_18_port, CK => CLOCK, 
                           Q => pipe1_3_18_port, QN => n_1214);
   pipe1_reg_3_17_inst : DFF_X1 port map( D => mux_out_7_17_port, CK => CLOCK, 
                           Q => pipe1_3_17_port, QN => n_1215);
   pipe1_reg_3_16_inst : DFF_X1 port map( D => mux_out_7_16_port, CK => CLOCK, 
                           Q => pipe1_3_16_port, QN => n_1216);
   pipe1_reg_3_15_inst : DFF_X1 port map( D => mux_out_7_15_port, CK => CLOCK, 
                           Q => pipe1_3_15_port, QN => n_1217);
   pipe1_reg_3_14_inst : DFF_X1 port map( D => mux_out_7_14_port, CK => CLOCK, 
                           Q => pipe1_3_14_port, QN => n_1218);
   pipe1_reg_3_13_inst : DFF_X1 port map( D => mux_out_7_13_port, CK => CLOCK, 
                           Q => pipe1_3_13_port, QN => n_1219);
   pipe1_reg_3_12_inst : DFF_X1 port map( D => mux_out_7_12_port, CK => CLOCK, 
                           Q => pipe1_3_12_port, QN => n_1220);
   pipe1_reg_3_11_inst : DFF_X1 port map( D => mux_out_7_11_port, CK => CLOCK, 
                           Q => pipe1_3_11_port, QN => n_1221);
   pipe1_reg_3_10_inst : DFF_X1 port map( D => mux_out_7_10_port, CK => CLOCK, 
                           Q => pipe1_3_10_port, QN => n_1222);
   pipe1_reg_3_9_inst : DFF_X1 port map( D => mux_out_7_9_port, CK => CLOCK, Q 
                           => pipe1_3_9_port, QN => n_1223);
   pipe1_reg_3_8_inst : DFF_X1 port map( D => mux_out_7_8_port, CK => CLOCK, Q 
                           => pipe1_3_8_port, QN => n_1224);
   pipe1_reg_3_7_inst : DFF_X1 port map( D => mux_out_7_7_port, CK => CLOCK, Q 
                           => pipe1_3_7_port, QN => n_1225);
   pipe1_reg_3_6_inst : DFF_X1 port map( D => mux_out_7_6_port, CK => CLOCK, Q 
                           => pipe1_3_6_port, QN => n_1226);
   pipe1_reg_3_5_inst : DFF_X1 port map( D => mux_out_7_5_port, CK => CLOCK, Q 
                           => pipe1_3_5_port, QN => n_1227);
   pipe1_reg_3_4_inst : DFF_X1 port map( D => mux_out_7_4_port, CK => CLOCK, Q 
                           => pipe1_3_4_port, QN => n_1228);
   pipe1_reg_3_3_inst : DFF_X1 port map( D => mux_out_7_3_port, CK => CLOCK, Q 
                           => pipe1_3_3_port, QN => n_1229);
   pipe1_reg_3_2_inst : DFF_X1 port map( D => mux_out_7_2_port, CK => CLOCK, Q 
                           => pipe1_3_2_port, QN => n_1230);
   pipe1_reg_3_1_inst : DFF_X1 port map( D => mux_out_7_1_port, CK => CLOCK, Q 
                           => pipe1_3_1_port, QN => n_1231);
   pipe1_reg_3_0_inst : DFF_X1 port map( D => mux_out_7_0_port, CK => CLOCK, Q 
                           => pipe1_3_0_port, QN => n_1232);
   pipe1_reg_2_31_inst : DFF_X1 port map( D => mux_out_6_31_port, CK => CLOCK, 
                           Q => pipe1_2_31_port, QN => n_1233);
   pipe1_reg_2_30_inst : DFF_X1 port map( D => mux_out_6_30_port, CK => CLOCK, 
                           Q => pipe1_2_30_port, QN => n_1234);
   pipe1_reg_2_29_inst : DFF_X1 port map( D => mux_out_6_29_port, CK => CLOCK, 
                           Q => pipe1_2_29_port, QN => n_1235);
   pipe1_reg_2_28_inst : DFF_X1 port map( D => mux_out_6_28_port, CK => CLOCK, 
                           Q => pipe1_2_28_port, QN => n_1236);
   pipe1_reg_2_27_inst : DFF_X1 port map( D => mux_out_6_27_port, CK => CLOCK, 
                           Q => pipe1_2_27_port, QN => n_1237);
   pipe1_reg_2_26_inst : DFF_X1 port map( D => mux_out_6_26_port, CK => CLOCK, 
                           Q => pipe1_2_26_port, QN => n_1238);
   pipe1_reg_2_25_inst : DFF_X1 port map( D => mux_out_6_25_port, CK => CLOCK, 
                           Q => pipe1_2_25_port, QN => n_1239);
   pipe1_reg_2_24_inst : DFF_X1 port map( D => mux_out_6_24_port, CK => CLOCK, 
                           Q => pipe1_2_24_port, QN => n_1240);
   pipe1_reg_2_23_inst : DFF_X1 port map( D => mux_out_6_23_port, CK => CLOCK, 
                           Q => pipe1_2_23_port, QN => n_1241);
   pipe1_reg_2_22_inst : DFF_X1 port map( D => mux_out_6_22_port, CK => CLOCK, 
                           Q => pipe1_2_22_port, QN => n_1242);
   pipe1_reg_2_21_inst : DFF_X1 port map( D => mux_out_6_21_port, CK => CLOCK, 
                           Q => pipe1_2_21_port, QN => n_1243);
   pipe1_reg_2_20_inst : DFF_X1 port map( D => mux_out_6_20_port, CK => CLOCK, 
                           Q => pipe1_2_20_port, QN => n_1244);
   pipe1_reg_2_19_inst : DFF_X1 port map( D => mux_out_6_19_port, CK => CLOCK, 
                           Q => pipe1_2_19_port, QN => n_1245);
   pipe1_reg_2_18_inst : DFF_X1 port map( D => mux_out_6_18_port, CK => CLOCK, 
                           Q => pipe1_2_18_port, QN => n_1246);
   pipe1_reg_2_17_inst : DFF_X1 port map( D => mux_out_6_17_port, CK => CLOCK, 
                           Q => pipe1_2_17_port, QN => n_1247);
   pipe1_reg_2_16_inst : DFF_X1 port map( D => mux_out_6_16_port, CK => CLOCK, 
                           Q => pipe1_2_16_port, QN => n_1248);
   pipe1_reg_2_15_inst : DFF_X1 port map( D => mux_out_6_15_port, CK => CLOCK, 
                           Q => pipe1_2_15_port, QN => n_1249);
   pipe1_reg_2_14_inst : DFF_X1 port map( D => mux_out_6_14_port, CK => CLOCK, 
                           Q => pipe1_2_14_port, QN => n_1250);
   pipe1_reg_2_13_inst : DFF_X1 port map( D => mux_out_6_13_port, CK => CLOCK, 
                           Q => pipe1_2_13_port, QN => n_1251);
   pipe1_reg_2_12_inst : DFF_X1 port map( D => mux_out_6_12_port, CK => CLOCK, 
                           Q => pipe1_2_12_port, QN => n_1252);
   pipe1_reg_2_11_inst : DFF_X1 port map( D => mux_out_6_11_port, CK => CLOCK, 
                           Q => pipe1_2_11_port, QN => n_1253);
   pipe1_reg_2_10_inst : DFF_X1 port map( D => mux_out_6_10_port, CK => CLOCK, 
                           Q => pipe1_2_10_port, QN => n_1254);
   pipe1_reg_2_9_inst : DFF_X1 port map( D => mux_out_6_9_port, CK => CLOCK, Q 
                           => pipe1_2_9_port, QN => n_1255);
   pipe1_reg_2_8_inst : DFF_X1 port map( D => mux_out_6_8_port, CK => CLOCK, Q 
                           => pipe1_2_8_port, QN => n_1256);
   pipe1_reg_2_7_inst : DFF_X1 port map( D => mux_out_6_7_port, CK => CLOCK, Q 
                           => pipe1_2_7_port, QN => n_1257);
   pipe1_reg_2_6_inst : DFF_X1 port map( D => mux_out_6_6_port, CK => CLOCK, Q 
                           => pipe1_2_6_port, QN => n_1258);
   pipe1_reg_2_5_inst : DFF_X1 port map( D => mux_out_6_5_port, CK => CLOCK, Q 
                           => pipe1_2_5_port, QN => n_1259);
   pipe1_reg_2_4_inst : DFF_X1 port map( D => mux_out_6_4_port, CK => CLOCK, Q 
                           => pipe1_2_4_port, QN => n_1260);
   pipe1_reg_2_3_inst : DFF_X1 port map( D => mux_out_6_3_port, CK => CLOCK, Q 
                           => pipe1_2_3_port, QN => n_1261);
   pipe1_reg_2_2_inst : DFF_X1 port map( D => mux_out_6_2_port, CK => CLOCK, Q 
                           => pipe1_2_2_port, QN => n_1262);
   pipe1_reg_2_1_inst : DFF_X1 port map( D => mux_out_6_1_port, CK => CLOCK, Q 
                           => pipe1_2_1_port, QN => n_1263);
   pipe1_reg_2_0_inst : DFF_X1 port map( D => mux_out_6_0_port, CK => CLOCK, Q 
                           => pipe1_2_0_port, QN => n_1264);
   pipe1_reg_1_31_inst : DFF_X1 port map( D => mux_out_5_31_port, CK => CLOCK, 
                           Q => pipe1_1_31_port, QN => n_1265);
   addends_reg_5_31_inst : DFF_X1 port map( D => pipe1_1_31_port, CK => CLOCK, 
                           Q => addends_5_31_port, QN => n_1266);
   pipe1_reg_1_30_inst : DFF_X1 port map( D => mux_out_5_30_port, CK => CLOCK, 
                           Q => pipe1_1_30_port, QN => n_1267);
   addends_reg_5_30_inst : DFF_X1 port map( D => pipe1_1_30_port, CK => CLOCK, 
                           Q => addends_5_30_port, QN => n_1268);
   pipe1_reg_1_29_inst : DFF_X1 port map( D => mux_out_5_29_port, CK => CLOCK, 
                           Q => pipe1_1_29_port, QN => n_1269);
   addends_reg_5_29_inst : DFF_X1 port map( D => pipe1_1_29_port, CK => CLOCK, 
                           Q => addends_5_29_port, QN => n_1270);
   pipe1_reg_1_28_inst : DFF_X1 port map( D => mux_out_5_28_port, CK => CLOCK, 
                           Q => pipe1_1_28_port, QN => n_1271);
   addends_reg_5_28_inst : DFF_X1 port map( D => pipe1_1_28_port, CK => CLOCK, 
                           Q => addends_5_28_port, QN => n_1272);
   pipe1_reg_1_27_inst : DFF_X1 port map( D => mux_out_5_27_port, CK => CLOCK, 
                           Q => pipe1_1_27_port, QN => n_1273);
   addends_reg_5_27_inst : DFF_X1 port map( D => pipe1_1_27_port, CK => CLOCK, 
                           Q => addends_5_27_port, QN => n_1274);
   pipe1_reg_1_26_inst : DFF_X1 port map( D => mux_out_5_26_port, CK => CLOCK, 
                           Q => pipe1_1_26_port, QN => n_1275);
   addends_reg_5_26_inst : DFF_X1 port map( D => pipe1_1_26_port, CK => CLOCK, 
                           Q => addends_5_26_port, QN => n_1276);
   pipe1_reg_1_25_inst : DFF_X1 port map( D => mux_out_5_25_port, CK => CLOCK, 
                           Q => pipe1_1_25_port, QN => n_1277);
   addends_reg_5_25_inst : DFF_X1 port map( D => pipe1_1_25_port, CK => CLOCK, 
                           Q => addends_5_25_port, QN => n_1278);
   pipe1_reg_1_24_inst : DFF_X1 port map( D => mux_out_5_24_port, CK => CLOCK, 
                           Q => pipe1_1_24_port, QN => n_1279);
   addends_reg_5_24_inst : DFF_X1 port map( D => pipe1_1_24_port, CK => CLOCK, 
                           Q => addends_5_24_port, QN => n_1280);
   pipe1_reg_1_23_inst : DFF_X1 port map( D => mux_out_5_23_port, CK => CLOCK, 
                           Q => pipe1_1_23_port, QN => n_1281);
   addends_reg_5_23_inst : DFF_X1 port map( D => pipe1_1_23_port, CK => CLOCK, 
                           Q => addends_5_23_port, QN => n_1282);
   pipe1_reg_1_22_inst : DFF_X1 port map( D => mux_out_5_22_port, CK => CLOCK, 
                           Q => pipe1_1_22_port, QN => n_1283);
   addends_reg_5_22_inst : DFF_X1 port map( D => pipe1_1_22_port, CK => CLOCK, 
                           Q => addends_5_22_port, QN => n_1284);
   pipe1_reg_1_21_inst : DFF_X1 port map( D => mux_out_5_21_port, CK => CLOCK, 
                           Q => pipe1_1_21_port, QN => n_1285);
   addends_reg_5_21_inst : DFF_X1 port map( D => pipe1_1_21_port, CK => CLOCK, 
                           Q => addends_5_21_port, QN => n_1286);
   pipe1_reg_1_20_inst : DFF_X1 port map( D => mux_out_5_20_port, CK => CLOCK, 
                           Q => pipe1_1_20_port, QN => n_1287);
   addends_reg_5_20_inst : DFF_X1 port map( D => pipe1_1_20_port, CK => CLOCK, 
                           Q => addends_5_20_port, QN => n_1288);
   pipe1_reg_1_19_inst : DFF_X1 port map( D => mux_out_5_19_port, CK => CLOCK, 
                           Q => pipe1_1_19_port, QN => n_1289);
   addends_reg_5_19_inst : DFF_X1 port map( D => pipe1_1_19_port, CK => CLOCK, 
                           Q => addends_5_19_port, QN => n_1290);
   pipe1_reg_1_18_inst : DFF_X1 port map( D => mux_out_5_18_port, CK => CLOCK, 
                           Q => pipe1_1_18_port, QN => n_1291);
   addends_reg_5_18_inst : DFF_X1 port map( D => pipe1_1_18_port, CK => CLOCK, 
                           Q => addends_5_18_port, QN => n_1292);
   pipe1_reg_1_17_inst : DFF_X1 port map( D => mux_out_5_17_port, CK => CLOCK, 
                           Q => pipe1_1_17_port, QN => n_1293);
   addends_reg_5_17_inst : DFF_X1 port map( D => pipe1_1_17_port, CK => CLOCK, 
                           Q => addends_5_17_port, QN => n_1294);
   pipe1_reg_1_16_inst : DFF_X1 port map( D => mux_out_5_16_port, CK => CLOCK, 
                           Q => pipe1_1_16_port, QN => n_1295);
   addends_reg_5_16_inst : DFF_X1 port map( D => pipe1_1_16_port, CK => CLOCK, 
                           Q => addends_5_16_port, QN => n_1296);
   pipe1_reg_1_15_inst : DFF_X1 port map( D => mux_out_5_15_port, CK => CLOCK, 
                           Q => pipe1_1_15_port, QN => n_1297);
   addends_reg_5_15_inst : DFF_X1 port map( D => pipe1_1_15_port, CK => CLOCK, 
                           Q => addends_5_15_port, QN => n_1298);
   pipe1_reg_1_14_inst : DFF_X1 port map( D => mux_out_5_14_port, CK => CLOCK, 
                           Q => pipe1_1_14_port, QN => n_1299);
   addends_reg_5_14_inst : DFF_X1 port map( D => pipe1_1_14_port, CK => CLOCK, 
                           Q => addends_5_14_port, QN => n_1300);
   pipe1_reg_1_13_inst : DFF_X1 port map( D => mux_out_5_13_port, CK => CLOCK, 
                           Q => pipe1_1_13_port, QN => n_1301);
   addends_reg_5_13_inst : DFF_X1 port map( D => pipe1_1_13_port, CK => CLOCK, 
                           Q => addends_5_13_port, QN => n_1302);
   pipe1_reg_1_12_inst : DFF_X1 port map( D => mux_out_5_12_port, CK => CLOCK, 
                           Q => pipe1_1_12_port, QN => n_1303);
   addends_reg_5_12_inst : DFF_X1 port map( D => pipe1_1_12_port, CK => CLOCK, 
                           Q => addends_5_12_port, QN => n_1304);
   pipe1_reg_1_11_inst : DFF_X1 port map( D => mux_out_5_11_port, CK => CLOCK, 
                           Q => pipe1_1_11_port, QN => n_1305);
   addends_reg_5_11_inst : DFF_X1 port map( D => pipe1_1_11_port, CK => CLOCK, 
                           Q => addends_5_11_port, QN => n_1306);
   pipe1_reg_1_10_inst : DFF_X1 port map( D => mux_out_5_10_port, CK => CLOCK, 
                           Q => pipe1_1_10_port, QN => n_1307);
   addends_reg_5_10_inst : DFF_X1 port map( D => pipe1_1_10_port, CK => CLOCK, 
                           Q => addends_5_10_port, QN => n_1308);
   pipe1_reg_1_9_inst : DFF_X1 port map( D => mux_out_5_9_port, CK => CLOCK, Q 
                           => pipe1_1_9_port, QN => n_1309);
   addends_reg_5_9_inst : DFF_X1 port map( D => pipe1_1_9_port, CK => CLOCK, Q 
                           => addends_5_9_port, QN => n_1310);
   pipe1_reg_1_8_inst : DFF_X1 port map( D => mux_out_5_8_port, CK => CLOCK, Q 
                           => pipe1_1_8_port, QN => n_1311);
   addends_reg_5_8_inst : DFF_X1 port map( D => pipe1_1_8_port, CK => CLOCK, Q 
                           => addends_5_8_port, QN => n_1312);
   pipe1_reg_1_7_inst : DFF_X1 port map( D => mux_out_5_7_port, CK => CLOCK, Q 
                           => pipe1_1_7_port, QN => n_1313);
   addends_reg_5_7_inst : DFF_X1 port map( D => pipe1_1_7_port, CK => CLOCK, Q 
                           => addends_5_7_port, QN => n_1314);
   pipe1_reg_1_6_inst : DFF_X1 port map( D => mux_out_5_6_port, CK => CLOCK, Q 
                           => pipe1_1_6_port, QN => n_1315);
   addends_reg_5_6_inst : DFF_X1 port map( D => pipe1_1_6_port, CK => CLOCK, Q 
                           => addends_5_6_port, QN => n_1316);
   pipe1_reg_1_5_inst : DFF_X1 port map( D => mux_out_5_5_port, CK => CLOCK, Q 
                           => pipe1_1_5_port, QN => n_1317);
   addends_reg_5_5_inst : DFF_X1 port map( D => pipe1_1_5_port, CK => CLOCK, Q 
                           => addends_5_5_port, QN => n_1318);
   pipe1_reg_1_4_inst : DFF_X1 port map( D => mux_out_5_4_port, CK => CLOCK, Q 
                           => pipe1_1_4_port, QN => n_1319);
   addends_reg_5_4_inst : DFF_X1 port map( D => pipe1_1_4_port, CK => CLOCK, Q 
                           => addends_5_4_port, QN => n_1320);
   pipe1_reg_1_3_inst : DFF_X1 port map( D => mux_out_5_3_port, CK => CLOCK, Q 
                           => pipe1_1_3_port, QN => n_1321);
   addends_reg_5_3_inst : DFF_X1 port map( D => pipe1_1_3_port, CK => CLOCK, Q 
                           => addends_5_3_port, QN => n_1322);
   pipe1_reg_1_2_inst : DFF_X1 port map( D => mux_out_5_2_port, CK => CLOCK, Q 
                           => pipe1_1_2_port, QN => n_1323);
   addends_reg_5_2_inst : DFF_X1 port map( D => pipe1_1_2_port, CK => CLOCK, Q 
                           => addends_5_2_port, QN => n_1324);
   pipe1_reg_1_1_inst : DFF_X1 port map( D => mux_out_5_1_port, CK => CLOCK, Q 
                           => pipe1_1_1_port, QN => n_1325);
   addends_reg_5_1_inst : DFF_X1 port map( D => pipe1_1_1_port, CK => CLOCK, Q 
                           => addends_5_1_port, QN => n_1326);
   pipe1_reg_1_0_inst : DFF_X1 port map( D => mux_out_5_0_port, CK => CLOCK, Q 
                           => pipe1_1_0_port, QN => n_1327);
   addends_reg_5_0_inst : DFF_X1 port map( D => pipe1_1_0_port, CK => CLOCK, Q 
                           => addends_5_0_port, QN => n_1328);
   pipe1_reg_0_31_inst : DFF_X1 port map( D => mux_out_4_31_port, CK => CLOCK, 
                           Q => pipe1_0_31_port, QN => n_1329);
   addends_reg_4_31_inst : DFF_X1 port map( D => pipe1_0_31_port, CK => CLOCK, 
                           Q => addends_4_31_port, QN => n_1330);
   pipe1_reg_0_30_inst : DFF_X1 port map( D => mux_out_4_30_port, CK => CLOCK, 
                           Q => pipe1_0_30_port, QN => n_1331);
   addends_reg_4_30_inst : DFF_X1 port map( D => pipe1_0_30_port, CK => CLOCK, 
                           Q => addends_4_30_port, QN => n_1332);
   pipe1_reg_0_29_inst : DFF_X1 port map( D => mux_out_4_29_port, CK => CLOCK, 
                           Q => pipe1_0_29_port, QN => n_1333);
   addends_reg_4_29_inst : DFF_X1 port map( D => pipe1_0_29_port, CK => CLOCK, 
                           Q => addends_4_29_port, QN => n_1334);
   pipe1_reg_0_28_inst : DFF_X1 port map( D => mux_out_4_28_port, CK => CLOCK, 
                           Q => pipe1_0_28_port, QN => n_1335);
   addends_reg_4_28_inst : DFF_X1 port map( D => pipe1_0_28_port, CK => CLOCK, 
                           Q => addends_4_28_port, QN => n_1336);
   pipe1_reg_0_27_inst : DFF_X1 port map( D => mux_out_4_27_port, CK => CLOCK, 
                           Q => pipe1_0_27_port, QN => n_1337);
   addends_reg_4_27_inst : DFF_X1 port map( D => pipe1_0_27_port, CK => CLOCK, 
                           Q => addends_4_27_port, QN => n_1338);
   pipe1_reg_0_26_inst : DFF_X1 port map( D => mux_out_4_26_port, CK => CLOCK, 
                           Q => pipe1_0_26_port, QN => n_1339);
   addends_reg_4_26_inst : DFF_X1 port map( D => pipe1_0_26_port, CK => CLOCK, 
                           Q => addends_4_26_port, QN => n_1340);
   pipe1_reg_0_25_inst : DFF_X1 port map( D => mux_out_4_25_port, CK => CLOCK, 
                           Q => pipe1_0_25_port, QN => n_1341);
   addends_reg_4_25_inst : DFF_X1 port map( D => pipe1_0_25_port, CK => CLOCK, 
                           Q => addends_4_25_port, QN => n_1342);
   pipe1_reg_0_24_inst : DFF_X1 port map( D => mux_out_4_24_port, CK => CLOCK, 
                           Q => pipe1_0_24_port, QN => n_1343);
   addends_reg_4_24_inst : DFF_X1 port map( D => pipe1_0_24_port, CK => CLOCK, 
                           Q => addends_4_24_port, QN => n_1344);
   pipe1_reg_0_23_inst : DFF_X1 port map( D => mux_out_4_23_port, CK => CLOCK, 
                           Q => pipe1_0_23_port, QN => n_1345);
   addends_reg_4_23_inst : DFF_X1 port map( D => pipe1_0_23_port, CK => CLOCK, 
                           Q => addends_4_23_port, QN => n_1346);
   pipe1_reg_0_22_inst : DFF_X1 port map( D => mux_out_4_22_port, CK => CLOCK, 
                           Q => pipe1_0_22_port, QN => n_1347);
   addends_reg_4_22_inst : DFF_X1 port map( D => pipe1_0_22_port, CK => CLOCK, 
                           Q => addends_4_22_port, QN => n_1348);
   pipe1_reg_0_21_inst : DFF_X1 port map( D => mux_out_4_21_port, CK => CLOCK, 
                           Q => pipe1_0_21_port, QN => n_1349);
   addends_reg_4_21_inst : DFF_X1 port map( D => pipe1_0_21_port, CK => CLOCK, 
                           Q => addends_4_21_port, QN => n_1350);
   pipe1_reg_0_20_inst : DFF_X1 port map( D => mux_out_4_20_port, CK => CLOCK, 
                           Q => pipe1_0_20_port, QN => n_1351);
   addends_reg_4_20_inst : DFF_X1 port map( D => pipe1_0_20_port, CK => CLOCK, 
                           Q => addends_4_20_port, QN => n_1352);
   pipe1_reg_0_19_inst : DFF_X1 port map( D => mux_out_4_19_port, CK => CLOCK, 
                           Q => pipe1_0_19_port, QN => n_1353);
   addends_reg_4_19_inst : DFF_X1 port map( D => pipe1_0_19_port, CK => CLOCK, 
                           Q => addends_4_19_port, QN => n_1354);
   pipe1_reg_0_18_inst : DFF_X1 port map( D => mux_out_4_18_port, CK => CLOCK, 
                           Q => pipe1_0_18_port, QN => n_1355);
   addends_reg_4_18_inst : DFF_X1 port map( D => pipe1_0_18_port, CK => CLOCK, 
                           Q => addends_4_18_port, QN => n_1356);
   pipe1_reg_0_17_inst : DFF_X1 port map( D => mux_out_4_17_port, CK => CLOCK, 
                           Q => pipe1_0_17_port, QN => n_1357);
   addends_reg_4_17_inst : DFF_X1 port map( D => pipe1_0_17_port, CK => CLOCK, 
                           Q => addends_4_17_port, QN => n_1358);
   pipe1_reg_0_16_inst : DFF_X1 port map( D => mux_out_4_16_port, CK => CLOCK, 
                           Q => pipe1_0_16_port, QN => n_1359);
   addends_reg_4_16_inst : DFF_X1 port map( D => pipe1_0_16_port, CK => CLOCK, 
                           Q => addends_4_16_port, QN => n_1360);
   pipe1_reg_0_15_inst : DFF_X1 port map( D => mux_out_4_15_port, CK => CLOCK, 
                           Q => pipe1_0_15_port, QN => n_1361);
   addends_reg_4_15_inst : DFF_X1 port map( D => pipe1_0_15_port, CK => CLOCK, 
                           Q => addends_4_15_port, QN => n_1362);
   pipe1_reg_0_14_inst : DFF_X1 port map( D => mux_out_4_14_port, CK => CLOCK, 
                           Q => pipe1_0_14_port, QN => n_1363);
   addends_reg_4_14_inst : DFF_X1 port map( D => pipe1_0_14_port, CK => CLOCK, 
                           Q => addends_4_14_port, QN => n_1364);
   pipe1_reg_0_13_inst : DFF_X1 port map( D => mux_out_4_13_port, CK => CLOCK, 
                           Q => pipe1_0_13_port, QN => n_1365);
   addends_reg_4_13_inst : DFF_X1 port map( D => pipe1_0_13_port, CK => CLOCK, 
                           Q => addends_4_13_port, QN => n_1366);
   pipe1_reg_0_12_inst : DFF_X1 port map( D => mux_out_4_12_port, CK => CLOCK, 
                           Q => pipe1_0_12_port, QN => n_1367);
   addends_reg_4_12_inst : DFF_X1 port map( D => pipe1_0_12_port, CK => CLOCK, 
                           Q => addends_4_12_port, QN => n_1368);
   pipe1_reg_0_11_inst : DFF_X1 port map( D => mux_out_4_11_port, CK => CLOCK, 
                           Q => pipe1_0_11_port, QN => n_1369);
   addends_reg_4_11_inst : DFF_X1 port map( D => pipe1_0_11_port, CK => CLOCK, 
                           Q => addends_4_11_port, QN => n_1370);
   pipe1_reg_0_10_inst : DFF_X1 port map( D => mux_out_4_10_port, CK => CLOCK, 
                           Q => pipe1_0_10_port, QN => n_1371);
   addends_reg_4_10_inst : DFF_X1 port map( D => pipe1_0_10_port, CK => CLOCK, 
                           Q => addends_4_10_port, QN => n_1372);
   pipe1_reg_0_9_inst : DFF_X1 port map( D => mux_out_4_9_port, CK => CLOCK, Q 
                           => pipe1_0_9_port, QN => n_1373);
   addends_reg_4_9_inst : DFF_X1 port map( D => pipe1_0_9_port, CK => CLOCK, Q 
                           => addends_4_9_port, QN => n_1374);
   pipe1_reg_0_8_inst : DFF_X1 port map( D => mux_out_4_8_port, CK => CLOCK, Q 
                           => pipe1_0_8_port, QN => n_1375);
   addends_reg_4_8_inst : DFF_X1 port map( D => pipe1_0_8_port, CK => CLOCK, Q 
                           => addends_4_8_port, QN => n_1376);
   pipe1_reg_0_7_inst : DFF_X1 port map( D => mux_out_4_7_port, CK => CLOCK, Q 
                           => pipe1_0_7_port, QN => n_1377);
   addends_reg_4_7_inst : DFF_X1 port map( D => pipe1_0_7_port, CK => CLOCK, Q 
                           => addends_4_7_port, QN => n_1378);
   pipe1_reg_0_6_inst : DFF_X1 port map( D => mux_out_4_6_port, CK => CLOCK, Q 
                           => pipe1_0_6_port, QN => n_1379);
   addends_reg_4_6_inst : DFF_X1 port map( D => pipe1_0_6_port, CK => CLOCK, Q 
                           => addends_4_6_port, QN => n_1380);
   pipe1_reg_0_5_inst : DFF_X1 port map( D => mux_out_4_5_port, CK => CLOCK, Q 
                           => pipe1_0_5_port, QN => n_1381);
   addends_reg_4_5_inst : DFF_X1 port map( D => pipe1_0_5_port, CK => CLOCK, Q 
                           => addends_4_5_port, QN => n_1382);
   pipe1_reg_0_4_inst : DFF_X1 port map( D => mux_out_4_4_port, CK => CLOCK, Q 
                           => pipe1_0_4_port, QN => n_1383);
   addends_reg_4_4_inst : DFF_X1 port map( D => pipe1_0_4_port, CK => CLOCK, Q 
                           => addends_4_4_port, QN => n_1384);
   pipe1_reg_0_3_inst : DFF_X1 port map( D => mux_out_4_3_port, CK => CLOCK, Q 
                           => pipe1_0_3_port, QN => n_1385);
   addends_reg_4_3_inst : DFF_X1 port map( D => pipe1_0_3_port, CK => CLOCK, Q 
                           => addends_4_3_port, QN => n_1386);
   pipe1_reg_0_2_inst : DFF_X1 port map( D => mux_out_4_2_port, CK => CLOCK, Q 
                           => pipe1_0_2_port, QN => n_1387);
   addends_reg_4_2_inst : DFF_X1 port map( D => pipe1_0_2_port, CK => CLOCK, Q 
                           => addends_4_2_port, QN => n_1388);
   pipe1_reg_0_1_inst : DFF_X1 port map( D => mux_out_4_1_port, CK => CLOCK, Q 
                           => pipe1_0_1_port, QN => n_1389);
   addends_reg_4_1_inst : DFF_X1 port map( D => pipe1_0_1_port, CK => CLOCK, Q 
                           => addends_4_1_port, QN => n_1390);
   pipe1_reg_0_0_inst : DFF_X1 port map( D => mux_out_4_0_port, CK => CLOCK, Q 
                           => pipe1_0_0_port, QN => n_1391);
   pipe2_reg_1_31_inst : DFF_X1 port map( D => pipe1_3_31_port, CK => CLOCK, Q 
                           => pipe2_1_31_port, QN => n_1392);
   addends_reg_7_31_inst : DFF_X1 port map( D => pipe2_1_31_port, CK => CLOCK, 
                           Q => addends_7_31_port, QN => n_1393);
   pipe2_reg_1_30_inst : DFF_X1 port map( D => pipe1_3_30_port, CK => CLOCK, Q 
                           => pipe2_1_30_port, QN => n_1394);
   addends_reg_7_30_inst : DFF_X1 port map( D => pipe2_1_30_port, CK => CLOCK, 
                           Q => addends_7_30_port, QN => n_1395);
   pipe2_reg_1_29_inst : DFF_X1 port map( D => pipe1_3_29_port, CK => CLOCK, Q 
                           => pipe2_1_29_port, QN => n_1396);
   addends_reg_7_29_inst : DFF_X1 port map( D => pipe2_1_29_port, CK => CLOCK, 
                           Q => addends_7_29_port, QN => n_1397);
   pipe2_reg_1_28_inst : DFF_X1 port map( D => pipe1_3_28_port, CK => CLOCK, Q 
                           => pipe2_1_28_port, QN => n_1398);
   addends_reg_7_28_inst : DFF_X1 port map( D => pipe2_1_28_port, CK => CLOCK, 
                           Q => addends_7_28_port, QN => n_1399);
   pipe2_reg_1_27_inst : DFF_X1 port map( D => pipe1_3_27_port, CK => CLOCK, Q 
                           => pipe2_1_27_port, QN => n_1400);
   addends_reg_7_27_inst : DFF_X1 port map( D => pipe2_1_27_port, CK => CLOCK, 
                           Q => addends_7_27_port, QN => n_1401);
   pipe2_reg_1_26_inst : DFF_X1 port map( D => pipe1_3_26_port, CK => CLOCK, Q 
                           => pipe2_1_26_port, QN => n_1402);
   addends_reg_7_26_inst : DFF_X1 port map( D => pipe2_1_26_port, CK => CLOCK, 
                           Q => addends_7_26_port, QN => n_1403);
   pipe2_reg_1_25_inst : DFF_X1 port map( D => pipe1_3_25_port, CK => CLOCK, Q 
                           => pipe2_1_25_port, QN => n_1404);
   addends_reg_7_25_inst : DFF_X1 port map( D => pipe2_1_25_port, CK => CLOCK, 
                           Q => addends_7_25_port, QN => n_1405);
   pipe2_reg_1_24_inst : DFF_X1 port map( D => pipe1_3_24_port, CK => CLOCK, Q 
                           => pipe2_1_24_port, QN => n_1406);
   addends_reg_7_24_inst : DFF_X1 port map( D => pipe2_1_24_port, CK => CLOCK, 
                           Q => addends_7_24_port, QN => n_1407);
   pipe2_reg_1_23_inst : DFF_X1 port map( D => pipe1_3_23_port, CK => CLOCK, Q 
                           => pipe2_1_23_port, QN => n_1408);
   addends_reg_7_23_inst : DFF_X1 port map( D => pipe2_1_23_port, CK => CLOCK, 
                           Q => addends_7_23_port, QN => n_1409);
   pipe2_reg_1_22_inst : DFF_X1 port map( D => pipe1_3_22_port, CK => CLOCK, Q 
                           => pipe2_1_22_port, QN => n_1410);
   addends_reg_7_22_inst : DFF_X1 port map( D => pipe2_1_22_port, CK => CLOCK, 
                           Q => addends_7_22_port, QN => n_1411);
   pipe2_reg_1_21_inst : DFF_X1 port map( D => pipe1_3_21_port, CK => CLOCK, Q 
                           => pipe2_1_21_port, QN => n_1412);
   addends_reg_7_21_inst : DFF_X1 port map( D => pipe2_1_21_port, CK => CLOCK, 
                           Q => addends_7_21_port, QN => n_1413);
   pipe2_reg_1_20_inst : DFF_X1 port map( D => pipe1_3_20_port, CK => CLOCK, Q 
                           => pipe2_1_20_port, QN => n_1414);
   addends_reg_7_20_inst : DFF_X1 port map( D => pipe2_1_20_port, CK => CLOCK, 
                           Q => addends_7_20_port, QN => n_1415);
   pipe2_reg_1_19_inst : DFF_X1 port map( D => pipe1_3_19_port, CK => CLOCK, Q 
                           => pipe2_1_19_port, QN => n_1416);
   addends_reg_7_19_inst : DFF_X1 port map( D => pipe2_1_19_port, CK => CLOCK, 
                           Q => addends_7_19_port, QN => n_1417);
   pipe2_reg_1_18_inst : DFF_X1 port map( D => pipe1_3_18_port, CK => CLOCK, Q 
                           => pipe2_1_18_port, QN => n_1418);
   addends_reg_7_18_inst : DFF_X1 port map( D => pipe2_1_18_port, CK => CLOCK, 
                           Q => addends_7_18_port, QN => n_1419);
   pipe2_reg_1_17_inst : DFF_X1 port map( D => pipe1_3_17_port, CK => CLOCK, Q 
                           => pipe2_1_17_port, QN => n_1420);
   addends_reg_7_17_inst : DFF_X1 port map( D => pipe2_1_17_port, CK => CLOCK, 
                           Q => addends_7_17_port, QN => n_1421);
   pipe2_reg_1_16_inst : DFF_X1 port map( D => pipe1_3_16_port, CK => CLOCK, Q 
                           => pipe2_1_16_port, QN => n_1422);
   addends_reg_7_16_inst : DFF_X1 port map( D => pipe2_1_16_port, CK => CLOCK, 
                           Q => addends_7_16_port, QN => n_1423);
   pipe2_reg_1_15_inst : DFF_X1 port map( D => pipe1_3_15_port, CK => CLOCK, Q 
                           => pipe2_1_15_port, QN => n_1424);
   addends_reg_7_15_inst : DFF_X1 port map( D => pipe2_1_15_port, CK => CLOCK, 
                           Q => addends_7_15_port, QN => n_1425);
   pipe2_reg_1_14_inst : DFF_X1 port map( D => pipe1_3_14_port, CK => CLOCK, Q 
                           => pipe2_1_14_port, QN => n_1426);
   addends_reg_7_14_inst : DFF_X1 port map( D => pipe2_1_14_port, CK => CLOCK, 
                           Q => addends_7_14_port, QN => n_1427);
   pipe2_reg_1_13_inst : DFF_X1 port map( D => pipe1_3_13_port, CK => CLOCK, Q 
                           => pipe2_1_13_port, QN => n_1428);
   addends_reg_7_13_inst : DFF_X1 port map( D => pipe2_1_13_port, CK => CLOCK, 
                           Q => addends_7_13_port, QN => n_1429);
   pipe2_reg_1_12_inst : DFF_X1 port map( D => pipe1_3_12_port, CK => CLOCK, Q 
                           => pipe2_1_12_port, QN => n_1430);
   addends_reg_7_12_inst : DFF_X1 port map( D => pipe2_1_12_port, CK => CLOCK, 
                           Q => addends_7_12_port, QN => n_1431);
   pipe2_reg_1_11_inst : DFF_X1 port map( D => pipe1_3_11_port, CK => CLOCK, Q 
                           => pipe2_1_11_port, QN => n_1432);
   addends_reg_7_11_inst : DFF_X1 port map( D => pipe2_1_11_port, CK => CLOCK, 
                           Q => addends_7_11_port, QN => n_1433);
   pipe2_reg_1_10_inst : DFF_X1 port map( D => pipe1_3_10_port, CK => CLOCK, Q 
                           => pipe2_1_10_port, QN => n_1434);
   addends_reg_7_10_inst : DFF_X1 port map( D => pipe2_1_10_port, CK => CLOCK, 
                           Q => addends_7_10_port, QN => n_1435);
   pipe2_reg_1_9_inst : DFF_X1 port map( D => pipe1_3_9_port, CK => CLOCK, Q =>
                           pipe2_1_9_port, QN => n_1436);
   addends_reg_7_9_inst : DFF_X1 port map( D => pipe2_1_9_port, CK => CLOCK, Q 
                           => addends_7_9_port, QN => n_1437);
   pipe2_reg_1_8_inst : DFF_X1 port map( D => pipe1_3_8_port, CK => CLOCK, Q =>
                           pipe2_1_8_port, QN => n_1438);
   addends_reg_7_8_inst : DFF_X1 port map( D => pipe2_1_8_port, CK => CLOCK, Q 
                           => addends_7_8_port, QN => n_1439);
   pipe2_reg_1_7_inst : DFF_X1 port map( D => pipe1_3_7_port, CK => CLOCK, Q =>
                           pipe2_1_7_port, QN => n_1440);
   addends_reg_7_7_inst : DFF_X1 port map( D => pipe2_1_7_port, CK => CLOCK, Q 
                           => addends_7_7_port, QN => n_1441);
   pipe2_reg_1_6_inst : DFF_X1 port map( D => pipe1_3_6_port, CK => CLOCK, Q =>
                           pipe2_1_6_port, QN => n_1442);
   addends_reg_7_6_inst : DFF_X1 port map( D => pipe2_1_6_port, CK => CLOCK, Q 
                           => addends_7_6_port, QN => n_1443);
   pipe2_reg_1_5_inst : DFF_X1 port map( D => pipe1_3_5_port, CK => CLOCK, Q =>
                           pipe2_1_5_port, QN => n_1444);
   addends_reg_7_5_inst : DFF_X1 port map( D => pipe2_1_5_port, CK => CLOCK, Q 
                           => addends_7_5_port, QN => n_1445);
   pipe2_reg_1_4_inst : DFF_X1 port map( D => pipe1_3_4_port, CK => CLOCK, Q =>
                           pipe2_1_4_port, QN => n_1446);
   addends_reg_7_4_inst : DFF_X1 port map( D => pipe2_1_4_port, CK => CLOCK, Q 
                           => addends_7_4_port, QN => n_1447);
   pipe2_reg_1_3_inst : DFF_X1 port map( D => pipe1_3_3_port, CK => CLOCK, Q =>
                           pipe2_1_3_port, QN => n_1448);
   addends_reg_7_3_inst : DFF_X1 port map( D => pipe2_1_3_port, CK => CLOCK, Q 
                           => addends_7_3_port, QN => n_1449);
   pipe2_reg_1_2_inst : DFF_X1 port map( D => pipe1_3_2_port, CK => CLOCK, Q =>
                           pipe2_1_2_port, QN => n_1450);
   addends_reg_7_2_inst : DFF_X1 port map( D => pipe2_1_2_port, CK => CLOCK, Q 
                           => addends_7_2_port, QN => n_1451);
   pipe2_reg_1_1_inst : DFF_X1 port map( D => pipe1_3_1_port, CK => CLOCK, Q =>
                           pipe2_1_1_port, QN => n_1452);
   addends_reg_7_1_inst : DFF_X1 port map( D => pipe2_1_1_port, CK => CLOCK, Q 
                           => addends_7_1_port, QN => n_1453);
   pipe2_reg_1_0_inst : DFF_X1 port map( D => pipe1_3_0_port, CK => CLOCK, Q =>
                           pipe2_1_0_port, QN => n_1454);
   addends_reg_7_0_inst : DFF_X1 port map( D => pipe2_1_0_port, CK => CLOCK, Q 
                           => addends_7_0_port, QN => n_1455);
   pipe2_reg_0_31_inst : DFF_X1 port map( D => pipe1_2_31_port, CK => CLOCK, Q 
                           => pipe2_0_31_port, QN => n_1456);
   addends_reg_6_31_inst : DFF_X1 port map( D => pipe2_0_31_port, CK => CLOCK, 
                           Q => addends_6_31_port, QN => n_1457);
   pipe2_reg_0_30_inst : DFF_X1 port map( D => pipe1_2_30_port, CK => CLOCK, Q 
                           => pipe2_0_30_port, QN => n_1458);
   addends_reg_6_30_inst : DFF_X1 port map( D => pipe2_0_30_port, CK => CLOCK, 
                           Q => addends_6_30_port, QN => n_1459);
   pipe2_reg_0_29_inst : DFF_X1 port map( D => pipe1_2_29_port, CK => CLOCK, Q 
                           => pipe2_0_29_port, QN => n_1460);
   addends_reg_6_29_inst : DFF_X1 port map( D => pipe2_0_29_port, CK => CLOCK, 
                           Q => addends_6_29_port, QN => n_1461);
   pipe2_reg_0_28_inst : DFF_X1 port map( D => pipe1_2_28_port, CK => CLOCK, Q 
                           => pipe2_0_28_port, QN => n_1462);
   addends_reg_6_28_inst : DFF_X1 port map( D => pipe2_0_28_port, CK => CLOCK, 
                           Q => addends_6_28_port, QN => n_1463);
   pipe2_reg_0_27_inst : DFF_X1 port map( D => pipe1_2_27_port, CK => CLOCK, Q 
                           => pipe2_0_27_port, QN => n_1464);
   addends_reg_6_27_inst : DFF_X1 port map( D => pipe2_0_27_port, CK => CLOCK, 
                           Q => addends_6_27_port, QN => n_1465);
   pipe2_reg_0_26_inst : DFF_X1 port map( D => pipe1_2_26_port, CK => CLOCK, Q 
                           => pipe2_0_26_port, QN => n_1466);
   addends_reg_6_26_inst : DFF_X1 port map( D => pipe2_0_26_port, CK => CLOCK, 
                           Q => addends_6_26_port, QN => n_1467);
   pipe2_reg_0_25_inst : DFF_X1 port map( D => pipe1_2_25_port, CK => CLOCK, Q 
                           => pipe2_0_25_port, QN => n_1468);
   addends_reg_6_25_inst : DFF_X1 port map( D => pipe2_0_25_port, CK => CLOCK, 
                           Q => addends_6_25_port, QN => n_1469);
   pipe2_reg_0_24_inst : DFF_X1 port map( D => pipe1_2_24_port, CK => CLOCK, Q 
                           => pipe2_0_24_port, QN => n_1470);
   addends_reg_6_24_inst : DFF_X1 port map( D => pipe2_0_24_port, CK => CLOCK, 
                           Q => addends_6_24_port, QN => n_1471);
   pipe2_reg_0_23_inst : DFF_X1 port map( D => pipe1_2_23_port, CK => CLOCK, Q 
                           => pipe2_0_23_port, QN => n_1472);
   addends_reg_6_23_inst : DFF_X1 port map( D => pipe2_0_23_port, CK => CLOCK, 
                           Q => addends_6_23_port, QN => n_1473);
   pipe2_reg_0_22_inst : DFF_X1 port map( D => pipe1_2_22_port, CK => CLOCK, Q 
                           => pipe2_0_22_port, QN => n_1474);
   addends_reg_6_22_inst : DFF_X1 port map( D => pipe2_0_22_port, CK => CLOCK, 
                           Q => addends_6_22_port, QN => n_1475);
   pipe2_reg_0_21_inst : DFF_X1 port map( D => pipe1_2_21_port, CK => CLOCK, Q 
                           => pipe2_0_21_port, QN => n_1476);
   addends_reg_6_21_inst : DFF_X1 port map( D => pipe2_0_21_port, CK => CLOCK, 
                           Q => addends_6_21_port, QN => n_1477);
   pipe2_reg_0_20_inst : DFF_X1 port map( D => pipe1_2_20_port, CK => CLOCK, Q 
                           => pipe2_0_20_port, QN => n_1478);
   addends_reg_6_20_inst : DFF_X1 port map( D => pipe2_0_20_port, CK => CLOCK, 
                           Q => addends_6_20_port, QN => n_1479);
   pipe2_reg_0_19_inst : DFF_X1 port map( D => pipe1_2_19_port, CK => CLOCK, Q 
                           => pipe2_0_19_port, QN => n_1480);
   addends_reg_6_19_inst : DFF_X1 port map( D => pipe2_0_19_port, CK => CLOCK, 
                           Q => addends_6_19_port, QN => n_1481);
   pipe2_reg_0_18_inst : DFF_X1 port map( D => pipe1_2_18_port, CK => CLOCK, Q 
                           => pipe2_0_18_port, QN => n_1482);
   addends_reg_6_18_inst : DFF_X1 port map( D => pipe2_0_18_port, CK => CLOCK, 
                           Q => addends_6_18_port, QN => n_1483);
   pipe2_reg_0_17_inst : DFF_X1 port map( D => pipe1_2_17_port, CK => CLOCK, Q 
                           => pipe2_0_17_port, QN => n_1484);
   addends_reg_6_17_inst : DFF_X1 port map( D => pipe2_0_17_port, CK => CLOCK, 
                           Q => addends_6_17_port, QN => n_1485);
   pipe2_reg_0_16_inst : DFF_X1 port map( D => pipe1_2_16_port, CK => CLOCK, Q 
                           => pipe2_0_16_port, QN => n_1486);
   addends_reg_6_16_inst : DFF_X1 port map( D => pipe2_0_16_port, CK => CLOCK, 
                           Q => addends_6_16_port, QN => n_1487);
   pipe2_reg_0_15_inst : DFF_X1 port map( D => pipe1_2_15_port, CK => CLOCK, Q 
                           => pipe2_0_15_port, QN => n_1488);
   addends_reg_6_15_inst : DFF_X1 port map( D => pipe2_0_15_port, CK => CLOCK, 
                           Q => addends_6_15_port, QN => n_1489);
   pipe2_reg_0_14_inst : DFF_X1 port map( D => pipe1_2_14_port, CK => CLOCK, Q 
                           => pipe2_0_14_port, QN => n_1490);
   addends_reg_6_14_inst : DFF_X1 port map( D => pipe2_0_14_port, CK => CLOCK, 
                           Q => addends_6_14_port, QN => n_1491);
   pipe2_reg_0_13_inst : DFF_X1 port map( D => pipe1_2_13_port, CK => CLOCK, Q 
                           => pipe2_0_13_port, QN => n_1492);
   addends_reg_6_13_inst : DFF_X1 port map( D => pipe2_0_13_port, CK => CLOCK, 
                           Q => addends_6_13_port, QN => n_1493);
   pipe2_reg_0_12_inst : DFF_X1 port map( D => pipe1_2_12_port, CK => CLOCK, Q 
                           => pipe2_0_12_port, QN => n_1494);
   addends_reg_6_12_inst : DFF_X1 port map( D => pipe2_0_12_port, CK => CLOCK, 
                           Q => addends_6_12_port, QN => n_1495);
   pipe2_reg_0_11_inst : DFF_X1 port map( D => pipe1_2_11_port, CK => CLOCK, Q 
                           => pipe2_0_11_port, QN => n_1496);
   addends_reg_6_11_inst : DFF_X1 port map( D => pipe2_0_11_port, CK => CLOCK, 
                           Q => addends_6_11_port, QN => n_1497);
   pipe2_reg_0_10_inst : DFF_X1 port map( D => pipe1_2_10_port, CK => CLOCK, Q 
                           => pipe2_0_10_port, QN => n_1498);
   addends_reg_6_10_inst : DFF_X1 port map( D => pipe2_0_10_port, CK => CLOCK, 
                           Q => addends_6_10_port, QN => n_1499);
   pipe2_reg_0_9_inst : DFF_X1 port map( D => pipe1_2_9_port, CK => CLOCK, Q =>
                           pipe2_0_9_port, QN => n_1500);
   addends_reg_6_9_inst : DFF_X1 port map( D => pipe2_0_9_port, CK => CLOCK, Q 
                           => addends_6_9_port, QN => n_1501);
   pipe2_reg_0_8_inst : DFF_X1 port map( D => pipe1_2_8_port, CK => CLOCK, Q =>
                           pipe2_0_8_port, QN => n_1502);
   addends_reg_6_8_inst : DFF_X1 port map( D => pipe2_0_8_port, CK => CLOCK, Q 
                           => addends_6_8_port, QN => n_1503);
   pipe2_reg_0_7_inst : DFF_X1 port map( D => pipe1_2_7_port, CK => CLOCK, Q =>
                           pipe2_0_7_port, QN => n_1504);
   addends_reg_6_7_inst : DFF_X1 port map( D => pipe2_0_7_port, CK => CLOCK, Q 
                           => addends_6_7_port, QN => n_1505);
   pipe2_reg_0_6_inst : DFF_X1 port map( D => pipe1_2_6_port, CK => CLOCK, Q =>
                           pipe2_0_6_port, QN => n_1506);
   addends_reg_6_6_inst : DFF_X1 port map( D => pipe2_0_6_port, CK => CLOCK, Q 
                           => addends_6_6_port, QN => n_1507);
   pipe2_reg_0_5_inst : DFF_X1 port map( D => pipe1_2_5_port, CK => CLOCK, Q =>
                           pipe2_0_5_port, QN => n_1508);
   addends_reg_6_5_inst : DFF_X1 port map( D => pipe2_0_5_port, CK => CLOCK, Q 
                           => addends_6_5_port, QN => n_1509);
   pipe2_reg_0_4_inst : DFF_X1 port map( D => pipe1_2_4_port, CK => CLOCK, Q =>
                           pipe2_0_4_port, QN => n_1510);
   addends_reg_6_4_inst : DFF_X1 port map( D => pipe2_0_4_port, CK => CLOCK, Q 
                           => addends_6_4_port, QN => n_1511);
   pipe2_reg_0_3_inst : DFF_X1 port map( D => pipe1_2_3_port, CK => CLOCK, Q =>
                           pipe2_0_3_port, QN => n_1512);
   pipe2_reg_0_2_inst : DFF_X1 port map( D => pipe1_2_2_port, CK => CLOCK, Q =>
                           pipe2_0_2_port, QN => n_1513);
   addends_reg_6_2_inst : DFF_X1 port map( D => pipe2_0_2_port, CK => CLOCK, Q 
                           => addends_6_2_port, QN => n_1514);
   pipe2_reg_0_1_inst : DFF_X1 port map( D => pipe1_2_1_port, CK => CLOCK, Q =>
                           pipe2_0_1_port, QN => n_1515);
   pipe2_reg_0_0_inst : DFF_X1 port map( D => pipe1_2_0_port, CK => CLOCK, Q =>
                           pipe2_0_0_port, QN => n_1516);
   addends_reg_6_1_inst : DFF_X1 port map( D => pipe2_0_1_port, CK => CLOCK, Q 
                           => addends_6_1_port, QN => n_1517);
   addends_reg_6_0_inst : DFF_X1 port map( D => pipe2_0_0_port, CK => CLOCK, Q 
                           => addends_6_0_port, QN => n_1518);
   addends_reg_4_0_inst : DFF_X1 port map( D => pipe1_0_0_port, CK => CLOCK, Q 
                           => addends_4_0_port, QN => n_1519);
   addends_reg_6_3_inst : DFF_X1 port map( D => pipe2_0_3_port, CK => CLOCK, Q 
                           => addends_6_3_port, QN => n_1520);
   n69 <= '0';
   U5 : XNOR2_X2 port map( A => n10, B => A(5), ZN => A_neg_9_14_port);
   U8 : XNOR2_X2 port map( A => n4, B => A(15), ZN => A_neg_9_24_port);
   enc_1 : ENCODER_0 port map( INPUT(2) => B(1), INPUT(1) => B(0), INPUT(0) => 
                           X_Logic0_port, OUTPUT(2) => selector_2_port, 
                           OUTPUT(1) => selector_1_port, OUTPUT(0) => 
                           selector_0_port);
   enc_2 : ENCODER_7 port map( INPUT(2) => B(3), INPUT(1) => B(2), INPUT(0) => 
                           B(1), OUTPUT(2) => selector_5_port, OUTPUT(1) => 
                           selector_4_port, OUTPUT(0) => selector_3_port);
   enc_3 : ENCODER_6 port map( INPUT(2) => B(5), INPUT(1) => B(4), INPUT(0) => 
                           B(3), OUTPUT(2) => selector_8_port, OUTPUT(1) => 
                           selector_7_port, OUTPUT(0) => selector_6_port);
   enc_4 : ENCODER_5 port map( INPUT(2) => B(7), INPUT(1) => B(6), INPUT(0) => 
                           B(5), OUTPUT(2) => selector_11_port, OUTPUT(1) => 
                           selector_10_port, OUTPUT(0) => selector_9_port);
   enc_5 : ENCODER_4 port map( INPUT(2) => B(9), INPUT(1) => B(8), INPUT(0) => 
                           B(7), OUTPUT(2) => selector_14_port, OUTPUT(1) => 
                           selector_13_port, OUTPUT(0) => selector_12_port);
   enc_6 : ENCODER_3 port map( INPUT(2) => B(11), INPUT(1) => B(10), INPUT(0) 
                           => B(9), OUTPUT(2) => selector_17_port, OUTPUT(1) =>
                           selector_16_port, OUTPUT(0) => selector_15_port);
   enc_7 : ENCODER_2 port map( INPUT(2) => B(13), INPUT(1) => B(12), INPUT(0) 
                           => B(11), OUTPUT(2) => selector_20_port, OUTPUT(1) 
                           => selector_19_port, OUTPUT(0) => selector_18_port);
   enc_8 : ENCODER_1 port map( INPUT(2) => B(15), INPUT(1) => B(14), INPUT(0) 
                           => B(13), OUTPUT(2) => selector_23_port, OUTPUT(1) 
                           => selector_22_port, OUTPUT(0) => selector_21_port);
   MUX_I_0 : MUX5to1_NBIT32_8 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => A(15), B(14) => A(14), B(13)
                           => A(13), B(12) => A(12), B(11) => A(11), B(10) => 
                           A(10), B(9) => A(9), B(8) => A(8), B(7) => A(7), 
                           B(6) => A(6), B(5) => A(5), B(4) => A(4), B(3) => 
                           A(3), B(2) => A(2), B(1) => A(1), B(0) => n96, C(31)
                           => n82, C(30) => n78, C(29) => n78, C(28) => n78, 
                           C(27) => n78, C(26) => n78, C(25) => n78, C(24) => 
                           n78, C(23) => n78, C(22) => n78, C(21) => n78, C(20)
                           => n78, C(19) => n78, C(18) => n79, C(17) => n79, 
                           C(16) => n79, C(15) => A_neg_9_24_port, C(14) => 
                           A_neg_9_23_port, C(13) => A_neg_9_22_port, C(12) => 
                           A_neg_9_21_port, C(11) => A_neg_9_20_port, C(10) => 
                           A_neg_9_19_port, C(9) => A_neg_9_18_port, C(8) => 
                           A_neg_9_17_port, C(7) => A_neg_9_16_port, C(6) => 
                           A_neg_9_15_port, C(5) => A_neg_9_14_port, C(4) => 
                           A_neg_9_13_port, C(3) => A_neg_9_12_port, C(2) => 
                           A_neg_9_11_port, C(1) => A_neg_9_10_port, C(0) => 
                           n95, D(31) => X_Logic0_port, D(30) => X_Logic0_port,
                           D(29) => X_Logic0_port, D(28) => X_Logic0_port, 
                           D(27) => X_Logic0_port, D(26) => X_Logic0_port, 
                           D(25) => X_Logic0_port, D(24) => X_Logic0_port, 
                           D(23) => X_Logic0_port, D(22) => X_Logic0_port, 
                           D(21) => X_Logic0_port, D(20) => X_Logic0_port, 
                           D(19) => X_Logic0_port, D(18) => X_Logic0_port, 
                           D(17) => X_Logic0_port, D(16) => A(15), D(15) => 
                           A(14), D(14) => A(13), D(13) => A(12), D(12) => 
                           A(11), D(11) => A(10), D(10) => A(9), D(9) => A(8), 
                           D(8) => A(7), D(7) => A(6), D(6) => A(5), D(5) => 
                           A(4), D(4) => A(3), D(3) => A(2), D(2) => A(1), D(1)
                           => n94, D(0) => X_Logic0_port, E(31) => n88, E(30) 
                           => n88, E(29) => n88, E(28) => n87, E(27) => n87, 
                           E(26) => n88, E(25) => n87, E(24) => n87, E(23) => 
                           n88, E(22) => n87, E(21) => n87, E(20) => n88, E(19)
                           => n88, E(18) => n87, E(17) => n87, E(16) => 
                           A_neg_9_24_port, E(15) => A_neg_9_23_port, E(14) => 
                           A_neg_9_22_port, E(13) => A_neg_9_21_port, E(12) => 
                           A_neg_9_20_port, E(11) => A_neg_9_19_port, E(10) => 
                           A_neg_9_18_port, E(9) => A_neg_9_17_port, E(8) => 
                           A_neg_9_16_port, E(7) => A_neg_9_15_port, E(6) => 
                           A_neg_9_14_port, E(5) => A_neg_9_13_port, E(4) => 
                           A_neg_9_12_port, E(3) => A_neg_9_11_port, E(2) => 
                           A_neg_9_10_port, E(1) => n95, E(0) => n69, SEL(2) =>
                           selector_2_port, SEL(1) => selector_1_port, SEL(0) 
                           => selector_0_port, Y(31) => addends_0_31_port, 
                           Y(30) => addends_0_30_port, Y(29) => 
                           addends_0_29_port, Y(28) => addends_0_28_port, Y(27)
                           => addends_0_27_port, Y(26) => addends_0_26_port, 
                           Y(25) => addends_0_25_port, Y(24) => 
                           addends_0_24_port, Y(23) => addends_0_23_port, Y(22)
                           => addends_0_22_port, Y(21) => addends_0_21_port, 
                           Y(20) => addends_0_20_port, Y(19) => 
                           addends_0_19_port, Y(18) => addends_0_18_port, Y(17)
                           => addends_0_17_port, Y(16) => addends_0_16_port, 
                           Y(15) => addends_0_15_port, Y(14) => 
                           addends_0_14_port, Y(13) => addends_0_13_port, Y(12)
                           => addends_0_12_port, Y(11) => addends_0_11_port, 
                           Y(10) => addends_0_10_port, Y(9) => addends_0_9_port
                           , Y(8) => addends_0_8_port, Y(7) => addends_0_7_port
                           , Y(6) => addends_0_6_port, Y(5) => addends_0_5_port
                           , Y(4) => addends_0_4_port, Y(3) => addends_0_3_port
                           , Y(2) => addends_0_2_port, Y(1) => addends_0_1_port
                           , Y(0) => addends_0_0_port);
   MUX_I_1 : MUX5to1_NBIT32_7 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => A(15), B(16) => A(14), B(15)
                           => A(13), B(14) => A(12), B(13) => A(11), B(12) => 
                           A(10), B(11) => A(9), B(10) => A(8), B(9) => A(7), 
                           B(8) => A(6), B(7) => A(5), B(6) => A(4), B(5) => 
                           A(3), B(4) => A(2), B(3) => A(1), B(2) => n96, B(1) 
                           => X_Logic0_port, B(0) => X_Logic0_port, C(31) => 
                           n79, C(30) => n79, C(29) => n79, C(28) => n79, C(27)
                           => n79, C(26) => n79, C(25) => n79, C(24) => n79, 
                           C(23) => n79, C(22) => n80, C(21) => n80, C(20) => 
                           n80, C(19) => n80, C(18) => n80, C(17) => 
                           A_neg_9_24_port, C(16) => A_neg_9_23_port, C(15) => 
                           A_neg_9_22_port, C(14) => A_neg_9_21_port, C(13) => 
                           A_neg_9_20_port, C(12) => A_neg_9_19_port, C(11) => 
                           A_neg_9_18_port, C(10) => A_neg_9_17_port, C(9) => 
                           A_neg_9_16_port, C(8) => A_neg_9_15_port, C(7) => 
                           A_neg_9_14_port, C(6) => A_neg_9_13_port, C(5) => 
                           A_neg_9_12_port, C(4) => A_neg_9_11_port, C(3) => 
                           A_neg_9_10_port, C(2) => n95, C(1) => n69, C(0) => 
                           n69, D(31) => X_Logic0_port, D(30) => X_Logic0_port,
                           D(29) => X_Logic0_port, D(28) => X_Logic0_port, 
                           D(27) => X_Logic0_port, D(26) => X_Logic0_port, 
                           D(25) => X_Logic0_port, D(24) => X_Logic0_port, 
                           D(23) => X_Logic0_port, D(22) => X_Logic0_port, 
                           D(21) => X_Logic0_port, D(20) => X_Logic0_port, 
                           D(19) => X_Logic0_port, D(18) => A(15), D(17) => 
                           A(14), D(16) => A(13), D(15) => A(12), D(14) => 
                           A(11), D(13) => A(10), D(12) => A(9), D(11) => A(8),
                           D(10) => A(7), D(9) => A(6), D(8) => A(5), D(7) => 
                           A(4), D(6) => A(3), D(5) => A(2), D(4) => A(1), D(3)
                           => n94, D(2) => X_Logic0_port, D(1) => X_Logic0_port
                           , D(0) => X_Logic0_port, E(31) => n86, E(30) => n86,
                           E(29) => n85, E(28) => n86, E(27) => n86, E(26) => 
                           n85, E(25) => n86, E(24) => n85, E(23) => n85, E(22)
                           => n86, E(21) => n85, E(20) => n87, E(19) => n86, 
                           E(18) => A_neg_9_24_port, E(17) => A_neg_9_23_port, 
                           E(16) => A_neg_9_22_port, E(15) => A_neg_9_21_port, 
                           E(14) => A_neg_9_20_port, E(13) => A_neg_9_19_port, 
                           E(12) => A_neg_9_18_port, E(11) => A_neg_9_17_port, 
                           E(10) => A_neg_9_16_port, E(9) => A_neg_9_15_port, 
                           E(8) => A_neg_9_14_port, E(7) => A_neg_9_13_port, 
                           E(6) => A_neg_9_12_port, E(5) => A_neg_9_11_port, 
                           E(4) => A_neg_9_10_port, E(3) => n95, E(2) => n69, 
                           E(1) => n69, E(0) => n69, SEL(2) => selector_5_port,
                           SEL(1) => selector_4_port, SEL(0) => selector_3_port
                           , Y(31) => addends_1_31_port, Y(30) => 
                           addends_1_30_port, Y(29) => addends_1_29_port, Y(28)
                           => addends_1_28_port, Y(27) => addends_1_27_port, 
                           Y(26) => addends_1_26_port, Y(25) => 
                           addends_1_25_port, Y(24) => addends_1_24_port, Y(23)
                           => addends_1_23_port, Y(22) => addends_1_22_port, 
                           Y(21) => addends_1_21_port, Y(20) => 
                           addends_1_20_port, Y(19) => addends_1_19_port, Y(18)
                           => addends_1_18_port, Y(17) => addends_1_17_port, 
                           Y(16) => addends_1_16_port, Y(15) => 
                           addends_1_15_port, Y(14) => addends_1_14_port, Y(13)
                           => addends_1_13_port, Y(12) => addends_1_12_port, 
                           Y(11) => addends_1_11_port, Y(10) => 
                           addends_1_10_port, Y(9) => addends_1_9_port, Y(8) =>
                           addends_1_8_port, Y(7) => addends_1_7_port, Y(6) => 
                           addends_1_6_port, Y(5) => addends_1_5_port, Y(4) => 
                           addends_1_4_port, Y(3) => addends_1_3_port, Y(2) => 
                           addends_1_2_port, Y(1) => addends_1_1_port, Y(0) => 
                           addends_1_0_port);
   MUX_I_2 : MUX5to1_NBIT32_6 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => A(15), B(18) => A(14), B(17)
                           => A(13), B(16) => A(12), B(15) => A(11), B(14) => 
                           A(10), B(13) => A(9), B(12) => A(8), B(11) => A(7), 
                           B(10) => A(6), B(9) => A(5), B(8) => A(4), B(7) => 
                           A(3), B(6) => A(2), B(5) => A(1), B(4) => n96, B(3) 
                           => X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n80, 
                           C(30) => n80, C(29) => n80, C(28) => n80, C(27) => 
                           n80, C(26) => n80, C(25) => n80, C(24) => n81, C(23)
                           => n81, C(22) => n81, C(21) => n81, C(20) => n81, 
                           C(19) => A_neg_9_24_port, C(18) => A_neg_9_23_port, 
                           C(17) => A_neg_9_22_port, C(16) => A_neg_9_21_port, 
                           C(15) => A_neg_9_20_port, C(14) => A_neg_9_19_port, 
                           C(13) => A_neg_9_18_port, C(12) => A_neg_9_17_port, 
                           C(11) => A_neg_9_16_port, C(10) => A_neg_9_15_port, 
                           C(9) => A_neg_9_14_port, C(8) => A_neg_9_13_port, 
                           C(7) => A_neg_9_12_port, C(6) => A_neg_9_11_port, 
                           C(5) => A_neg_9_10_port, C(4) => n94, C(3) => n69, 
                           C(2) => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => A(15), D(19) => A(14), D(18)
                           => A(13), D(17) => A(12), D(16) => A(11), D(15) => 
                           A(10), D(14) => A(9), D(13) => A(8), D(12) => A(7), 
                           D(11) => A(6), D(10) => A(5), D(9) => A(4), D(8) => 
                           A(3), D(7) => A(2), D(6) => A(1), D(5) => n94, D(4) 
                           => X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n85, E(30) => n84, E(29) => 
                           n85, E(28) => n84, E(27) => n84, E(26) => n85, E(25)
                           => n84, E(24) => n85, E(23) => n85, E(22) => n84, 
                           E(21) => n84, E(20) => A_neg_9_24_port, E(19) => 
                           A_neg_9_23_port, E(18) => A_neg_9_22_port, E(17) => 
                           A_neg_9_21_port, E(16) => A_neg_9_20_port, E(15) => 
                           A_neg_9_19_port, E(14) => A_neg_9_18_port, E(13) => 
                           A_neg_9_17_port, E(12) => A_neg_9_16_port, E(11) => 
                           A_neg_9_15_port, E(10) => A_neg_9_14_port, E(9) => 
                           A_neg_9_13_port, E(8) => A_neg_9_12_port, E(7) => 
                           A_neg_9_11_port, E(6) => A_neg_9_10_port, E(5) => 
                           n95, E(4) => n69, E(3) => n69, E(2) => n69, E(1) => 
                           n69, E(0) => n69, SEL(2) => selector_8_port, SEL(1) 
                           => selector_7_port, SEL(0) => selector_6_port, Y(31)
                           => mux_out_2_31_port, Y(30) => mux_out_2_30_port, 
                           Y(29) => mux_out_2_29_port, Y(28) => 
                           mux_out_2_28_port, Y(27) => mux_out_2_27_port, Y(26)
                           => mux_out_2_26_port, Y(25) => mux_out_2_25_port, 
                           Y(24) => mux_out_2_24_port, Y(23) => 
                           mux_out_2_23_port, Y(22) => mux_out_2_22_port, Y(21)
                           => mux_out_2_21_port, Y(20) => mux_out_2_20_port, 
                           Y(19) => mux_out_2_19_port, Y(18) => 
                           mux_out_2_18_port, Y(17) => mux_out_2_17_port, Y(16)
                           => mux_out_2_16_port, Y(15) => mux_out_2_15_port, 
                           Y(14) => mux_out_2_14_port, Y(13) => 
                           mux_out_2_13_port, Y(12) => mux_out_2_12_port, Y(11)
                           => mux_out_2_11_port, Y(10) => mux_out_2_10_port, 
                           Y(9) => mux_out_2_9_port, Y(8) => mux_out_2_8_port, 
                           Y(7) => mux_out_2_7_port, Y(6) => mux_out_2_6_port, 
                           Y(5) => mux_out_2_5_port, Y(4) => mux_out_2_4_port, 
                           Y(3) => mux_out_2_3_port, Y(2) => mux_out_2_2_port, 
                           Y(1) => mux_out_2_1_port, Y(0) => mux_out_2_0_port);
   MUX_I_3 : MUX5to1_NBIT32_5 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => A(15), B(20) => A(14), B(19)
                           => A(13), B(18) => A(12), B(17) => A(11), B(16) => 
                           A(10), B(15) => A(9), B(14) => A(8), B(13) => A(7), 
                           B(12) => A(6), B(11) => A(5), B(10) => A(4), B(9) =>
                           A(3), B(8) => A(2), B(7) => A(1), B(6) => n96, B(5) 
                           => X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n81, 
                           C(30) => n81, C(29) => n81, C(28) => n81, C(27) => 
                           n81, C(26) => n81, C(25) => n81, C(24) => n82, C(23)
                           => n82, C(22) => n82, C(21) => A_neg_9_24_port, 
                           C(20) => A_neg_9_23_port, C(19) => A_neg_9_22_port, 
                           C(18) => A_neg_9_21_port, C(17) => A_neg_9_20_port, 
                           C(16) => A_neg_9_19_port, C(15) => A_neg_9_18_port, 
                           C(14) => A_neg_9_17_port, C(13) => A_neg_9_16_port, 
                           C(12) => A_neg_9_15_port, C(11) => A_neg_9_14_port, 
                           C(10) => A_neg_9_13_port, C(9) => A_neg_9_12_port, 
                           C(8) => A_neg_9_11_port, C(7) => A_neg_9_10_port, 
                           C(6) => n94, C(5) => n69, C(4) => n69, C(3) => n69, 
                           C(2) => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => A(15), D(21) => A(14), D(20)
                           => A(13), D(19) => A(12), D(18) => A(11), D(17) => 
                           A(10), D(16) => A(9), D(15) => A(8), D(14) => A(7), 
                           D(13) => A(6), D(12) => A(5), D(11) => A(4), D(10) 
                           => A(3), D(9) => A(2), D(8) => A(1), D(7) => n94, 
                           D(6) => X_Logic0_port, D(5) => X_Logic0_port, D(4) 
                           => X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n84, E(30) => n84, E(29) => 
                           n84, E(28) => n85, E(27) => n86, E(26) => n84, E(25)
                           => n85, E(24) => n84, E(23) => n84, E(22) => 
                           A_neg_9_24_port, E(21) => A_neg_9_23_port, E(20) => 
                           A_neg_9_22_port, E(19) => A_neg_9_21_port, E(18) => 
                           A_neg_9_20_port, E(17) => A_neg_9_19_port, E(16) => 
                           A_neg_9_18_port, E(15) => A_neg_9_17_port, E(14) => 
                           A_neg_9_16_port, E(13) => A_neg_9_15_port, E(12) => 
                           A_neg_9_14_port, E(11) => A_neg_9_13_port, E(10) => 
                           A_neg_9_12_port, E(9) => A_neg_9_11_port, E(8) => 
                           A_neg_9_10_port, E(7) => n95, E(6) => n69, E(5) => 
                           n69, E(4) => n69, E(3) => n69, E(2) => n69, E(1) => 
                           n69, E(0) => n69, SEL(2) => selector_11_port, SEL(1)
                           => selector_10_port, SEL(0) => selector_9_port, 
                           Y(31) => mux_out_3_31_port, Y(30) => 
                           mux_out_3_30_port, Y(29) => mux_out_3_29_port, Y(28)
                           => mux_out_3_28_port, Y(27) => mux_out_3_27_port, 
                           Y(26) => mux_out_3_26_port, Y(25) => 
                           mux_out_3_25_port, Y(24) => mux_out_3_24_port, Y(23)
                           => mux_out_3_23_port, Y(22) => mux_out_3_22_port, 
                           Y(21) => mux_out_3_21_port, Y(20) => 
                           mux_out_3_20_port, Y(19) => mux_out_3_19_port, Y(18)
                           => mux_out_3_18_port, Y(17) => mux_out_3_17_port, 
                           Y(16) => mux_out_3_16_port, Y(15) => 
                           mux_out_3_15_port, Y(14) => mux_out_3_14_port, Y(13)
                           => mux_out_3_13_port, Y(12) => mux_out_3_12_port, 
                           Y(11) => mux_out_3_11_port, Y(10) => 
                           mux_out_3_10_port, Y(9) => mux_out_3_9_port, Y(8) =>
                           mux_out_3_8_port, Y(7) => mux_out_3_7_port, Y(6) => 
                           mux_out_3_6_port, Y(5) => mux_out_3_5_port, Y(4) => 
                           mux_out_3_4_port, Y(3) => mux_out_3_3_port, Y(2) => 
                           mux_out_3_2_port, Y(1) => mux_out_3_1_port, Y(0) => 
                           mux_out_3_0_port);
   MUX_I_4 : MUX5to1_NBIT32_4 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => A(15), B(22) => A(14), B(21)
                           => A(13), B(20) => A(12), B(19) => A(11), B(18) => 
                           A(10), B(17) => A(9), B(16) => A(8), B(15) => A(7), 
                           B(14) => A(6), B(13) => A(5), B(12) => A(4), B(11) 
                           => A(3), B(10) => A(2), B(9) => A(1), B(8) => n96, 
                           B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) 
                           => X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n82, 
                           C(30) => n83, C(29) => n83, C(28) => n82, C(27) => 
                           n83, C(26) => n83, C(25) => n83, C(24) => n83, C(23)
                           => A_neg_9_24_port, C(22) => A_neg_9_23_port, C(21) 
                           => A_neg_9_22_port, C(20) => A_neg_9_21_port, C(19) 
                           => A_neg_9_20_port, C(18) => A_neg_9_19_port, C(17) 
                           => A_neg_9_18_port, C(16) => A_neg_9_17_port, C(15) 
                           => A_neg_9_16_port, C(14) => A_neg_9_15_port, C(13) 
                           => A_neg_9_14_port, C(12) => A_neg_9_13_port, C(11) 
                           => A_neg_9_12_port, C(10) => A_neg_9_11_port, C(9) 
                           => A_neg_9_10_port, C(8) => n94, C(7) => n69, C(6) 
                           => n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) 
                           => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => A(15), D(23) => A(14), D(22)
                           => A(13), D(21) => A(12), D(20) => A(11), D(19) => 
                           A(10), D(18) => A(9), D(17) => A(8), D(16) => A(7), 
                           D(15) => A(6), D(14) => A(5), D(13) => A(4), D(12) 
                           => A(3), D(11) => A(2), D(10) => A(1), D(9) => n94, 
                           D(8) => X_Logic0_port, D(7) => X_Logic0_port, D(6) 
                           => X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n87, E(30) => n86, E(29) => 
                           n86, E(28) => n87, E(27) => n86, E(26) => n86, E(25)
                           => n87, E(24) => A_neg_9_24_port, E(23) => 
                           A_neg_9_23_port, E(22) => A_neg_9_22_port, E(21) => 
                           A_neg_9_21_port, E(20) => A_neg_9_20_port, E(19) => 
                           A_neg_9_19_port, E(18) => A_neg_9_18_port, E(17) => 
                           A_neg_9_17_port, E(16) => A_neg_9_16_port, E(15) => 
                           A_neg_9_15_port, E(14) => A_neg_9_14_port, E(13) => 
                           A_neg_9_13_port, E(12) => A_neg_9_12_port, E(11) => 
                           A_neg_9_11_port, E(10) => A_neg_9_10_port, E(9) => 
                           n95, E(8) => n69, E(7) => n69, E(6) => n69, E(5) => 
                           n69, E(4) => n69, E(3) => n69, E(2) => n69, E(1) => 
                           n69, E(0) => n69, SEL(2) => selector_14_port, SEL(1)
                           => selector_13_port, SEL(0) => selector_12_port, 
                           Y(31) => mux_out_4_31_port, Y(30) => 
                           mux_out_4_30_port, Y(29) => mux_out_4_29_port, Y(28)
                           => mux_out_4_28_port, Y(27) => mux_out_4_27_port, 
                           Y(26) => mux_out_4_26_port, Y(25) => 
                           mux_out_4_25_port, Y(24) => mux_out_4_24_port, Y(23)
                           => mux_out_4_23_port, Y(22) => mux_out_4_22_port, 
                           Y(21) => mux_out_4_21_port, Y(20) => 
                           mux_out_4_20_port, Y(19) => mux_out_4_19_port, Y(18)
                           => mux_out_4_18_port, Y(17) => mux_out_4_17_port, 
                           Y(16) => mux_out_4_16_port, Y(15) => 
                           mux_out_4_15_port, Y(14) => mux_out_4_14_port, Y(13)
                           => mux_out_4_13_port, Y(12) => mux_out_4_12_port, 
                           Y(11) => mux_out_4_11_port, Y(10) => 
                           mux_out_4_10_port, Y(9) => mux_out_4_9_port, Y(8) =>
                           mux_out_4_8_port, Y(7) => mux_out_4_7_port, Y(6) => 
                           mux_out_4_6_port, Y(5) => mux_out_4_5_port, Y(4) => 
                           mux_out_4_4_port, Y(3) => mux_out_4_3_port, Y(2) => 
                           mux_out_4_2_port, Y(1) => mux_out_4_1_port, Y(0) => 
                           mux_out_4_0_port);
   MUX_I_5 : MUX5to1_NBIT32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => A(15), B(24) => A(14), B(23)
                           => A(13), B(22) => A(12), B(21) => A(11), B(20) => 
                           A(10), B(19) => A(9), B(18) => A(8), B(17) => A(7), 
                           B(16) => A(6), B(15) => A(5), B(14) => A(4), B(13) 
                           => A(3), B(12) => A(2), B(11) => A(1), B(10) => n96,
                           B(9) => X_Logic0_port, B(8) => X_Logic0_port, B(7) 
                           => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n82, 
                           C(30) => n82, C(29) => n82, C(28) => n83, C(27) => 
                           n83, C(26) => n82, C(25) => A_neg_9_24_port, C(24) 
                           => A_neg_9_23_port, C(23) => A_neg_9_22_port, C(22) 
                           => A_neg_9_21_port, C(21) => A_neg_9_20_port, C(20) 
                           => A_neg_9_19_port, C(19) => A_neg_9_18_port, C(18) 
                           => A_neg_9_17_port, C(17) => A_neg_9_16_port, C(16) 
                           => A_neg_9_15_port, C(15) => A_neg_9_14_port, C(14) 
                           => A_neg_9_13_port, C(13) => A_neg_9_12_port, C(12) 
                           => A_neg_9_11_port, C(11) => A_neg_9_10_port, C(10) 
                           => n95, C(9) => n69, C(8) => n69, C(7) => n69, C(6) 
                           => n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) 
                           => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => A(15), D(25) => A(14), D(24)
                           => A(13), D(23) => A(12), D(22) => A(11), D(21) => 
                           A(10), D(20) => A(9), D(19) => A(8), D(18) => A(7), 
                           D(17) => A(6), D(16) => A(5), D(15) => A(4), D(14) 
                           => A(3), D(13) => A(2), D(12) => A(1), D(11) => n94,
                           D(10) => X_Logic0_port, D(9) => X_Logic0_port, D(8) 
                           => X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n88, E(30) => n88, E(29) => 
                           n88, E(28) => n88, E(27) => n88, E(26) => 
                           A_neg_9_24_port, E(25) => A_neg_9_23_port, E(24) => 
                           A_neg_9_22_port, E(23) => A_neg_9_21_port, E(22) => 
                           A_neg_9_20_port, E(21) => A_neg_9_19_port, E(20) => 
                           A_neg_9_18_port, E(19) => A_neg_9_17_port, E(18) => 
                           A_neg_9_16_port, E(17) => A_neg_9_15_port, E(16) => 
                           A_neg_9_14_port, E(15) => A_neg_9_13_port, E(14) => 
                           A_neg_9_12_port, E(13) => A_neg_9_11_port, E(12) => 
                           A_neg_9_10_port, E(11) => n95, E(10) => n69, E(9) =>
                           n69, E(8) => n69, E(7) => n69, E(6) => n69, E(5) => 
                           n69, E(4) => n69, E(3) => n69, E(2) => n69, E(1) => 
                           n69, E(0) => n69, SEL(2) => selector_17_port, SEL(1)
                           => selector_16_port, SEL(0) => selector_15_port, 
                           Y(31) => mux_out_5_31_port, Y(30) => 
                           mux_out_5_30_port, Y(29) => mux_out_5_29_port, Y(28)
                           => mux_out_5_28_port, Y(27) => mux_out_5_27_port, 
                           Y(26) => mux_out_5_26_port, Y(25) => 
                           mux_out_5_25_port, Y(24) => mux_out_5_24_port, Y(23)
                           => mux_out_5_23_port, Y(22) => mux_out_5_22_port, 
                           Y(21) => mux_out_5_21_port, Y(20) => 
                           mux_out_5_20_port, Y(19) => mux_out_5_19_port, Y(18)
                           => mux_out_5_18_port, Y(17) => mux_out_5_17_port, 
                           Y(16) => mux_out_5_16_port, Y(15) => 
                           mux_out_5_15_port, Y(14) => mux_out_5_14_port, Y(13)
                           => mux_out_5_13_port, Y(12) => mux_out_5_12_port, 
                           Y(11) => mux_out_5_11_port, Y(10) => 
                           mux_out_5_10_port, Y(9) => mux_out_5_9_port, Y(8) =>
                           mux_out_5_8_port, Y(7) => mux_out_5_7_port, Y(6) => 
                           mux_out_5_6_port, Y(5) => mux_out_5_5_port, Y(4) => 
                           mux_out_5_4_port, Y(3) => mux_out_5_3_port, Y(2) => 
                           mux_out_5_2_port, Y(1) => mux_out_5_1_port, Y(0) => 
                           mux_out_5_0_port);
   MUX_I_6 : MUX5to1_NBIT32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => A(15), B(26) => A(14), B(25)
                           => A(13), B(24) => A(12), B(23) => A(11), B(22) => 
                           A(10), B(21) => A(9), B(20) => A(8), B(19) => A(7), 
                           B(18) => A(6), B(17) => A(5), B(16) => A(4), B(15) 
                           => A(3), B(14) => A(2), B(13) => A(1), B(12) => n96,
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n82, 
                           C(30) => n83, C(29) => n82, C(28) => n83, C(27) => 
                           A_neg_9_24_port, C(26) => A_neg_9_23_port, C(25) => 
                           A_neg_9_22_port, C(24) => A_neg_9_21_port, C(23) => 
                           A_neg_9_20_port, C(22) => A_neg_9_19_port, C(21) => 
                           A_neg_9_18_port, C(20) => A_neg_9_17_port, C(19) => 
                           A_neg_9_16_port, C(18) => A_neg_9_15_port, C(17) => 
                           A_neg_9_14_port, C(16) => A_neg_9_13_port, C(15) => 
                           A_neg_9_12_port, C(14) => A_neg_9_11_port, C(13) => 
                           A_neg_9_10_port, C(12) => n95, C(11) => n69, C(10) 
                           => n69, C(9) => n69, C(8) => n69, C(7) => n69, C(6) 
                           => n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) 
                           => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => A(15), D(27) => A(14), D(26)
                           => A(13), D(25) => A(12), D(24) => A(11), D(23) => 
                           A(10), D(22) => A(9), D(21) => A(8), D(20) => A(7), 
                           D(19) => A(6), D(18) => A(5), D(17) => A(4), D(16) 
                           => A(3), D(15) => A(2), D(14) => A(1), D(13) => n94,
                           D(12) => X_Logic0_port, D(11) => X_Logic0_port, 
                           D(10) => X_Logic0_port, D(9) => X_Logic0_port, D(8) 
                           => X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n89, E(30) => n89, E(29) => 
                           n89, E(28) => A_neg_9_24_port, E(27) => 
                           A_neg_9_23_port, E(26) => A_neg_9_22_port, E(25) => 
                           A_neg_9_21_port, E(24) => A_neg_9_20_port, E(23) => 
                           A_neg_9_19_port, E(22) => A_neg_9_18_port, E(21) => 
                           A_neg_9_17_port, E(20) => A_neg_9_16_port, E(19) => 
                           A_neg_9_15_port, E(18) => A_neg_9_14_port, E(17) => 
                           A_neg_9_13_port, E(16) => A_neg_9_12_port, E(15) => 
                           A_neg_9_11_port, E(14) => A_neg_9_10_port, E(13) => 
                           n96, E(12) => n69, E(11) => n69, E(10) => n69, E(9) 
                           => n69, E(8) => n69, E(7) => n69, E(6) => n69, E(5) 
                           => n69, E(4) => n69, E(3) => n69, E(2) => n69, E(1) 
                           => n69, E(0) => n69, SEL(2) => selector_20_port, 
                           SEL(1) => selector_19_port, SEL(0) => 
                           selector_18_port, Y(31) => mux_out_6_31_port, Y(30) 
                           => mux_out_6_30_port, Y(29) => mux_out_6_29_port, 
                           Y(28) => mux_out_6_28_port, Y(27) => 
                           mux_out_6_27_port, Y(26) => mux_out_6_26_port, Y(25)
                           => mux_out_6_25_port, Y(24) => mux_out_6_24_port, 
                           Y(23) => mux_out_6_23_port, Y(22) => 
                           mux_out_6_22_port, Y(21) => mux_out_6_21_port, Y(20)
                           => mux_out_6_20_port, Y(19) => mux_out_6_19_port, 
                           Y(18) => mux_out_6_18_port, Y(17) => 
                           mux_out_6_17_port, Y(16) => mux_out_6_16_port, Y(15)
                           => mux_out_6_15_port, Y(14) => mux_out_6_14_port, 
                           Y(13) => mux_out_6_13_port, Y(12) => 
                           mux_out_6_12_port, Y(11) => mux_out_6_11_port, Y(10)
                           => mux_out_6_10_port, Y(9) => mux_out_6_9_port, Y(8)
                           => mux_out_6_8_port, Y(7) => mux_out_6_7_port, Y(6) 
                           => mux_out_6_6_port, Y(5) => mux_out_6_5_port, Y(4) 
                           => mux_out_6_4_port, Y(3) => mux_out_6_3_port, Y(2) 
                           => mux_out_6_2_port, Y(1) => mux_out_6_1_port, Y(0) 
                           => mux_out_6_0_port);
   MUX_I_7 : MUX5to1_NBIT32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => A(15), B(28) => A(14), B(27)
                           => A(13), B(26) => A(12), B(25) => A(11), B(24) => 
                           A(10), B(23) => A(9), B(22) => A(8), B(21) => A(7), 
                           B(20) => A(6), B(19) => A(5), B(18) => A(4), B(17) 
                           => A(3), B(16) => A(2), B(15) => A(1), B(14) => n96,
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n83, 
                           C(30) => n83, C(29) => A_neg_9_24_port, C(28) => 
                           A_neg_9_23_port, C(27) => A_neg_9_22_port, C(26) => 
                           A_neg_9_21_port, C(25) => A_neg_9_20_port, C(24) => 
                           A_neg_9_19_port, C(23) => A_neg_9_18_port, C(22) => 
                           A_neg_9_17_port, C(21) => A_neg_9_16_port, C(20) => 
                           A_neg_9_15_port, C(19) => A_neg_9_14_port, C(18) => 
                           A_neg_9_13_port, C(17) => A_neg_9_12_port, C(16) => 
                           A_neg_9_11_port, C(15) => A_neg_9_10_port, C(14) => 
                           n95, C(13) => n69, C(12) => n69, C(11) => n69, C(10)
                           => n69, C(9) => n69, C(8) => n69, C(7) => n69, C(6) 
                           => n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) 
                           => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => A(15), D(29) => A(14), D(28)
                           => A(13), D(27) => A(12), D(26) => A(11), D(25) => 
                           A(10), D(24) => A(9), D(23) => A(8), D(22) => A(7), 
                           D(21) => A(6), D(20) => A(5), D(19) => A(4), D(18) 
                           => A(3), D(17) => A(2), D(16) => A(1), D(15) => n94,
                           D(14) => X_Logic0_port, D(13) => X_Logic0_port, 
                           D(12) => X_Logic0_port, D(11) => X_Logic0_port, 
                           D(10) => X_Logic0_port, D(9) => X_Logic0_port, D(8) 
                           => X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n89, E(30) => 
                           A_neg_9_24_port, E(29) => A_neg_9_23_port, E(28) => 
                           A_neg_9_22_port, E(27) => A_neg_9_21_port, E(26) => 
                           A_neg_9_20_port, E(25) => A_neg_9_19_port, E(24) => 
                           A_neg_9_18_port, E(23) => A_neg_9_17_port, E(22) => 
                           A_neg_9_16_port, E(21) => A_neg_9_15_port, E(20) => 
                           A_neg_9_14_port, E(19) => A_neg_9_13_port, E(18) => 
                           A_neg_9_12_port, E(17) => A_neg_9_11_port, E(16) => 
                           A_neg_9_10_port, E(15) => n95, E(14) => n69, E(13) 
                           => n69, E(12) => n69, E(11) => n69, E(10) => n69, 
                           E(9) => n69, E(8) => n69, E(7) => n69, E(6) => n69, 
                           E(5) => n69, E(4) => n69, E(3) => n69, E(2) => n69, 
                           E(1) => n69, E(0) => n69, SEL(2) => selector_23_port
                           , SEL(1) => selector_22_port, SEL(0) => 
                           selector_21_port, Y(31) => mux_out_7_31_port, Y(30) 
                           => mux_out_7_30_port, Y(29) => mux_out_7_29_port, 
                           Y(28) => mux_out_7_28_port, Y(27) => 
                           mux_out_7_27_port, Y(26) => mux_out_7_26_port, Y(25)
                           => mux_out_7_25_port, Y(24) => mux_out_7_24_port, 
                           Y(23) => mux_out_7_23_port, Y(22) => 
                           mux_out_7_22_port, Y(21) => mux_out_7_21_port, Y(20)
                           => mux_out_7_20_port, Y(19) => mux_out_7_19_port, 
                           Y(18) => mux_out_7_18_port, Y(17) => 
                           mux_out_7_17_port, Y(16) => mux_out_7_16_port, Y(15)
                           => mux_out_7_15_port, Y(14) => mux_out_7_14_port, 
                           Y(13) => mux_out_7_13_port, Y(12) => 
                           mux_out_7_12_port, Y(11) => mux_out_7_11_port, Y(10)
                           => mux_out_7_10_port, Y(9) => mux_out_7_9_port, Y(8)
                           => mux_out_7_8_port, Y(7) => mux_out_7_7_port, Y(6) 
                           => mux_out_7_6_port, Y(5) => mux_out_7_5_port, Y(4) 
                           => mux_out_7_4_port, Y(3) => mux_out_7_3_port, Y(2) 
                           => mux_out_7_2_port, Y(1) => mux_out_7_1_port, Y(0) 
                           => mux_out_7_0_port);
   ADD0 : ADDER_NBIT32_NBIT_PER_BLOCK4_7 port map( A(31) => addends_0_31_port, 
                           A(30) => addends_0_30_port, A(29) => 
                           addends_0_29_port, A(28) => addends_0_28_port, A(27)
                           => addends_0_27_port, A(26) => addends_0_26_port, 
                           A(25) => addends_0_25_port, A(24) => 
                           addends_0_24_port, A(23) => addends_0_23_port, A(22)
                           => addends_0_22_port, A(21) => addends_0_21_port, 
                           A(20) => addends_0_20_port, A(19) => 
                           addends_0_19_port, A(18) => addends_0_18_port, A(17)
                           => addends_0_17_port, A(16) => addends_0_16_port, 
                           A(15) => addends_0_15_port, A(14) => 
                           addends_0_14_port, A(13) => addends_0_13_port, A(12)
                           => addends_0_12_port, A(11) => addends_0_11_port, 
                           A(10) => addends_0_10_port, A(9) => addends_0_9_port
                           , A(8) => addends_0_8_port, A(7) => addends_0_7_port
                           , A(6) => addends_0_6_port, A(5) => addends_0_5_port
                           , A(4) => addends_0_4_port, A(3) => addends_0_3_port
                           , A(2) => addends_0_2_port, A(1) => addends_0_1_port
                           , A(0) => addends_0_0_port, B(31) => 
                           addends_1_31_port, B(30) => addends_1_30_port, B(29)
                           => addends_1_29_port, B(28) => addends_1_28_port, 
                           B(27) => addends_1_27_port, B(26) => 
                           addends_1_26_port, B(25) => addends_1_25_port, B(24)
                           => addends_1_24_port, B(23) => addends_1_23_port, 
                           B(22) => addends_1_22_port, B(21) => 
                           addends_1_21_port, B(20) => addends_1_20_port, B(19)
                           => addends_1_19_port, B(18) => addends_1_18_port, 
                           B(17) => addends_1_17_port, B(16) => 
                           addends_1_16_port, B(15) => addends_1_15_port, B(14)
                           => addends_1_14_port, B(13) => addends_1_13_port, 
                           B(12) => addends_1_12_port, B(11) => 
                           addends_1_11_port, B(10) => addends_1_10_port, B(9) 
                           => addends_1_9_port, B(8) => addends_1_8_port, B(7) 
                           => addends_1_7_port, B(6) => addends_1_6_port, B(5) 
                           => addends_1_5_port, B(4) => addends_1_4_port, B(3) 
                           => addends_1_3_port, B(2) => addends_1_2_port, B(1) 
                           => addends_1_1_port, B(0) => addends_1_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_0_31_port, S(30) => reg_in_0_30_port
                           , S(29) => reg_in_0_29_port, S(28) => 
                           reg_in_0_28_port, S(27) => reg_in_0_27_port, S(26) 
                           => reg_in_0_26_port, S(25) => reg_in_0_25_port, 
                           S(24) => reg_in_0_24_port, S(23) => reg_in_0_23_port
                           , S(22) => reg_in_0_22_port, S(21) => 
                           reg_in_0_21_port, S(20) => reg_in_0_20_port, S(19) 
                           => reg_in_0_19_port, S(18) => reg_in_0_18_port, 
                           S(17) => reg_in_0_17_port, S(16) => reg_in_0_16_port
                           , S(15) => reg_in_0_15_port, S(14) => 
                           reg_in_0_14_port, S(13) => reg_in_0_13_port, S(12) 
                           => reg_in_0_12_port, S(11) => reg_in_0_11_port, 
                           S(10) => reg_in_0_10_port, S(9) => reg_in_0_9_port, 
                           S(8) => reg_in_0_8_port, S(7) => reg_in_0_7_port, 
                           S(6) => reg_in_0_6_port, S(5) => reg_in_0_5_port, 
                           S(4) => reg_in_0_4_port, S(3) => reg_in_0_3_port, 
                           S(2) => reg_in_0_2_port, S(1) => reg_in_0_1_port, 
                           S(0) => reg_in_0_0_port, Cout => n_1521);
   REG0 : REG_NBIT32_3 port map( clk => CLOCK, reset => X_Logic0_port, enable 
                           => X_Logic1_port, data_in(31) => reg_in_0_31_port, 
                           data_in(30) => reg_in_0_30_port, data_in(29) => 
                           reg_in_0_29_port, data_in(28) => reg_in_0_28_port, 
                           data_in(27) => reg_in_0_27_port, data_in(26) => 
                           reg_in_0_26_port, data_in(25) => reg_in_0_25_port, 
                           data_in(24) => reg_in_0_24_port, data_in(23) => 
                           reg_in_0_23_port, data_in(22) => reg_in_0_22_port, 
                           data_in(21) => reg_in_0_21_port, data_in(20) => 
                           reg_in_0_20_port, data_in(19) => reg_in_0_19_port, 
                           data_in(18) => reg_in_0_18_port, data_in(17) => 
                           reg_in_0_17_port, data_in(16) => reg_in_0_16_port, 
                           data_in(15) => reg_in_0_15_port, data_in(14) => 
                           reg_in_0_14_port, data_in(13) => reg_in_0_13_port, 
                           data_in(12) => reg_in_0_12_port, data_in(11) => 
                           reg_in_0_11_port, data_in(10) => reg_in_0_10_port, 
                           data_in(9) => reg_in_0_9_port, data_in(8) => 
                           reg_in_0_8_port, data_in(7) => reg_in_0_7_port, 
                           data_in(6) => reg_in_0_6_port, data_in(5) => 
                           reg_in_0_5_port, data_in(4) => reg_in_0_4_port, 
                           data_in(3) => reg_in_0_3_port, data_in(2) => 
                           reg_in_0_2_port, data_in(1) => reg_in_0_1_port, 
                           data_in(0) => reg_in_0_0_port, data_out(31) => 
                           reg_out_0_31_port, data_out(30) => reg_out_0_30_port
                           , data_out(29) => reg_out_0_29_port, data_out(28) =>
                           reg_out_0_28_port, data_out(27) => reg_out_0_27_port
                           , data_out(26) => reg_out_0_26_port, data_out(25) =>
                           reg_out_0_25_port, data_out(24) => reg_out_0_24_port
                           , data_out(23) => reg_out_0_23_port, data_out(22) =>
                           reg_out_0_22_port, data_out(21) => reg_out_0_21_port
                           , data_out(20) => reg_out_0_20_port, data_out(19) =>
                           reg_out_0_19_port, data_out(18) => reg_out_0_18_port
                           , data_out(17) => reg_out_0_17_port, data_out(16) =>
                           reg_out_0_16_port, data_out(15) => reg_out_0_15_port
                           , data_out(14) => reg_out_0_14_port, data_out(13) =>
                           reg_out_0_13_port, data_out(12) => reg_out_0_12_port
                           , data_out(11) => reg_out_0_11_port, data_out(10) =>
                           reg_out_0_10_port, data_out(9) => reg_out_0_9_port, 
                           data_out(8) => reg_out_0_8_port, data_out(7) => 
                           reg_out_0_7_port, data_out(6) => reg_out_0_6_port, 
                           data_out(5) => reg_out_0_5_port, data_out(4) => 
                           reg_out_0_4_port, data_out(3) => reg_out_0_3_port, 
                           data_out(2) => reg_out_0_2_port, data_out(1) => 
                           reg_out_0_1_port, data_out(0) => reg_out_0_0_port);
   ADD_0i_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_6 port map( A(31) => 
                           reg_out_0_31_port, A(30) => reg_out_0_30_port, A(29)
                           => reg_out_0_29_port, A(28) => reg_out_0_28_port, 
                           A(27) => reg_out_0_27_port, A(26) => 
                           reg_out_0_26_port, A(25) => reg_out_0_25_port, A(24)
                           => reg_out_0_24_port, A(23) => reg_out_0_23_port, 
                           A(22) => reg_out_0_22_port, A(21) => 
                           reg_out_0_21_port, A(20) => reg_out_0_20_port, A(19)
                           => reg_out_0_19_port, A(18) => reg_out_0_18_port, 
                           A(17) => reg_out_0_17_port, A(16) => 
                           reg_out_0_16_port, A(15) => reg_out_0_15_port, A(14)
                           => reg_out_0_14_port, A(13) => reg_out_0_13_port, 
                           A(12) => reg_out_0_12_port, A(11) => 
                           reg_out_0_11_port, A(10) => reg_out_0_10_port, A(9) 
                           => reg_out_0_9_port, A(8) => reg_out_0_8_port, A(7) 
                           => reg_out_0_7_port, A(6) => reg_out_0_6_port, A(5) 
                           => reg_out_0_5_port, A(4) => reg_out_0_4_port, A(3) 
                           => reg_out_0_3_port, A(2) => reg_out_0_2_port, A(1) 
                           => reg_out_0_1_port, A(0) => reg_out_0_0_port, B(31)
                           => addends_2_31_port, B(30) => addends_2_30_port, 
                           B(29) => addends_2_29_port, B(28) => 
                           addends_2_28_port, B(27) => addends_2_27_port, B(26)
                           => addends_2_26_port, B(25) => addends_2_25_port, 
                           B(24) => addends_2_24_port, B(23) => 
                           addends_2_23_port, B(22) => addends_2_22_port, B(21)
                           => addends_2_21_port, B(20) => addends_2_20_port, 
                           B(19) => addends_2_19_port, B(18) => 
                           addends_2_18_port, B(17) => addends_2_17_port, B(16)
                           => addends_2_16_port, B(15) => addends_2_15_port, 
                           B(14) => addends_2_14_port, B(13) => 
                           addends_2_13_port, B(12) => addends_2_12_port, B(11)
                           => addends_2_11_port, B(10) => addends_2_10_port, 
                           B(9) => addends_2_9_port, B(8) => addends_2_8_port, 
                           B(7) => addends_2_7_port, B(6) => addends_2_6_port, 
                           B(5) => addends_2_5_port, B(4) => addends_2_4_port, 
                           B(3) => addends_2_3_port, B(2) => addends_2_2_port, 
                           B(1) => addends_2_1_port, B(0) => addends_2_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_0_31_port, S(30) => 
                           add_out_0_30_port, S(29) => add_out_0_29_port, S(28)
                           => add_out_0_28_port, S(27) => add_out_0_27_port, 
                           S(26) => add_out_0_26_port, S(25) => 
                           add_out_0_25_port, S(24) => add_out_0_24_port, S(23)
                           => add_out_0_23_port, S(22) => add_out_0_22_port, 
                           S(21) => add_out_0_21_port, S(20) => 
                           add_out_0_20_port, S(19) => add_out_0_19_port, S(18)
                           => add_out_0_18_port, S(17) => add_out_0_17_port, 
                           S(16) => add_out_0_16_port, S(15) => 
                           add_out_0_15_port, S(14) => add_out_0_14_port, S(13)
                           => add_out_0_13_port, S(12) => add_out_0_12_port, 
                           S(11) => add_out_0_11_port, S(10) => 
                           add_out_0_10_port, S(9) => add_out_0_9_port, S(8) =>
                           add_out_0_8_port, S(7) => add_out_0_7_port, S(6) => 
                           add_out_0_6_port, S(5) => add_out_0_5_port, S(4) => 
                           add_out_0_4_port, S(3) => add_out_0_3_port, S(2) => 
                           add_out_0_2_port, S(1) => add_out_0_1_port, S(0) => 
                           add_out_0_0_port, Cout => n_1522);
   ADD_1i_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_5 port map( A(31) => 
                           add_out_0_31_port, A(30) => add_out_0_30_port, A(29)
                           => add_out_0_29_port, A(28) => add_out_0_28_port, 
                           A(27) => add_out_0_27_port, A(26) => 
                           add_out_0_26_port, A(25) => add_out_0_25_port, A(24)
                           => add_out_0_24_port, A(23) => add_out_0_23_port, 
                           A(22) => add_out_0_22_port, A(21) => 
                           add_out_0_21_port, A(20) => add_out_0_20_port, A(19)
                           => add_out_0_19_port, A(18) => add_out_0_18_port, 
                           A(17) => add_out_0_17_port, A(16) => 
                           add_out_0_16_port, A(15) => add_out_0_15_port, A(14)
                           => add_out_0_14_port, A(13) => add_out_0_13_port, 
                           A(12) => add_out_0_12_port, A(11) => 
                           add_out_0_11_port, A(10) => add_out_0_10_port, A(9) 
                           => add_out_0_9_port, A(8) => add_out_0_8_port, A(7) 
                           => add_out_0_7_port, A(6) => add_out_0_6_port, A(5) 
                           => add_out_0_5_port, A(4) => add_out_0_4_port, A(3) 
                           => add_out_0_3_port, A(2) => add_out_0_2_port, A(1) 
                           => add_out_0_1_port, A(0) => add_out_0_0_port, B(31)
                           => addends_3_31_port, B(30) => addends_3_30_port, 
                           B(29) => addends_3_29_port, B(28) => 
                           addends_3_28_port, B(27) => addends_3_27_port, B(26)
                           => addends_3_26_port, B(25) => addends_3_25_port, 
                           B(24) => addends_3_24_port, B(23) => 
                           addends_3_23_port, B(22) => addends_3_22_port, B(21)
                           => addends_3_21_port, B(20) => addends_3_20_port, 
                           B(19) => addends_3_19_port, B(18) => 
                           addends_3_18_port, B(17) => addends_3_17_port, B(16)
                           => addends_3_16_port, B(15) => addends_3_15_port, 
                           B(14) => addends_3_14_port, B(13) => 
                           addends_3_13_port, B(12) => addends_3_12_port, B(11)
                           => addends_3_11_port, B(10) => addends_3_10_port, 
                           B(9) => addends_3_9_port, B(8) => addends_3_8_port, 
                           B(7) => addends_3_7_port, B(6) => addends_3_6_port, 
                           B(5) => addends_3_5_port, B(4) => addends_3_4_port, 
                           B(3) => addends_3_3_port, B(2) => addends_3_2_port, 
                           B(1) => addends_3_1_port, B(0) => addends_3_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_1_31_port, S(30) => reg_in_1_30_port
                           , S(29) => reg_in_1_29_port, S(28) => 
                           reg_in_1_28_port, S(27) => reg_in_1_27_port, S(26) 
                           => reg_in_1_26_port, S(25) => reg_in_1_25_port, 
                           S(24) => reg_in_1_24_port, S(23) => reg_in_1_23_port
                           , S(22) => reg_in_1_22_port, S(21) => 
                           reg_in_1_21_port, S(20) => reg_in_1_20_port, S(19) 
                           => reg_in_1_19_port, S(18) => reg_in_1_18_port, 
                           S(17) => reg_in_1_17_port, S(16) => reg_in_1_16_port
                           , S(15) => reg_in_1_15_port, S(14) => 
                           reg_in_1_14_port, S(13) => reg_in_1_13_port, S(12) 
                           => reg_in_1_12_port, S(11) => reg_in_1_11_port, 
                           S(10) => reg_in_1_10_port, S(9) => reg_in_1_9_port, 
                           S(8) => reg_in_1_8_port, S(7) => reg_in_1_7_port, 
                           S(6) => reg_in_1_6_port, S(5) => reg_in_1_5_port, 
                           S(4) => reg_in_1_4_port, S(3) => reg_in_1_3_port, 
                           S(2) => reg_in_1_2_port, S(1) => reg_in_1_1_port, 
                           S(0) => reg_in_1_0_port, Cout => n_1523);
   REG_i_1 : REG_NBIT32_2 port map( clk => CLOCK, reset => X_Logic0_port, 
                           enable => X_Logic1_port, data_in(31) => 
                           reg_in_1_31_port, data_in(30) => reg_in_1_30_port, 
                           data_in(29) => reg_in_1_29_port, data_in(28) => 
                           reg_in_1_28_port, data_in(27) => reg_in_1_27_port, 
                           data_in(26) => reg_in_1_26_port, data_in(25) => 
                           reg_in_1_25_port, data_in(24) => reg_in_1_24_port, 
                           data_in(23) => reg_in_1_23_port, data_in(22) => 
                           reg_in_1_22_port, data_in(21) => reg_in_1_21_port, 
                           data_in(20) => reg_in_1_20_port, data_in(19) => 
                           reg_in_1_19_port, data_in(18) => reg_in_1_18_port, 
                           data_in(17) => reg_in_1_17_port, data_in(16) => 
                           reg_in_1_16_port, data_in(15) => reg_in_1_15_port, 
                           data_in(14) => reg_in_1_14_port, data_in(13) => 
                           reg_in_1_13_port, data_in(12) => reg_in_1_12_port, 
                           data_in(11) => reg_in_1_11_port, data_in(10) => 
                           reg_in_1_10_port, data_in(9) => reg_in_1_9_port, 
                           data_in(8) => reg_in_1_8_port, data_in(7) => 
                           reg_in_1_7_port, data_in(6) => reg_in_1_6_port, 
                           data_in(5) => reg_in_1_5_port, data_in(4) => 
                           reg_in_1_4_port, data_in(3) => reg_in_1_3_port, 
                           data_in(2) => reg_in_1_2_port, data_in(1) => 
                           reg_in_1_1_port, data_in(0) => reg_in_1_0_port, 
                           data_out(31) => reg_out_1_31_port, data_out(30) => 
                           reg_out_1_30_port, data_out(29) => reg_out_1_29_port
                           , data_out(28) => reg_out_1_28_port, data_out(27) =>
                           reg_out_1_27_port, data_out(26) => reg_out_1_26_port
                           , data_out(25) => reg_out_1_25_port, data_out(24) =>
                           reg_out_1_24_port, data_out(23) => reg_out_1_23_port
                           , data_out(22) => reg_out_1_22_port, data_out(21) =>
                           reg_out_1_21_port, data_out(20) => reg_out_1_20_port
                           , data_out(19) => reg_out_1_19_port, data_out(18) =>
                           reg_out_1_18_port, data_out(17) => reg_out_1_17_port
                           , data_out(16) => reg_out_1_16_port, data_out(15) =>
                           reg_out_1_15_port, data_out(14) => reg_out_1_14_port
                           , data_out(13) => reg_out_1_13_port, data_out(12) =>
                           reg_out_1_12_port, data_out(11) => reg_out_1_11_port
                           , data_out(10) => reg_out_1_10_port, data_out(9) => 
                           reg_out_1_9_port, data_out(8) => reg_out_1_8_port, 
                           data_out(7) => reg_out_1_7_port, data_out(6) => 
                           reg_out_1_6_port, data_out(5) => reg_out_1_5_port, 
                           data_out(4) => reg_out_1_4_port, data_out(3) => 
                           reg_out_1_3_port, data_out(2) => reg_out_1_2_port, 
                           data_out(1) => reg_out_1_1_port, data_out(0) => 
                           reg_out_1_0_port);
   ADD_0i_2 : ADDER_NBIT32_NBIT_PER_BLOCK4_4 port map( A(31) => 
                           reg_out_1_31_port, A(30) => reg_out_1_30_port, A(29)
                           => reg_out_1_29_port, A(28) => reg_out_1_28_port, 
                           A(27) => reg_out_1_27_port, A(26) => 
                           reg_out_1_26_port, A(25) => reg_out_1_25_port, A(24)
                           => reg_out_1_24_port, A(23) => reg_out_1_23_port, 
                           A(22) => reg_out_1_22_port, A(21) => 
                           reg_out_1_21_port, A(20) => reg_out_1_20_port, A(19)
                           => reg_out_1_19_port, A(18) => reg_out_1_18_port, 
                           A(17) => reg_out_1_17_port, A(16) => 
                           reg_out_1_16_port, A(15) => reg_out_1_15_port, A(14)
                           => reg_out_1_14_port, A(13) => reg_out_1_13_port, 
                           A(12) => reg_out_1_12_port, A(11) => 
                           reg_out_1_11_port, A(10) => reg_out_1_10_port, A(9) 
                           => reg_out_1_9_port, A(8) => reg_out_1_8_port, A(7) 
                           => reg_out_1_7_port, A(6) => reg_out_1_6_port, A(5) 
                           => reg_out_1_5_port, A(4) => reg_out_1_4_port, A(3) 
                           => reg_out_1_3_port, A(2) => reg_out_1_2_port, A(1) 
                           => reg_out_1_1_port, A(0) => reg_out_1_0_port, B(31)
                           => addends_4_31_port, B(30) => addends_4_30_port, 
                           B(29) => addends_4_29_port, B(28) => 
                           addends_4_28_port, B(27) => addends_4_27_port, B(26)
                           => addends_4_26_port, B(25) => addends_4_25_port, 
                           B(24) => addends_4_24_port, B(23) => 
                           addends_4_23_port, B(22) => addends_4_22_port, B(21)
                           => addends_4_21_port, B(20) => addends_4_20_port, 
                           B(19) => addends_4_19_port, B(18) => 
                           addends_4_18_port, B(17) => addends_4_17_port, B(16)
                           => addends_4_16_port, B(15) => addends_4_15_port, 
                           B(14) => addends_4_14_port, B(13) => 
                           addends_4_13_port, B(12) => addends_4_12_port, B(11)
                           => addends_4_11_port, B(10) => addends_4_10_port, 
                           B(9) => addends_4_9_port, B(8) => addends_4_8_port, 
                           B(7) => addends_4_7_port, B(6) => addends_4_6_port, 
                           B(5) => addends_4_5_port, B(4) => addends_4_4_port, 
                           B(3) => addends_4_3_port, B(2) => addends_4_2_port, 
                           B(1) => addends_4_1_port, B(0) => addends_4_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_1_31_port, S(30) => 
                           add_out_1_30_port, S(29) => add_out_1_29_port, S(28)
                           => add_out_1_28_port, S(27) => add_out_1_27_port, 
                           S(26) => add_out_1_26_port, S(25) => 
                           add_out_1_25_port, S(24) => add_out_1_24_port, S(23)
                           => add_out_1_23_port, S(22) => add_out_1_22_port, 
                           S(21) => add_out_1_21_port, S(20) => 
                           add_out_1_20_port, S(19) => add_out_1_19_port, S(18)
                           => add_out_1_18_port, S(17) => add_out_1_17_port, 
                           S(16) => add_out_1_16_port, S(15) => 
                           add_out_1_15_port, S(14) => add_out_1_14_port, S(13)
                           => add_out_1_13_port, S(12) => add_out_1_12_port, 
                           S(11) => add_out_1_11_port, S(10) => 
                           add_out_1_10_port, S(9) => add_out_1_9_port, S(8) =>
                           add_out_1_8_port, S(7) => add_out_1_7_port, S(6) => 
                           add_out_1_6_port, S(5) => add_out_1_5_port, S(4) => 
                           add_out_1_4_port, S(3) => add_out_1_3_port, S(2) => 
                           add_out_1_2_port, S(1) => add_out_1_1_port, S(0) => 
                           add_out_1_0_port, Cout => n_1524);
   ADD_1i_2 : ADDER_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => 
                           add_out_1_31_port, A(30) => add_out_1_30_port, A(29)
                           => add_out_1_29_port, A(28) => add_out_1_28_port, 
                           A(27) => add_out_1_27_port, A(26) => 
                           add_out_1_26_port, A(25) => add_out_1_25_port, A(24)
                           => add_out_1_24_port, A(23) => add_out_1_23_port, 
                           A(22) => add_out_1_22_port, A(21) => 
                           add_out_1_21_port, A(20) => add_out_1_20_port, A(19)
                           => add_out_1_19_port, A(18) => add_out_1_18_port, 
                           A(17) => add_out_1_17_port, A(16) => 
                           add_out_1_16_port, A(15) => add_out_1_15_port, A(14)
                           => add_out_1_14_port, A(13) => add_out_1_13_port, 
                           A(12) => add_out_1_12_port, A(11) => 
                           add_out_1_11_port, A(10) => add_out_1_10_port, A(9) 
                           => add_out_1_9_port, A(8) => add_out_1_8_port, A(7) 
                           => add_out_1_7_port, A(6) => add_out_1_6_port, A(5) 
                           => add_out_1_5_port, A(4) => add_out_1_4_port, A(3) 
                           => add_out_1_3_port, A(2) => add_out_1_2_port, A(1) 
                           => add_out_1_1_port, A(0) => add_out_1_0_port, B(31)
                           => addends_5_31_port, B(30) => addends_5_30_port, 
                           B(29) => addends_5_29_port, B(28) => 
                           addends_5_28_port, B(27) => addends_5_27_port, B(26)
                           => addends_5_26_port, B(25) => addends_5_25_port, 
                           B(24) => addends_5_24_port, B(23) => 
                           addends_5_23_port, B(22) => addends_5_22_port, B(21)
                           => addends_5_21_port, B(20) => addends_5_20_port, 
                           B(19) => addends_5_19_port, B(18) => 
                           addends_5_18_port, B(17) => addends_5_17_port, B(16)
                           => addends_5_16_port, B(15) => addends_5_15_port, 
                           B(14) => addends_5_14_port, B(13) => 
                           addends_5_13_port, B(12) => addends_5_12_port, B(11)
                           => addends_5_11_port, B(10) => addends_5_10_port, 
                           B(9) => addends_5_9_port, B(8) => addends_5_8_port, 
                           B(7) => addends_5_7_port, B(6) => addends_5_6_port, 
                           B(5) => addends_5_5_port, B(4) => addends_5_4_port, 
                           B(3) => addends_5_3_port, B(2) => addends_5_2_port, 
                           B(1) => addends_5_1_port, B(0) => addends_5_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_2_31_port, S(30) => reg_in_2_30_port
                           , S(29) => reg_in_2_29_port, S(28) => 
                           reg_in_2_28_port, S(27) => reg_in_2_27_port, S(26) 
                           => reg_in_2_26_port, S(25) => reg_in_2_25_port, 
                           S(24) => reg_in_2_24_port, S(23) => reg_in_2_23_port
                           , S(22) => reg_in_2_22_port, S(21) => 
                           reg_in_2_21_port, S(20) => reg_in_2_20_port, S(19) 
                           => reg_in_2_19_port, S(18) => reg_in_2_18_port, 
                           S(17) => reg_in_2_17_port, S(16) => reg_in_2_16_port
                           , S(15) => reg_in_2_15_port, S(14) => 
                           reg_in_2_14_port, S(13) => reg_in_2_13_port, S(12) 
                           => reg_in_2_12_port, S(11) => reg_in_2_11_port, 
                           S(10) => reg_in_2_10_port, S(9) => reg_in_2_9_port, 
                           S(8) => reg_in_2_8_port, S(7) => reg_in_2_7_port, 
                           S(6) => reg_in_2_6_port, S(5) => reg_in_2_5_port, 
                           S(4) => reg_in_2_4_port, S(3) => reg_in_2_3_port, 
                           S(2) => reg_in_2_2_port, S(1) => reg_in_2_1_port, 
                           S(0) => reg_in_2_0_port, Cout => n_1525);
   REG_i_2 : REG_NBIT32_1 port map( clk => CLOCK, reset => X_Logic0_port, 
                           enable => X_Logic1_port, data_in(31) => 
                           reg_in_2_31_port, data_in(30) => reg_in_2_30_port, 
                           data_in(29) => reg_in_2_29_port, data_in(28) => 
                           reg_in_2_28_port, data_in(27) => reg_in_2_27_port, 
                           data_in(26) => reg_in_2_26_port, data_in(25) => 
                           reg_in_2_25_port, data_in(24) => reg_in_2_24_port, 
                           data_in(23) => reg_in_2_23_port, data_in(22) => 
                           reg_in_2_22_port, data_in(21) => reg_in_2_21_port, 
                           data_in(20) => reg_in_2_20_port, data_in(19) => 
                           reg_in_2_19_port, data_in(18) => reg_in_2_18_port, 
                           data_in(17) => reg_in_2_17_port, data_in(16) => 
                           reg_in_2_16_port, data_in(15) => reg_in_2_15_port, 
                           data_in(14) => reg_in_2_14_port, data_in(13) => 
                           reg_in_2_13_port, data_in(12) => reg_in_2_12_port, 
                           data_in(11) => reg_in_2_11_port, data_in(10) => 
                           reg_in_2_10_port, data_in(9) => reg_in_2_9_port, 
                           data_in(8) => reg_in_2_8_port, data_in(7) => 
                           reg_in_2_7_port, data_in(6) => reg_in_2_6_port, 
                           data_in(5) => reg_in_2_5_port, data_in(4) => 
                           reg_in_2_4_port, data_in(3) => reg_in_2_3_port, 
                           data_in(2) => reg_in_2_2_port, data_in(1) => 
                           reg_in_2_1_port, data_in(0) => reg_in_2_0_port, 
                           data_out(31) => reg_out_2_31_port, data_out(30) => 
                           reg_out_2_30_port, data_out(29) => reg_out_2_29_port
                           , data_out(28) => reg_out_2_28_port, data_out(27) =>
                           reg_out_2_27_port, data_out(26) => reg_out_2_26_port
                           , data_out(25) => reg_out_2_25_port, data_out(24) =>
                           reg_out_2_24_port, data_out(23) => reg_out_2_23_port
                           , data_out(22) => reg_out_2_22_port, data_out(21) =>
                           reg_out_2_21_port, data_out(20) => reg_out_2_20_port
                           , data_out(19) => reg_out_2_19_port, data_out(18) =>
                           reg_out_2_18_port, data_out(17) => reg_out_2_17_port
                           , data_out(16) => reg_out_2_16_port, data_out(15) =>
                           reg_out_2_15_port, data_out(14) => reg_out_2_14_port
                           , data_out(13) => reg_out_2_13_port, data_out(12) =>
                           reg_out_2_12_port, data_out(11) => reg_out_2_11_port
                           , data_out(10) => reg_out_2_10_port, data_out(9) => 
                           reg_out_2_9_port, data_out(8) => reg_out_2_8_port, 
                           data_out(7) => reg_out_2_7_port, data_out(6) => 
                           reg_out_2_6_port, data_out(5) => reg_out_2_5_port, 
                           data_out(4) => reg_out_2_4_port, data_out(3) => 
                           reg_out_2_3_port, data_out(2) => reg_out_2_2_port, 
                           data_out(1) => reg_out_2_1_port, data_out(0) => 
                           reg_out_2_0_port);
   ADD_N_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => 
                           reg_out_2_31_port, A(30) => reg_out_2_30_port, A(29)
                           => reg_out_2_29_port, A(28) => reg_out_2_28_port, 
                           A(27) => reg_out_2_27_port, A(26) => 
                           reg_out_2_26_port, A(25) => reg_out_2_25_port, A(24)
                           => reg_out_2_24_port, A(23) => reg_out_2_23_port, 
                           A(22) => reg_out_2_22_port, A(21) => 
                           reg_out_2_21_port, A(20) => reg_out_2_20_port, A(19)
                           => reg_out_2_19_port, A(18) => reg_out_2_18_port, 
                           A(17) => reg_out_2_17_port, A(16) => 
                           reg_out_2_16_port, A(15) => reg_out_2_15_port, A(14)
                           => reg_out_2_14_port, A(13) => reg_out_2_13_port, 
                           A(12) => reg_out_2_12_port, A(11) => 
                           reg_out_2_11_port, A(10) => reg_out_2_10_port, A(9) 
                           => reg_out_2_9_port, A(8) => reg_out_2_8_port, A(7) 
                           => reg_out_2_7_port, A(6) => reg_out_2_6_port, A(5) 
                           => reg_out_2_5_port, A(4) => reg_out_2_4_port, A(3) 
                           => reg_out_2_3_port, A(2) => reg_out_2_2_port, A(1) 
                           => reg_out_2_1_port, A(0) => reg_out_2_0_port, B(31)
                           => addends_6_31_port, B(30) => addends_6_30_port, 
                           B(29) => addends_6_29_port, B(28) => 
                           addends_6_28_port, B(27) => addends_6_27_port, B(26)
                           => addends_6_26_port, B(25) => addends_6_25_port, 
                           B(24) => addends_6_24_port, B(23) => 
                           addends_6_23_port, B(22) => addends_6_22_port, B(21)
                           => addends_6_21_port, B(20) => addends_6_20_port, 
                           B(19) => addends_6_19_port, B(18) => 
                           addends_6_18_port, B(17) => addends_6_17_port, B(16)
                           => addends_6_16_port, B(15) => addends_6_15_port, 
                           B(14) => addends_6_14_port, B(13) => 
                           addends_6_13_port, B(12) => addends_6_12_port, B(11)
                           => addends_6_11_port, B(10) => addends_6_10_port, 
                           B(9) => addends_6_9_port, B(8) => addends_6_8_port, 
                           B(7) => addends_6_7_port, B(6) => addends_6_6_port, 
                           B(5) => addends_6_5_port, B(4) => addends_6_4_port, 
                           B(3) => addends_6_3_port, B(2) => addends_6_2_port, 
                           B(1) => addends_6_1_port, B(0) => addends_6_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_2_31_port, S(30) => 
                           add_out_2_30_port, S(29) => add_out_2_29_port, S(28)
                           => add_out_2_28_port, S(27) => add_out_2_27_port, 
                           S(26) => add_out_2_26_port, S(25) => 
                           add_out_2_25_port, S(24) => add_out_2_24_port, S(23)
                           => add_out_2_23_port, S(22) => add_out_2_22_port, 
                           S(21) => add_out_2_21_port, S(20) => 
                           add_out_2_20_port, S(19) => add_out_2_19_port, S(18)
                           => add_out_2_18_port, S(17) => add_out_2_17_port, 
                           S(16) => add_out_2_16_port, S(15) => 
                           add_out_2_15_port, S(14) => add_out_2_14_port, S(13)
                           => add_out_2_13_port, S(12) => add_out_2_12_port, 
                           S(11) => add_out_2_11_port, S(10) => 
                           add_out_2_10_port, S(9) => add_out_2_9_port, S(8) =>
                           add_out_2_8_port, S(7) => add_out_2_7_port, S(6) => 
                           add_out_2_6_port, S(5) => add_out_2_5_port, S(4) => 
                           add_out_2_4_port, S(3) => add_out_2_3_port, S(2) => 
                           add_out_2_2_port, S(1) => add_out_2_1_port, S(0) => 
                           add_out_2_0_port, Cout => n_1526);
   ADD_N : ADDER_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => add_out_2_31_port,
                           A(30) => add_out_2_30_port, A(29) => 
                           add_out_2_29_port, A(28) => add_out_2_28_port, A(27)
                           => add_out_2_27_port, A(26) => add_out_2_26_port, 
                           A(25) => add_out_2_25_port, A(24) => 
                           add_out_2_24_port, A(23) => add_out_2_23_port, A(22)
                           => add_out_2_22_port, A(21) => add_out_2_21_port, 
                           A(20) => add_out_2_20_port, A(19) => 
                           add_out_2_19_port, A(18) => add_out_2_18_port, A(17)
                           => add_out_2_17_port, A(16) => add_out_2_16_port, 
                           A(15) => add_out_2_15_port, A(14) => 
                           add_out_2_14_port, A(13) => add_out_2_13_port, A(12)
                           => add_out_2_12_port, A(11) => add_out_2_11_port, 
                           A(10) => add_out_2_10_port, A(9) => add_out_2_9_port
                           , A(8) => add_out_2_8_port, A(7) => add_out_2_7_port
                           , A(6) => add_out_2_6_port, A(5) => add_out_2_5_port
                           , A(4) => add_out_2_4_port, A(3) => add_out_2_3_port
                           , A(2) => add_out_2_2_port, A(1) => add_out_2_1_port
                           , A(0) => add_out_2_0_port, B(31) => 
                           addends_7_31_port, B(30) => addends_7_30_port, B(29)
                           => addends_7_29_port, B(28) => addends_7_28_port, 
                           B(27) => addends_7_27_port, B(26) => 
                           addends_7_26_port, B(25) => addends_7_25_port, B(24)
                           => addends_7_24_port, B(23) => addends_7_23_port, 
                           B(22) => addends_7_22_port, B(21) => 
                           addends_7_21_port, B(20) => addends_7_20_port, B(19)
                           => addends_7_19_port, B(18) => addends_7_18_port, 
                           B(17) => addends_7_17_port, B(16) => 
                           addends_7_16_port, B(15) => addends_7_15_port, B(14)
                           => addends_7_14_port, B(13) => addends_7_13_port, 
                           B(12) => addends_7_12_port, B(11) => 
                           addends_7_11_port, B(10) => addends_7_10_port, B(9) 
                           => addends_7_9_port, B(8) => addends_7_8_port, B(7) 
                           => addends_7_7_port, B(6) => addends_7_6_port, B(5) 
                           => addends_7_5_port, B(4) => addends_7_4_port, B(3) 
                           => addends_7_3_port, B(2) => addends_7_2_port, B(1) 
                           => addends_7_1_port, B(0) => addends_7_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => Y(31), S(30) => Y(30), S(29) => Y(29), 
                           S(28) => Y(28), S(27) => Y(27), S(26) => Y(26), 
                           S(25) => Y(25), S(24) => Y(24), S(23) => Y(23), 
                           S(22) => Y(22), S(21) => Y(21), S(20) => Y(20), 
                           S(19) => Y(19), S(18) => Y(18), S(17) => Y(17), 
                           S(16) => Y(16), S(15) => Y(15), S(14) => Y(14), 
                           S(13) => Y(13), S(12) => Y(12), S(11) => Y(11), 
                           S(10) => Y(10), S(9) => Y(9), S(8) => Y(8), S(7) => 
                           Y(7), S(6) => Y(6), S(5) => Y(5), S(4) => Y(4), S(3)
                           => Y(3), S(2) => Y(2), S(1) => Y(1), S(0) => Y(0), 
                           Cout => n_1527);
   U3 : XNOR2_X2 port map( A => n72, B => A(8), ZN => A_neg_9_17_port);
   U4 : XNOR2_X2 port map( A => n74, B => A(14), ZN => A_neg_9_23_port);
   U6 : XNOR2_X2 port map( A => n73, B => A(12), ZN => A_neg_9_21_port);
   U7 : XNOR2_X2 port map( A => n71, B => A(4), ZN => A_neg_9_13_port);
   U9 : XNOR2_X2 port map( A => n70, B => A(2), ZN => A_neg_9_11_port);
   U10 : XOR2_X2 port map( A => n7, B => A(7), Z => A_neg_9_16_port);
   U11 : XOR2_X2 port map( A => n14, B => A(13), Z => A_neg_9_22_port);
   U12 : XOR2_X2 port map( A => n16, B => A(11), Z => A_neg_9_20_port);
   U13 : XOR2_X2 port map( A => n5, B => A(9), Z => A_neg_9_18_port);
   U14 : XOR2_X2 port map( A => n8, B => A(6), Z => A_neg_9_15_port);
   U15 : XOR2_X2 port map( A => n12, B => A(3), Z => A_neg_9_12_port);
   U16 : XOR2_X2 port map( A => A(1), B => n96, Z => A_neg_9_10_port);
   U17 : BUF_X1 port map( A => n75, Z => n91);
   U18 : BUF_X1 port map( A => n75, Z => n92);
   U19 : BUF_X1 port map( A => n75, Z => n90);
   U20 : BUF_X1 port map( A => n77, Z => n75);
   U21 : BUF_X1 port map( A => n76, Z => n93);
   U22 : BUF_X1 port map( A => A(0), Z => n97);
   U23 : BUF_X1 port map( A => n92, Z => n83);
   U24 : BUF_X1 port map( A => n92, Z => n81);
   U25 : BUF_X1 port map( A => n92, Z => n82);
   U26 : BUF_X1 port map( A => n91, Z => n84);
   U27 : BUF_X1 port map( A => n91, Z => n85);
   U28 : BUF_X1 port map( A => n91, Z => n86);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n90, Z => n89);
   U32 : BUF_X1 port map( A => n93, Z => n80);
   U33 : BUF_X1 port map( A => n93, Z => n79);
   U34 : BUF_X1 port map( A => n93, Z => n78);
   U35 : BUF_X1 port map( A => n77, Z => n76);
   U36 : NOR2_X1 port map( A1 => n96, A2 => A(1), ZN => n70);
   U37 : NOR2_X1 port map( A1 => n12, A2 => A(3), ZN => n71);
   U38 : NOR2_X1 port map( A1 => n7, A2 => A(7), ZN => n72);
   U39 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n73);
   U40 : NOR2_X1 port map( A1 => n14, A2 => A(13), ZN => n74);
   U41 : OAI21_X2 port map( B1 => n18, B2 => n99, A => n19, ZN => 
                           A_neg_9_19_port);
   U42 : OAI21_X1 port map( B1 => A(9), B2 => n5, A => n99, ZN => n19);
   U43 : INV_X1 port map( A => A(10), ZN => n99);
   U44 : NOR3_X1 port map( A1 => A(3), A2 => A(4), A3 => n12, ZN => n10);
   U45 : NOR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n14, ZN => n4);
   U46 : NAND2_X1 port map( A1 => n10, A2 => n100, ZN => n8);
   U47 : INV_X1 port map( A => A(5), ZN => n100);
   U48 : OR2_X1 port map( A1 => n5, A2 => A(9), ZN => n18);
   U49 : OR2_X1 port map( A1 => n18, A2 => A(10), ZN => n16);
   U50 : OR2_X1 port map( A1 => n8, A2 => A(6), ZN => n7);
   U51 : OR3_X1 port map( A1 => A(11), A2 => A(12), A3 => n16, ZN => n14);
   U52 : OR3_X1 port map( A1 => A(2), A2 => n94, A3 => A(1), ZN => n12);
   U53 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n7, ZN => n5);
   U54 : BUF_X1 port map( A => n9, Z => n77);
   U55 : NAND2_X1 port map( A1 => n4, A2 => n98, ZN => n9);
   U56 : INV_X1 port map( A => A(15), ZN => n98);
   U57 : BUF_X1 port map( A => n97, Z => n94);
   U58 : BUF_X1 port map( A => n97, Z => n95);
   U59 : BUF_X1 port map( A => n97, Z => n96);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CMP_NBIT32 is

   port( SUM : in std_logic_vector (31 downto 0);  Cout : in std_logic;  A_L_B,
         A_LE_B, A_G_B, A_GE_B, A_E_B, A_NE_B : out std_logic);

end CMP_NBIT32;

architecture SYN_structural of CMP_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal A_L_B_port, A_LE_B_port, N29, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      A_E_B_port : std_logic;

begin
   A_L_B <= A_L_B_port;
   A_LE_B <= A_LE_B_port;
   A_E_B <= A_E_B_port;
   A_NE_B <= N29;
   
   U1 : NOR2_X1 port map( A1 => Cout, A2 => A_E_B_port, ZN => A_L_B_port);
   U2 : NAND2_X1 port map( A1 => Cout, A2 => N29, ZN => A_LE_B_port);
   U3 : INV_X1 port map( A => N29, ZN => A_E_B_port);
   U4 : NAND4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => N29);
   U5 : AND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n7);
   U6 : NOR4_X1 port map( A1 => SUM(19), A2 => SUM(18), A3 => SUM(17), A4 => 
                           SUM(16), ZN => n4);
   U7 : NOR4_X1 port map( A1 => SUM(22), A2 => SUM(21), A3 => SUM(20), A4 => 
                           SUM(1), ZN => n5);
   U8 : NOR4_X1 port map( A1 => SUM(9), A2 => SUM(8), A3 => SUM(7), A4 => 
                           SUM(6), ZN => n11);
   U9 : NOR4_X1 port map( A1 => SUM(5), A2 => SUM(4), A3 => SUM(3), A4 => 
                           SUM(30), ZN => n10);
   U10 : NOR4_X1 port map( A1 => n12, A2 => SUM(0), A3 => SUM(11), A4 => 
                           SUM(10), ZN => n6);
   U11 : NOR4_X1 port map( A1 => SUM(2), A2 => SUM(29), A3 => SUM(28), A4 => 
                           SUM(27), ZN => n9);
   U12 : NOR4_X1 port map( A1 => SUM(26), A2 => SUM(25), A3 => SUM(24), A4 => 
                           SUM(23), ZN => n8);
   U13 : OR4_X1 port map( A1 => SUM(13), A2 => SUM(12), A3 => SUM(15), A4 => 
                           SUM(14), ZN => n12);
   U14 : INV_X1 port map( A => A_LE_B_port, ZN => A_G_B);
   U15 : INV_X1 port map( A => A_L_B_port, ZN => A_GE_B);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LOGIC_NBIT32_N_SELECTOR4 is

   port( S : in std_logic_vector (3 downto 0);  A, B : in std_logic_vector (31 
         downto 0);  O : out std_logic_vector (31 downto 0));

end LOGIC_NBIT32_N_SELECTOR4;

architecture SYN_structural of LOGIC_NBIT32_N_SELECTOR4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4_1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_2
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_3
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_4
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_2
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_5
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_6
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_7
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_8
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_3
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_9
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_10
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_11
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_12
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_4
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_13
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_14
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_15
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_16
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_5
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_17
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_18
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_19
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_20
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_6
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_21
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_22
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_23
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_24
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_7
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_25
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_26
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_27
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_28
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_8
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_29
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_30
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_31
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_32
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_9
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_33
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_34
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_35
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_36
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_10
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_37
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_38
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_39
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_40
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_11
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_41
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_42
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_43
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_44
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_12
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_45
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_46
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_47
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_48
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_13
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_49
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_50
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_51
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_52
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_14
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_53
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_54
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_55
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_56
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_15
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_57
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_58
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_59
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_60
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_16
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_61
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_62
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_63
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_64
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_17
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_65
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_66
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_67
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_68
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_18
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_69
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_70
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_71
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_72
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_19
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_73
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_74
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_75
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_76
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_20
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_77
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_78
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_79
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_80
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_21
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_81
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_82
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_83
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_84
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_22
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_85
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_86
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_87
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_88
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_23
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_89
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_90
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_91
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_92
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_24
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_93
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_94
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_95
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_96
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_25
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_97
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_98
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_99
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_100
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_26
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_101
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_102
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_103
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_104
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_27
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_105
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_106
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_107
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_108
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_28
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_109
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_110
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_111
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_112
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_29
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_113
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_114
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_115
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_116
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_30
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_117
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_118
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_119
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_120
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_31
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_121
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_122
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_123
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_124
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_0
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_125
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_126
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_127
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_0
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal An_31_port, An_30_port, An_29_port, An_28_port, An_27_port, 
      An_26_port, An_25_port, An_24_port, An_23_port, An_22_port, An_21_port, 
      An_20_port, An_19_port, An_18_port, An_17_port, An_16_port, An_15_port, 
      An_14_port, An_13_port, An_12_port, An_11_port, An_10_port, An_9_port, 
      An_8_port, An_7_port, An_6_port, An_5_port, An_4_port, An_3_port, 
      An_2_port, An_1_port, An_0_port, Bn_31_port, Bn_30_port, Bn_29_port, 
      Bn_28_port, Bn_27_port, Bn_26_port, Bn_25_port, Bn_24_port, Bn_23_port, 
      Bn_22_port, Bn_21_port, Bn_20_port, Bn_19_port, Bn_18_port, Bn_17_port, 
      Bn_16_port, Bn_15_port, Bn_14_port, Bn_13_port, Bn_12_port, Bn_11_port, 
      Bn_10_port, Bn_9_port, Bn_8_port, Bn_7_port, Bn_6_port, Bn_5_port, 
      Bn_4_port, Bn_3_port, Bn_2_port, Bn_1_port, Bn_0_port, l0_31_port, 
      l0_30_port, l0_29_port, l0_28_port, l0_27_port, l0_26_port, l0_25_port, 
      l0_24_port, l0_23_port, l0_22_port, l0_21_port, l0_20_port, l0_19_port, 
      l0_18_port, l0_17_port, l0_16_port, l0_15_port, l0_14_port, l0_13_port, 
      l0_12_port, l0_11_port, l0_10_port, l0_9_port, l0_8_port, l0_7_port, 
      l0_6_port, l0_5_port, l0_4_port, l0_3_port, l0_2_port, l0_1_port, 
      l0_0_port, l1_31_port, l1_30_port, l1_29_port, l1_28_port, l1_27_port, 
      l1_26_port, l1_25_port, l1_24_port, l1_23_port, l1_22_port, l1_21_port, 
      l1_20_port, l1_19_port, l1_18_port, l1_17_port, l1_16_port, l1_15_port, 
      l1_14_port, l1_13_port, l1_12_port, l1_11_port, l1_10_port, l1_9_port, 
      l1_8_port, l1_7_port, l1_6_port, l1_5_port, l1_4_port, l1_3_port, 
      l1_2_port, l1_1_port, l1_0_port, l2_31_port, l2_30_port, l2_29_port, 
      l2_28_port, l2_27_port, l2_26_port, l2_25_port, l2_24_port, l2_23_port, 
      l2_22_port, l2_21_port, l2_20_port, l2_19_port, l2_18_port, l2_17_port, 
      l2_16_port, l2_15_port, l2_14_port, l2_13_port, l2_12_port, l2_11_port, 
      l2_10_port, l2_9_port, l2_8_port, l2_7_port, l2_6_port, l2_5_port, 
      l2_4_port, l2_3_port, l2_2_port, l2_1_port, l2_0_port, l3_31_port, 
      l3_30_port, l3_29_port, l3_28_port, l3_27_port, l3_26_port, l3_25_port, 
      l3_24_port, l3_23_port, l3_22_port, l3_21_port, l3_20_port, l3_19_port, 
      l3_18_port, l3_17_port, l3_16_port, l3_15_port, l3_14_port, l3_13_port, 
      l3_12_port, l3_11_port, l3_10_port, l3_9_port, l3_8_port, l3_7_port, 
      l3_6_port, l3_5_port, l3_4_port, l3_3_port, l3_2_port, l3_1_port, 
      l3_0_port, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32 : std_logic;

begin
   
   A_i_0 : IV_0 port map( A => A(0), Y => An_0_port);
   A_i_1 : IV_63 port map( A => A(1), Y => An_1_port);
   A_i_2 : IV_62 port map( A => A(2), Y => An_2_port);
   A_i_3 : IV_61 port map( A => A(3), Y => An_3_port);
   A_i_4 : IV_60 port map( A => A(4), Y => An_4_port);
   A_i_5 : IV_59 port map( A => A(5), Y => An_5_port);
   A_i_6 : IV_58 port map( A => A(6), Y => An_6_port);
   A_i_7 : IV_57 port map( A => A(7), Y => An_7_port);
   A_i_8 : IV_56 port map( A => A(8), Y => An_8_port);
   A_i_9 : IV_55 port map( A => A(9), Y => An_9_port);
   A_i_10 : IV_54 port map( A => A(10), Y => An_10_port);
   A_i_11 : IV_53 port map( A => A(11), Y => An_11_port);
   A_i_12 : IV_52 port map( A => A(12), Y => An_12_port);
   A_i_13 : IV_51 port map( A => A(13), Y => An_13_port);
   A_i_14 : IV_50 port map( A => A(14), Y => An_14_port);
   A_i_15 : IV_49 port map( A => A(15), Y => An_15_port);
   A_i_16 : IV_48 port map( A => A(16), Y => An_16_port);
   A_i_17 : IV_47 port map( A => A(17), Y => An_17_port);
   A_i_18 : IV_46 port map( A => A(18), Y => An_18_port);
   A_i_19 : IV_45 port map( A => A(19), Y => An_19_port);
   A_i_20 : IV_44 port map( A => A(20), Y => An_20_port);
   A_i_21 : IV_43 port map( A => A(21), Y => An_21_port);
   A_i_22 : IV_42 port map( A => A(22), Y => An_22_port);
   A_i_23 : IV_41 port map( A => A(23), Y => An_23_port);
   A_i_24 : IV_40 port map( A => A(24), Y => An_24_port);
   A_i_25 : IV_39 port map( A => A(25), Y => An_25_port);
   A_i_26 : IV_38 port map( A => A(26), Y => An_26_port);
   A_i_27 : IV_37 port map( A => A(27), Y => An_27_port);
   A_i_28 : IV_36 port map( A => A(28), Y => An_28_port);
   A_i_29 : IV_35 port map( A => A(29), Y => An_29_port);
   A_i_30 : IV_34 port map( A => A(30), Y => An_30_port);
   A_i_31 : IV_33 port map( A => A(31), Y => An_31_port);
   B_i_0 : IV_32 port map( A => B(0), Y => Bn_0_port);
   B_i_1 : IV_31 port map( A => B(1), Y => Bn_1_port);
   B_i_2 : IV_30 port map( A => B(2), Y => Bn_2_port);
   B_i_3 : IV_29 port map( A => B(3), Y => Bn_3_port);
   B_i_4 : IV_28 port map( A => B(4), Y => Bn_4_port);
   B_i_5 : IV_27 port map( A => B(5), Y => Bn_5_port);
   B_i_6 : IV_26 port map( A => B(6), Y => Bn_6_port);
   B_i_7 : IV_25 port map( A => B(7), Y => Bn_7_port);
   B_i_8 : IV_24 port map( A => B(8), Y => Bn_8_port);
   B_i_9 : IV_23 port map( A => B(9), Y => Bn_9_port);
   B_i_10 : IV_22 port map( A => B(10), Y => Bn_10_port);
   B_i_11 : IV_21 port map( A => B(11), Y => Bn_11_port);
   B_i_12 : IV_20 port map( A => B(12), Y => Bn_12_port);
   B_i_13 : IV_19 port map( A => B(13), Y => Bn_13_port);
   B_i_14 : IV_18 port map( A => B(14), Y => Bn_14_port);
   B_i_15 : IV_17 port map( A => B(15), Y => Bn_15_port);
   B_i_16 : IV_16 port map( A => B(16), Y => Bn_16_port);
   B_i_17 : IV_15 port map( A => B(17), Y => Bn_17_port);
   B_i_18 : IV_14 port map( A => B(18), Y => Bn_18_port);
   B_i_19 : IV_13 port map( A => B(19), Y => Bn_19_port);
   B_i_20 : IV_12 port map( A => B(20), Y => Bn_20_port);
   B_i_21 : IV_11 port map( A => B(21), Y => Bn_21_port);
   B_i_22 : IV_10 port map( A => B(22), Y => Bn_22_port);
   B_i_23 : IV_9 port map( A => B(23), Y => Bn_23_port);
   B_i_24 : IV_8 port map( A => B(24), Y => Bn_24_port);
   B_i_25 : IV_7 port map( A => B(25), Y => Bn_25_port);
   B_i_26 : IV_6 port map( A => B(26), Y => Bn_26_port);
   B_i_27 : IV_5 port map( A => B(27), Y => Bn_27_port);
   B_i_28 : IV_4 port map( A => B(28), Y => Bn_28_port);
   B_i_29 : IV_3 port map( A => B(29), Y => Bn_29_port);
   B_i_30 : IV_2 port map( A => B(30), Y => Bn_30_port);
   B_i_31 : IV_1 port map( A => B(31), Y => Bn_31_port);
   U0_0 : ND3_0 port map( A => n19, B => An_0_port, C => Bn_0_port, Y => 
                           l0_0_port);
   U1_0 : ND3_127 port map( A => n21, B => An_0_port, C => B(0), Y => l1_0_port
                           );
   U2_0 : ND3_126 port map( A => n25, B => A(0), C => Bn_0_port, Y => l2_0_port
                           );
   U3_0 : ND3_125 port map( A => n29, B => A(0), C => B(0), Y => l3_0_port);
   U4_0 : ND4_0 port map( A => l0_0_port, B => l1_0_port, C => l2_0_port, D => 
                           l3_0_port, Y => O(0));
   U0_1 : ND3_124 port map( A => n17, B => An_1_port, C => Bn_1_port, Y => 
                           l0_1_port);
   U1_1 : ND3_123 port map( A => n21, B => An_1_port, C => B(1), Y => l1_1_port
                           );
   U2_1 : ND3_122 port map( A => n25, B => A(1), C => Bn_1_port, Y => l2_1_port
                           );
   U3_1 : ND3_121 port map( A => n29, B => A(1), C => B(1), Y => l3_1_port);
   U4_1 : ND4_31 port map( A => l0_1_port, B => l1_1_port, C => l2_1_port, D =>
                           l3_1_port, Y => O(1));
   U0_2 : ND3_120 port map( A => n17, B => An_2_port, C => Bn_2_port, Y => 
                           l0_2_port);
   U1_2 : ND3_119 port map( A => n21, B => An_2_port, C => B(2), Y => l1_2_port
                           );
   U2_2 : ND3_118 port map( A => n25, B => A(2), C => Bn_2_port, Y => l2_2_port
                           );
   U3_2 : ND3_117 port map( A => n29, B => A(2), C => B(2), Y => l3_2_port);
   U4_2 : ND4_30 port map( A => l0_2_port, B => l1_2_port, C => l2_2_port, D =>
                           l3_2_port, Y => O(2));
   U0_3 : ND3_116 port map( A => n17, B => An_3_port, C => Bn_3_port, Y => 
                           l0_3_port);
   U1_3 : ND3_115 port map( A => n21, B => An_3_port, C => B(3), Y => l1_3_port
                           );
   U2_3 : ND3_114 port map( A => n25, B => A(3), C => Bn_3_port, Y => l2_3_port
                           );
   U3_3 : ND3_113 port map( A => n29, B => A(3), C => B(3), Y => l3_3_port);
   U4_3 : ND4_29 port map( A => l0_3_port, B => l1_3_port, C => l2_3_port, D =>
                           l3_3_port, Y => O(3));
   U0_4 : ND3_112 port map( A => n17, B => An_4_port, C => Bn_4_port, Y => 
                           l0_4_port);
   U1_4 : ND3_111 port map( A => n21, B => An_4_port, C => B(4), Y => l1_4_port
                           );
   U2_4 : ND3_110 port map( A => n25, B => A(4), C => Bn_4_port, Y => l2_4_port
                           );
   U3_4 : ND3_109 port map( A => n29, B => A(4), C => B(4), Y => l3_4_port);
   U4_4 : ND4_28 port map( A => l0_4_port, B => l1_4_port, C => l2_4_port, D =>
                           l3_4_port, Y => O(4));
   U0_5 : ND3_108 port map( A => n17, B => An_5_port, C => Bn_5_port, Y => 
                           l0_5_port);
   U1_5 : ND3_107 port map( A => n21, B => An_5_port, C => B(5), Y => l1_5_port
                           );
   U2_5 : ND3_106 port map( A => n25, B => A(5), C => Bn_5_port, Y => l2_5_port
                           );
   U3_5 : ND3_105 port map( A => n29, B => A(5), C => B(5), Y => l3_5_port);
   U4_5 : ND4_27 port map( A => l0_5_port, B => l1_5_port, C => l2_5_port, D =>
                           l3_5_port, Y => O(5));
   U0_6 : ND3_104 port map( A => n17, B => An_6_port, C => Bn_6_port, Y => 
                           l0_6_port);
   U1_6 : ND3_103 port map( A => n21, B => An_6_port, C => B(6), Y => l1_6_port
                           );
   U2_6 : ND3_102 port map( A => n25, B => A(6), C => Bn_6_port, Y => l2_6_port
                           );
   U3_6 : ND3_101 port map( A => n29, B => A(6), C => B(6), Y => l3_6_port);
   U4_6 : ND4_26 port map( A => l0_6_port, B => l1_6_port, C => l2_6_port, D =>
                           l3_6_port, Y => O(6));
   U0_7 : ND3_100 port map( A => n17, B => An_7_port, C => Bn_7_port, Y => 
                           l0_7_port);
   U1_7 : ND3_99 port map( A => n21, B => An_7_port, C => B(7), Y => l1_7_port)
                           ;
   U2_7 : ND3_98 port map( A => n25, B => A(7), C => Bn_7_port, Y => l2_7_port)
                           ;
   U3_7 : ND3_97 port map( A => n29, B => A(7), C => B(7), Y => l3_7_port);
   U4_7 : ND4_25 port map( A => l0_7_port, B => l1_7_port, C => l2_7_port, D =>
                           l3_7_port, Y => O(7));
   U0_8 : ND3_96 port map( A => n17, B => An_8_port, C => Bn_8_port, Y => 
                           l0_8_port);
   U1_8 : ND3_95 port map( A => n21, B => An_8_port, C => B(8), Y => l1_8_port)
                           ;
   U2_8 : ND3_94 port map( A => n25, B => A(8), C => Bn_8_port, Y => l2_8_port)
                           ;
   U3_8 : ND3_93 port map( A => n29, B => A(8), C => B(8), Y => l3_8_port);
   U4_8 : ND4_24 port map( A => l0_8_port, B => l1_8_port, C => l2_8_port, D =>
                           l3_8_port, Y => O(8));
   U0_9 : ND3_92 port map( A => n17, B => An_9_port, C => Bn_9_port, Y => 
                           l0_9_port);
   U1_9 : ND3_91 port map( A => n21, B => An_9_port, C => B(9), Y => l1_9_port)
                           ;
   U2_9 : ND3_90 port map( A => n25, B => A(9), C => Bn_9_port, Y => l2_9_port)
                           ;
   U3_9 : ND3_89 port map( A => n29, B => A(9), C => B(9), Y => l3_9_port);
   U4_9 : ND4_23 port map( A => l0_9_port, B => l1_9_port, C => l2_9_port, D =>
                           l3_9_port, Y => O(9));
   U0_10 : ND3_88 port map( A => n17, B => An_10_port, C => Bn_10_port, Y => 
                           l0_10_port);
   U1_10 : ND3_87 port map( A => n21, B => An_10_port, C => B(10), Y => 
                           l1_10_port);
   U2_10 : ND3_86 port map( A => n25, B => A(10), C => Bn_10_port, Y => 
                           l2_10_port);
   U3_10 : ND3_85 port map( A => n29, B => A(10), C => B(10), Y => l3_10_port);
   U4_10 : ND4_22 port map( A => l0_10_port, B => l1_10_port, C => l2_10_port, 
                           D => l3_10_port, Y => O(10));
   U0_11 : ND3_84 port map( A => n17, B => An_11_port, C => Bn_11_port, Y => 
                           l0_11_port);
   U1_11 : ND3_83 port map( A => n21, B => An_11_port, C => B(11), Y => 
                           l1_11_port);
   U2_11 : ND3_82 port map( A => n25, B => A(11), C => Bn_11_port, Y => 
                           l2_11_port);
   U3_11 : ND3_81 port map( A => n29, B => A(11), C => B(11), Y => l3_11_port);
   U4_11 : ND4_21 port map( A => l0_11_port, B => l1_11_port, C => l2_11_port, 
                           D => l3_11_port, Y => O(11));
   U0_12 : ND3_80 port map( A => n17, B => An_12_port, C => Bn_12_port, Y => 
                           l0_12_port);
   U1_12 : ND3_79 port map( A => n22, B => An_12_port, C => B(12), Y => 
                           l1_12_port);
   U2_12 : ND3_78 port map( A => n26, B => A(12), C => Bn_12_port, Y => 
                           l2_12_port);
   U3_12 : ND3_77 port map( A => n30, B => A(12), C => B(12), Y => l3_12_port);
   U4_12 : ND4_20 port map( A => l0_12_port, B => l1_12_port, C => l2_12_port, 
                           D => l3_12_port, Y => O(12));
   U0_13 : ND3_76 port map( A => n18, B => An_13_port, C => Bn_13_port, Y => 
                           l0_13_port);
   U1_13 : ND3_75 port map( A => n22, B => An_13_port, C => B(13), Y => 
                           l1_13_port);
   U2_13 : ND3_74 port map( A => n26, B => A(13), C => Bn_13_port, Y => 
                           l2_13_port);
   U3_13 : ND3_73 port map( A => n30, B => A(13), C => B(13), Y => l3_13_port);
   U4_13 : ND4_19 port map( A => l0_13_port, B => l1_13_port, C => l2_13_port, 
                           D => l3_13_port, Y => O(13));
   U0_14 : ND3_72 port map( A => n18, B => An_14_port, C => Bn_14_port, Y => 
                           l0_14_port);
   U1_14 : ND3_71 port map( A => n22, B => An_14_port, C => B(14), Y => 
                           l1_14_port);
   U2_14 : ND3_70 port map( A => n26, B => A(14), C => Bn_14_port, Y => 
                           l2_14_port);
   U3_14 : ND3_69 port map( A => n30, B => A(14), C => B(14), Y => l3_14_port);
   U4_14 : ND4_18 port map( A => l0_14_port, B => l1_14_port, C => l2_14_port, 
                           D => l3_14_port, Y => O(14));
   U0_15 : ND3_68 port map( A => n18, B => An_15_port, C => Bn_15_port, Y => 
                           l0_15_port);
   U1_15 : ND3_67 port map( A => n22, B => An_15_port, C => B(15), Y => 
                           l1_15_port);
   U2_15 : ND3_66 port map( A => n26, B => A(15), C => Bn_15_port, Y => 
                           l2_15_port);
   U3_15 : ND3_65 port map( A => n30, B => A(15), C => B(15), Y => l3_15_port);
   U4_15 : ND4_17 port map( A => l0_15_port, B => l1_15_port, C => l2_15_port, 
                           D => l3_15_port, Y => O(15));
   U0_16 : ND3_64 port map( A => n18, B => An_16_port, C => Bn_16_port, Y => 
                           l0_16_port);
   U1_16 : ND3_63 port map( A => n22, B => An_16_port, C => B(16), Y => 
                           l1_16_port);
   U2_16 : ND3_62 port map( A => n26, B => A(16), C => Bn_16_port, Y => 
                           l2_16_port);
   U3_16 : ND3_61 port map( A => n30, B => A(16), C => B(16), Y => l3_16_port);
   U4_16 : ND4_16 port map( A => l0_16_port, B => l1_16_port, C => l2_16_port, 
                           D => l3_16_port, Y => O(16));
   U0_17 : ND3_60 port map( A => n18, B => An_17_port, C => Bn_17_port, Y => 
                           l0_17_port);
   U1_17 : ND3_59 port map( A => n22, B => An_17_port, C => B(17), Y => 
                           l1_17_port);
   U2_17 : ND3_58 port map( A => n26, B => A(17), C => Bn_17_port, Y => 
                           l2_17_port);
   U3_17 : ND3_57 port map( A => n30, B => A(17), C => B(17), Y => l3_17_port);
   U4_17 : ND4_15 port map( A => l0_17_port, B => l1_17_port, C => l2_17_port, 
                           D => l3_17_port, Y => O(17));
   U0_18 : ND3_56 port map( A => n18, B => An_18_port, C => Bn_18_port, Y => 
                           l0_18_port);
   U1_18 : ND3_55 port map( A => n22, B => An_18_port, C => B(18), Y => 
                           l1_18_port);
   U2_18 : ND3_54 port map( A => n26, B => A(18), C => Bn_18_port, Y => 
                           l2_18_port);
   U3_18 : ND3_53 port map( A => n30, B => A(18), C => B(18), Y => l3_18_port);
   U4_18 : ND4_14 port map( A => l0_18_port, B => l1_18_port, C => l2_18_port, 
                           D => l3_18_port, Y => O(18));
   U0_19 : ND3_52 port map( A => n18, B => An_19_port, C => Bn_19_port, Y => 
                           l0_19_port);
   U1_19 : ND3_51 port map( A => n22, B => An_19_port, C => B(19), Y => 
                           l1_19_port);
   U2_19 : ND3_50 port map( A => n26, B => A(19), C => Bn_19_port, Y => 
                           l2_19_port);
   U3_19 : ND3_49 port map( A => n30, B => A(19), C => B(19), Y => l3_19_port);
   U4_19 : ND4_13 port map( A => l0_19_port, B => l1_19_port, C => l2_19_port, 
                           D => l3_19_port, Y => O(19));
   U0_20 : ND3_48 port map( A => n18, B => An_20_port, C => Bn_20_port, Y => 
                           l0_20_port);
   U1_20 : ND3_47 port map( A => n22, B => An_20_port, C => B(20), Y => 
                           l1_20_port);
   U2_20 : ND3_46 port map( A => n26, B => A(20), C => Bn_20_port, Y => 
                           l2_20_port);
   U3_20 : ND3_45 port map( A => n30, B => A(20), C => B(20), Y => l3_20_port);
   U4_20 : ND4_12 port map( A => l0_20_port, B => l1_20_port, C => l2_20_port, 
                           D => l3_20_port, Y => O(20));
   U0_21 : ND3_44 port map( A => n18, B => An_21_port, C => Bn_21_port, Y => 
                           l0_21_port);
   U1_21 : ND3_43 port map( A => n22, B => An_21_port, C => B(21), Y => 
                           l1_21_port);
   U2_21 : ND3_42 port map( A => n26, B => A(21), C => Bn_21_port, Y => 
                           l2_21_port);
   U3_21 : ND3_41 port map( A => n30, B => A(21), C => B(21), Y => l3_21_port);
   U4_21 : ND4_11 port map( A => l0_21_port, B => l1_21_port, C => l2_21_port, 
                           D => l3_21_port, Y => O(21));
   U0_22 : ND3_40 port map( A => n18, B => An_22_port, C => Bn_22_port, Y => 
                           l0_22_port);
   U1_22 : ND3_39 port map( A => n22, B => An_22_port, C => B(22), Y => 
                           l1_22_port);
   U2_22 : ND3_38 port map( A => n26, B => A(22), C => Bn_22_port, Y => 
                           l2_22_port);
   U3_22 : ND3_37 port map( A => n30, B => A(22), C => B(22), Y => l3_22_port);
   U4_22 : ND4_10 port map( A => l0_22_port, B => l1_22_port, C => l2_22_port, 
                           D => l3_22_port, Y => O(22));
   U0_23 : ND3_36 port map( A => n18, B => An_23_port, C => Bn_23_port, Y => 
                           l0_23_port);
   U1_23 : ND3_35 port map( A => n22, B => An_23_port, C => B(23), Y => 
                           l1_23_port);
   U2_23 : ND3_34 port map( A => n26, B => A(23), C => Bn_23_port, Y => 
                           l2_23_port);
   U3_23 : ND3_33 port map( A => n30, B => A(23), C => B(23), Y => l3_23_port);
   U4_23 : ND4_9 port map( A => l0_23_port, B => l1_23_port, C => l2_23_port, D
                           => l3_23_port, Y => O(23));
   U0_24 : ND3_32 port map( A => n18, B => An_24_port, C => Bn_24_port, Y => 
                           l0_24_port);
   U1_24 : ND3_31 port map( A => n23, B => An_24_port, C => B(24), Y => 
                           l1_24_port);
   U2_24 : ND3_30 port map( A => n27, B => A(24), C => Bn_24_port, Y => 
                           l2_24_port);
   U3_24 : ND3_29 port map( A => n31, B => A(24), C => B(24), Y => l3_24_port);
   U4_24 : ND4_8 port map( A => l0_24_port, B => l1_24_port, C => l2_24_port, D
                           => l3_24_port, Y => O(24));
   U0_25 : ND3_28 port map( A => n19, B => An_25_port, C => Bn_25_port, Y => 
                           l0_25_port);
   U1_25 : ND3_27 port map( A => n23, B => An_25_port, C => B(25), Y => 
                           l1_25_port);
   U2_25 : ND3_26 port map( A => n27, B => A(25), C => Bn_25_port, Y => 
                           l2_25_port);
   U3_25 : ND3_25 port map( A => n31, B => A(25), C => B(25), Y => l3_25_port);
   U4_25 : ND4_7 port map( A => l0_25_port, B => l1_25_port, C => l2_25_port, D
                           => l3_25_port, Y => O(25));
   U0_26 : ND3_24 port map( A => n19, B => An_26_port, C => Bn_26_port, Y => 
                           l0_26_port);
   U1_26 : ND3_23 port map( A => n23, B => An_26_port, C => B(26), Y => 
                           l1_26_port);
   U2_26 : ND3_22 port map( A => n27, B => A(26), C => Bn_26_port, Y => 
                           l2_26_port);
   U3_26 : ND3_21 port map( A => n31, B => A(26), C => B(26), Y => l3_26_port);
   U4_26 : ND4_6 port map( A => l0_26_port, B => l1_26_port, C => l2_26_port, D
                           => l3_26_port, Y => O(26));
   U0_27 : ND3_20 port map( A => n19, B => An_27_port, C => Bn_27_port, Y => 
                           l0_27_port);
   U1_27 : ND3_19 port map( A => n23, B => An_27_port, C => B(27), Y => 
                           l1_27_port);
   U2_27 : ND3_18 port map( A => n27, B => A(27), C => Bn_27_port, Y => 
                           l2_27_port);
   U3_27 : ND3_17 port map( A => n31, B => A(27), C => B(27), Y => l3_27_port);
   U4_27 : ND4_5 port map( A => l0_27_port, B => l1_27_port, C => l2_27_port, D
                           => l3_27_port, Y => O(27));
   U0_28 : ND3_16 port map( A => n19, B => An_28_port, C => Bn_28_port, Y => 
                           l0_28_port);
   U1_28 : ND3_15 port map( A => n23, B => An_28_port, C => B(28), Y => 
                           l1_28_port);
   U2_28 : ND3_14 port map( A => n27, B => A(28), C => Bn_28_port, Y => 
                           l2_28_port);
   U3_28 : ND3_13 port map( A => n31, B => A(28), C => B(28), Y => l3_28_port);
   U4_28 : ND4_4 port map( A => l0_28_port, B => l1_28_port, C => l2_28_port, D
                           => l3_28_port, Y => O(28));
   U0_29 : ND3_12 port map( A => n19, B => An_29_port, C => Bn_29_port, Y => 
                           l0_29_port);
   U1_29 : ND3_11 port map( A => n23, B => An_29_port, C => B(29), Y => 
                           l1_29_port);
   U2_29 : ND3_10 port map( A => n27, B => A(29), C => Bn_29_port, Y => 
                           l2_29_port);
   U3_29 : ND3_9 port map( A => n31, B => A(29), C => B(29), Y => l3_29_port);
   U4_29 : ND4_3 port map( A => l0_29_port, B => l1_29_port, C => l2_29_port, D
                           => l3_29_port, Y => O(29));
   U0_30 : ND3_8 port map( A => n19, B => An_30_port, C => Bn_30_port, Y => 
                           l0_30_port);
   U1_30 : ND3_7 port map( A => n23, B => An_30_port, C => B(30), Y => 
                           l1_30_port);
   U2_30 : ND3_6 port map( A => n27, B => A(30), C => Bn_30_port, Y => 
                           l2_30_port);
   U3_30 : ND3_5 port map( A => n31, B => A(30), C => B(30), Y => l3_30_port);
   U4_30 : ND4_2 port map( A => l0_30_port, B => l1_30_port, C => l2_30_port, D
                           => l3_30_port, Y => O(30));
   U0_31 : ND3_4 port map( A => n19, B => An_31_port, C => Bn_31_port, Y => 
                           l0_31_port);
   U1_31 : ND3_3 port map( A => n23, B => An_31_port, C => B(31), Y => 
                           l1_31_port);
   U2_31 : ND3_2 port map( A => n27, B => A(31), C => Bn_31_port, Y => 
                           l2_31_port);
   U3_31 : ND3_1 port map( A => n31, B => A(31), C => B(31), Y => l3_31_port);
   U4_31 : ND4_1 port map( A => l0_31_port, B => l1_31_port, C => l2_31_port, D
                           => l3_31_port, Y => O(31));
   U1 : BUF_X1 port map( A => S(0), Z => n20);
   U2 : BUF_X1 port map( A => S(1), Z => n24);
   U3 : BUF_X1 port map( A => S(2), Z => n28);
   U4 : BUF_X1 port map( A => S(3), Z => n32);
   U5 : BUF_X1 port map( A => n24, Z => n21);
   U6 : BUF_X1 port map( A => n28, Z => n25);
   U7 : BUF_X1 port map( A => n32, Z => n29);
   U8 : BUF_X1 port map( A => n20, Z => n17);
   U9 : BUF_X1 port map( A => n24, Z => n22);
   U10 : BUF_X1 port map( A => n28, Z => n26);
   U11 : BUF_X1 port map( A => n32, Z => n30);
   U12 : BUF_X1 port map( A => n20, Z => n18);
   U13 : BUF_X1 port map( A => n20, Z => n19);
   U14 : BUF_X1 port map( A => n24, Z => n23);
   U15 : BUF_X1 port map( A => n28, Z => n27);
   U16 : BUF_X1 port map( A => n32, Z => n31);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SHIFTER is

   port( data_in : in std_logic_vector (31 downto 0);  R : in std_logic_vector 
         (4 downto 0);  conf : in std_logic_vector (1 downto 0);  data_out : 
         out std_logic_vector (31 downto 0));

end SHIFTER;

architecture SYN_Behavioral of SHIFTER is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal mask_0_39_port, mask_0_38_port, mask_0_37_port, mask_0_36_port, 
      mask_0_35_port, mask_0_34_port, mask_0_33_port, mask_0_32_port, 
      mask_0_31_port, mask_0_30_port, mask_0_29_port, mask_0_28_port, 
      mask_0_27_port, mask_0_26_port, mask_0_25_port, mask_0_24_port, 
      mask_0_23_port, mask_0_22_port, mask_0_21_port, mask_0_20_port, 
      mask_0_19_port, mask_0_18_port, mask_0_17_port, mask_0_16_port, 
      mask_0_15_port, mask_0_14_port, mask_0_13_port, mask_0_12_port, 
      mask_0_11_port, mask_0_10_port, mask_0_9_port, mask_0_8_port, 
      mask_0_7_port, mask_0_6_port, mask_0_5_port, mask_0_4_port, mask_0_3_port
      , mask_0_2_port, mask_0_1_port, mask_0_0_port, mask_1_39_port, 
      mask_1_38_port, mask_1_37_port, mask_1_36_port, mask_1_35_port, 
      mask_1_34_port, mask_1_33_port, mask_1_32_port, mask_1_31_port, 
      mask_1_30_port, mask_1_29_port, mask_1_28_port, mask_1_27_port, 
      mask_1_26_port, mask_1_25_port, mask_1_24_port, mask_1_23_port, 
      mask_1_22_port, mask_1_21_port, mask_1_20_port, mask_1_19_port, 
      mask_1_18_port, mask_1_17_port, mask_1_16_port, mask_1_15_port, 
      mask_1_14_port, mask_1_13_port, mask_1_12_port, mask_1_11_port, 
      mask_1_10_port, mask_1_9_port, mask_1_8_port, mask_1_7_port, 
      mask_1_6_port, mask_1_5_port, mask_1_4_port, mask_1_3_port, mask_1_2_port
      , mask_1_1_port, mask_1_0_port, mask_2_39_port, mask_2_38_port, 
      mask_2_37_port, mask_2_36_port, mask_2_35_port, mask_2_34_port, 
      mask_2_33_port, mask_2_32_port, mask_2_31_port, mask_2_30_port, 
      mask_2_29_port, mask_2_28_port, mask_2_27_port, mask_2_26_port, 
      mask_2_25_port, mask_2_24_port, mask_2_23_port, mask_2_22_port, 
      mask_2_21_port, mask_2_20_port, mask_2_19_port, mask_2_18_port, 
      mask_2_17_port, mask_2_16_port, mask_2_15_port, mask_2_14_port, 
      mask_2_13_port, mask_2_12_port, mask_2_11_port, mask_2_10_port, 
      mask_2_9_port, mask_2_8_port, mask_2_7_port, mask_2_6_port, mask_2_5_port
      , mask_2_4_port, mask_2_3_port, mask_2_2_port, mask_2_1_port, 
      mask_2_0_port, mask_3_39_port, mask_3_38_port, mask_3_37_port, 
      mask_3_36_port, mask_3_35_port, mask_3_34_port, mask_3_33_port, 
      mask_3_32_port, mask_3_31_port, mask_3_30_port, mask_3_29_port, 
      mask_3_28_port, mask_3_27_port, mask_3_26_port, mask_3_25_port, 
      mask_3_24_port, mask_3_23_port, mask_3_22_port, mask_3_21_port, 
      mask_3_20_port, mask_3_19_port, mask_3_18_port, mask_3_17_port, 
      mask_3_16_port, mask_3_15_port, mask_3_14_port, mask_3_13_port, 
      mask_3_12_port, mask_3_11_port, mask_3_10_port, mask_3_9_port, 
      mask_3_8_port, mask_3_7_port, mask_3_6_port, mask_3_5_port, mask_3_4_port
      , mask_3_3_port, mask_3_2_port, mask_3_1_port, mask_3_0_port, N28, N35, 
      N37, N38, N39, N40, N41, N42, N43, N45, N46, N47, N48, N49, N50, N51, N53
      , N54, N55, N56, N57, N58, N59, N60, N68, N69, N70, N71, N72, N73, N74, 
      N75, N76, N77, N78, N79, N80, N81, N82, N83, N85, N86, N87, N88, N89, N90
      , N91, N92, N93, N94, N95, N96, N97, N98, N99, N108, N109, N110, N111, 
      N112, N113, N114, N115, N116, n9, n128, n129, n131, n132, n135, n137, 
      n138, n139, n140, n143, n144, n145, n146, n147, n148, n149, n151, n152, 
      n153, n154, n155, n156, n157, n159, n160, n161, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
      n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n629, n630, n631, 
      n632, n633, n634, n635, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
      n742 : std_logic;

begin
   
   mask_reg_0_39_inst : DLH_X1 port map( G => n619, D => n473, Q => 
                           mask_0_39_port);
   mask_reg_0_38_inst : DLH_X1 port map( G => n619, D => n482, Q => 
                           mask_0_38_port);
   mask_reg_0_37_inst : DLH_X1 port map( G => n619, D => n481, Q => 
                           mask_0_37_port);
   mask_reg_0_36_inst : DLH_X1 port map( G => n619, D => n480, Q => 
                           mask_0_36_port);
   mask_reg_0_35_inst : DLH_X1 port map( G => n619, D => n479, Q => 
                           mask_0_35_port);
   mask_reg_0_34_inst : DLH_X1 port map( G => n619, D => n478, Q => 
                           mask_0_34_port);
   mask_reg_0_33_inst : DLH_X1 port map( G => n618, D => n477, Q => 
                           mask_0_33_port);
   mask_reg_0_32_inst : DLH_X1 port map( G => n618, D => n476, Q => 
                           mask_0_32_port);
   mask_reg_0_31_inst : DLH_X1 port map( G => n618, D => N116, Q => 
                           mask_0_31_port);
   mask_reg_0_30_inst : DLH_X1 port map( G => n618, D => N115, Q => 
                           mask_0_30_port);
   mask_reg_0_29_inst : DLH_X1 port map( G => n618, D => N114, Q => 
                           mask_0_29_port);
   mask_reg_0_28_inst : DLH_X1 port map( G => n618, D => N113, Q => 
                           mask_0_28_port);
   mask_reg_0_27_inst : DLH_X1 port map( G => n618, D => N112, Q => 
                           mask_0_27_port);
   mask_reg_0_26_inst : DLH_X1 port map( G => n618, D => N111, Q => 
                           mask_0_26_port);
   mask_reg_0_25_inst : DLH_X1 port map( G => n618, D => N110, Q => 
                           mask_0_25_port);
   mask_reg_0_24_inst : DLH_X1 port map( G => n618, D => N109, Q => 
                           mask_0_24_port);
   mask_reg_0_23_inst : DLH_X1 port map( G => n618, D => N108, Q => 
                           mask_0_23_port);
   mask_reg_0_22_inst : DLH_X1 port map( G => n617, D => n484, Q => 
                           mask_0_22_port);
   mask_reg_0_21_inst : DLH_X1 port map( G => n617, D => n485, Q => 
                           mask_0_21_port);
   mask_reg_0_20_inst : DLH_X1 port map( G => n617, D => n486, Q => 
                           mask_0_20_port);
   mask_reg_0_19_inst : DLH_X1 port map( G => n617, D => n487, Q => 
                           mask_0_19_port);
   mask_reg_0_18_inst : DLH_X1 port map( G => n617, D => n488, Q => 
                           mask_0_18_port);
   mask_reg_0_17_inst : DLH_X1 port map( G => n617, D => n489, Q => 
                           mask_0_17_port);
   mask_reg_0_16_inst : DLH_X1 port map( G => n617, D => n490, Q => 
                           mask_0_16_port);
   mask_reg_0_15_inst : DLH_X1 port map( G => n617, D => n491, Q => 
                           mask_0_15_port);
   mask_reg_0_14_inst : DLH_X1 port map( G => n617, D => N99, Q => 
                           mask_0_14_port);
   mask_reg_0_13_inst : DLH_X1 port map( G => n617, D => N98, Q => 
                           mask_0_13_port);
   mask_reg_0_12_inst : DLH_X1 port map( G => n617, D => N97, Q => 
                           mask_0_12_port);
   mask_reg_0_11_inst : DLH_X1 port map( G => n616, D => N96, Q => 
                           mask_0_11_port);
   mask_reg_0_10_inst : DLH_X1 port map( G => n616, D => N95, Q => 
                           mask_0_10_port);
   mask_reg_0_9_inst : DLH_X1 port map( G => n616, D => N94, Q => mask_0_9_port
                           );
   mask_reg_0_8_inst : DLH_X1 port map( G => n616, D => N93, Q => mask_0_8_port
                           );
   mask_reg_0_7_inst : DLH_X1 port map( G => n616, D => N92, Q => mask_0_7_port
                           );
   mask_reg_0_6_inst : DLH_X1 port map( G => n616, D => N91, Q => mask_0_6_port
                           );
   mask_reg_0_5_inst : DLH_X1 port map( G => n616, D => N90, Q => mask_0_5_port
                           );
   mask_reg_0_4_inst : DLH_X1 port map( G => n616, D => N89, Q => mask_0_4_port
                           );
   mask_reg_0_3_inst : DLH_X1 port map( G => n616, D => N88, Q => mask_0_3_port
                           );
   mask_reg_0_2_inst : DLH_X1 port map( G => n616, D => N87, Q => mask_0_2_port
                           );
   mask_reg_0_1_inst : DLH_X1 port map( G => n616, D => N86, Q => mask_0_1_port
                           );
   mask_reg_0_0_inst : DLH_X1 port map( G => n615, D => N85, Q => mask_0_0_port
                           );
   mask_reg_1_39_inst : DLH_X1 port map( G => n615, D => n475, Q => 
                           mask_1_39_port);
   mask_reg_1_38_inst : DLH_X1 port map( G => n615, D => N83, Q => 
                           mask_1_38_port);
   mask_reg_1_37_inst : DLH_X1 port map( G => n615, D => N82, Q => 
                           mask_1_37_port);
   mask_reg_1_36_inst : DLH_X1 port map( G => n615, D => N81, Q => 
                           mask_1_36_port);
   mask_reg_1_35_inst : DLH_X1 port map( G => n615, D => N80, Q => 
                           mask_1_35_port);
   mask_reg_1_34_inst : DLH_X1 port map( G => n615, D => N79, Q => 
                           mask_1_34_port);
   mask_reg_1_33_inst : DLH_X1 port map( G => n615, D => N78, Q => 
                           mask_1_33_port);
   mask_reg_1_32_inst : DLH_X1 port map( G => n615, D => N77, Q => 
                           mask_1_32_port);
   mask_reg_1_31_inst : DLH_X1 port map( G => n615, D => N60, Q => 
                           mask_1_31_port);
   mask_reg_1_30_inst : DLH_X1 port map( G => n615, D => N59, Q => 
                           mask_1_30_port);
   mask_reg_1_29_inst : DLH_X1 port map( G => n614, D => N58, Q => 
                           mask_1_29_port);
   mask_reg_1_28_inst : DLH_X1 port map( G => n614, D => N57, Q => 
                           mask_1_28_port);
   mask_reg_1_27_inst : DLH_X1 port map( G => n614, D => N56, Q => 
                           mask_1_27_port);
   mask_reg_1_26_inst : DLH_X1 port map( G => n614, D => N55, Q => 
                           mask_1_26_port);
   mask_reg_1_25_inst : DLH_X1 port map( G => n614, D => N54, Q => 
                           mask_1_25_port);
   mask_reg_1_24_inst : DLH_X1 port map( G => n614, D => N53, Q => 
                           mask_1_24_port);
   mask_reg_1_23_inst : DLH_X1 port map( G => n614, D => N76, Q => 
                           mask_1_23_port);
   mask_reg_1_22_inst : DLH_X1 port map( G => n614, D => N75, Q => 
                           mask_1_22_port);
   mask_reg_1_21_inst : DLH_X1 port map( G => n614, D => N74, Q => 
                           mask_1_21_port);
   mask_reg_1_20_inst : DLH_X1 port map( G => n614, D => N73, Q => 
                           mask_1_20_port);
   mask_reg_1_19_inst : DLH_X1 port map( G => n614, D => N72, Q => 
                           mask_1_19_port);
   mask_reg_1_18_inst : DLH_X1 port map( G => n613, D => N71, Q => 
                           mask_1_18_port);
   mask_reg_1_17_inst : DLH_X1 port map( G => n613, D => N70, Q => 
                           mask_1_17_port);
   mask_reg_1_16_inst : DLH_X1 port map( G => n613, D => N69, Q => 
                           mask_1_16_port);
   mask_reg_1_15_inst : DLH_X1 port map( G => n613, D => n483, Q => 
                           mask_1_15_port);
   mask_reg_1_14_inst : DLH_X1 port map( G => n613, D => N51, Q => 
                           mask_1_14_port);
   mask_reg_1_13_inst : DLH_X1 port map( G => n613, D => N50, Q => 
                           mask_1_13_port);
   mask_reg_1_12_inst : DLH_X1 port map( G => n613, D => N49, Q => 
                           mask_1_12_port);
   mask_reg_1_11_inst : DLH_X1 port map( G => n613, D => N48, Q => 
                           mask_1_11_port);
   mask_reg_1_10_inst : DLH_X1 port map( G => n613, D => N47, Q => 
                           mask_1_10_port);
   mask_reg_1_9_inst : DLH_X1 port map( G => n613, D => N46, Q => mask_1_9_port
                           );
   mask_reg_1_8_inst : DLH_X1 port map( G => n613, D => N45, Q => mask_1_8_port
                           );
   mask_reg_1_7_inst : DLH_X1 port map( G => n612, D => N68, Q => mask_1_7_port
                           );
   mask_reg_1_6_inst : DLH_X1 port map( G => n612, D => n492, Q => 
                           mask_1_6_port);
   mask_reg_1_5_inst : DLH_X1 port map( G => n612, D => n493, Q => 
                           mask_1_5_port);
   mask_reg_1_4_inst : DLH_X1 port map( G => n612, D => n494, Q => 
                           mask_1_4_port);
   mask_reg_1_3_inst : DLH_X1 port map( G => n612, D => n495, Q => 
                           mask_1_3_port);
   mask_reg_1_2_inst : DLH_X1 port map( G => n612, D => n496, Q => 
                           mask_1_2_port);
   mask_reg_1_1_inst : DLH_X1 port map( G => n612, D => n497, Q => 
                           mask_1_1_port);
   mask_reg_1_0_inst : DLH_X1 port map( G => n612, D => n498, Q => 
                           mask_1_0_port);
   mask_reg_2_39_inst : DLH_X1 port map( G => n612, D => N60, Q => 
                           mask_2_39_port);
   mask_reg_2_38_inst : DLH_X1 port map( G => n612, D => N59, Q => 
                           mask_2_38_port);
   mask_reg_2_37_inst : DLH_X1 port map( G => n612, D => N58, Q => 
                           mask_2_37_port);
   mask_reg_2_36_inst : DLH_X1 port map( G => n611, D => N57, Q => 
                           mask_2_36_port);
   mask_reg_2_35_inst : DLH_X1 port map( G => n611, D => N56, Q => 
                           mask_2_35_port);
   mask_reg_2_34_inst : DLH_X1 port map( G => n611, D => N55, Q => 
                           mask_2_34_port);
   mask_reg_2_33_inst : DLH_X1 port map( G => n611, D => N54, Q => 
                           mask_2_33_port);
   mask_reg_2_32_inst : DLH_X1 port map( G => n611, D => N53, Q => 
                           mask_2_32_port);
   mask_reg_2_31_inst : DLH_X1 port map( G => n611, D => n474, Q => 
                           mask_2_31_port);
   mask_reg_2_30_inst : DLH_X1 port map( G => n611, D => N43, Q => 
                           mask_2_30_port);
   mask_reg_2_29_inst : DLH_X1 port map( G => n611, D => N42, Q => 
                           mask_2_29_port);
   mask_reg_2_28_inst : DLH_X1 port map( G => n611, D => N41, Q => 
                           mask_2_28_port);
   mask_reg_2_27_inst : DLH_X1 port map( G => n611, D => N40, Q => 
                           mask_2_27_port);
   mask_reg_2_26_inst : DLH_X1 port map( G => n611, D => N39, Q => 
                           mask_2_26_port);
   mask_reg_2_25_inst : DLH_X1 port map( G => n610, D => N38, Q => 
                           mask_2_25_port);
   mask_reg_2_24_inst : DLH_X1 port map( G => n610, D => N37, Q => 
                           mask_2_24_port);
   mask_reg_2_23_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_23_port);
   mask_reg_2_22_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_22_port);
   mask_reg_2_21_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_21_port);
   mask_reg_2_20_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_20_port);
   mask_reg_2_19_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_19_port);
   mask_reg_2_18_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_18_port);
   mask_reg_2_17_inst : DLH_X1 port map( G => n610, D => n536, Q => 
                           mask_2_17_port);
   mask_reg_2_16_inst : DLH_X1 port map( G => n610, D => n537, Q => 
                           mask_2_16_port);
   mask_reg_2_15_inst : DLH_X1 port map( G => n610, D => N35, Q => 
                           mask_2_15_port);
   mask_reg_2_14_inst : DLH_X1 port map( G => n609, D => n715, Q => 
                           mask_2_14_port);
   mask_reg_2_13_inst : DLH_X1 port map( G => n609, D => n714, Q => 
                           mask_2_13_port);
   mask_reg_2_12_inst : DLH_X1 port map( G => n609, D => n713, Q => 
                           mask_2_12_port);
   mask_reg_2_11_inst : DLH_X1 port map( G => n609, D => n712, Q => 
                           mask_2_11_port);
   mask_reg_2_10_inst : DLH_X1 port map( G => n609, D => n711, Q => 
                           mask_2_10_port);
   mask_reg_2_9_inst : DLH_X1 port map( G => n609, D => n710, Q => 
                           mask_2_9_port);
   mask_reg_2_8_inst : DLH_X1 port map( G => n609, D => n709, Q => 
                           mask_2_8_port);
   mask_reg_2_7_inst : DLH_X1 port map( G => n609, D => n483, Q => 
                           mask_2_7_port);
   mask_reg_2_6_inst : DLH_X1 port map( G => n609, D => N51, Q => mask_2_6_port
                           );
   mask_reg_2_5_inst : DLH_X1 port map( G => n609, D => N50, Q => mask_2_5_port
                           );
   mask_reg_2_4_inst : DLH_X1 port map( G => n609, D => N49, Q => mask_2_4_port
                           );
   mask_reg_2_3_inst : DLH_X1 port map( G => n608, D => N48, Q => mask_2_3_port
                           );
   mask_reg_2_2_inst : DLH_X1 port map( G => n608, D => N47, Q => mask_2_2_port
                           );
   mask_reg_2_1_inst : DLH_X1 port map( G => n608, D => N46, Q => mask_2_1_port
                           );
   mask_reg_2_0_inst : DLH_X1 port map( G => n608, D => N45, Q => mask_2_0_port
                           );
   mask_reg_3_39_inst : DLH_X1 port map( G => n608, D => n474, Q => 
                           mask_3_39_port);
   mask_reg_3_38_inst : DLH_X1 port map( G => n608, D => N43, Q => 
                           mask_3_38_port);
   mask_reg_3_37_inst : DLH_X1 port map( G => n608, D => N42, Q => 
                           mask_3_37_port);
   mask_reg_3_36_inst : DLH_X1 port map( G => n608, D => N41, Q => 
                           mask_3_36_port);
   mask_reg_3_35_inst : DLH_X1 port map( G => n608, D => N40, Q => 
                           mask_3_35_port);
   mask_reg_3_34_inst : DLH_X1 port map( G => n608, D => N39, Q => 
                           mask_3_34_port);
   mask_reg_3_33_inst : DLH_X1 port map( G => n608, D => N38, Q => 
                           mask_3_33_port);
   mask_reg_3_32_inst : DLH_X1 port map( G => n607, D => N37, Q => 
                           mask_3_32_port);
   mask_reg_3_31_inst : DLH_X1 port map( G => n607, D => n537, Q => 
                           mask_3_31_port);
   mask_reg_3_30_inst : DLH_X1 port map( G => n607, D => n537, Q => 
                           mask_3_30_port);
   mask_reg_3_29_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_29_port);
   mask_reg_3_28_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_28_port);
   mask_reg_3_27_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_27_port);
   mask_reg_3_26_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_26_port);
   mask_reg_3_25_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_25_port);
   mask_reg_3_24_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_24_port);
   mask_reg_3_23_inst : DLH_X1 port map( G => n607, D => n538, Q => 
                           mask_3_23_port);
   mask_reg_3_22_inst : DLH_X1 port map( G => n607, D => n536, Q => 
                           mask_3_22_port);
   mask_reg_3_21_inst : DLH_X1 port map( G => n606, D => n536, Q => 
                           mask_3_21_port);
   mask_reg_3_20_inst : DLH_X1 port map( G => n606, D => n536, Q => 
                           mask_3_20_port);
   mask_reg_3_19_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_19_port);
   mask_reg_3_18_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_18_port);
   mask_reg_3_17_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_17_port);
   mask_reg_3_16_inst : DLH_X1 port map( G => n606, D => n538, Q => 
                           mask_3_16_port);
   mask_reg_3_15_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_15_port);
   mask_reg_3_14_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_14_port);
   mask_reg_3_13_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_13_port);
   mask_reg_3_12_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_12_port);
   mask_reg_3_11_inst : DLH_X1 port map( G => n606, D => n537, Q => 
                           mask_3_11_port);
   mask_reg_3_10_inst : DLH_X1 port map( G => n605, D => n538, Q => 
                           mask_3_10_port);
   mask_reg_3_9_inst : DLH_X1 port map( G => n605, D => n538, Q => 
                           mask_3_9_port);
   mask_reg_3_8_inst : DLH_X1 port map( G => n605, D => n536, Q => 
                           mask_3_8_port);
   mask_reg_3_7_inst : DLH_X1 port map( G => n605, D => N35, Q => mask_3_7_port
                           );
   mask_reg_3_6_inst : DLH_X1 port map( G => n605, D => n715, Q => 
                           mask_3_6_port);
   mask_reg_3_5_inst : DLH_X1 port map( G => n605, D => n714, Q => 
                           mask_3_5_port);
   mask_reg_3_4_inst : DLH_X1 port map( G => n605, D => n713, Q => 
                           mask_3_4_port);
   mask_reg_3_3_inst : DLH_X1 port map( G => n605, D => n712, Q => 
                           mask_3_3_port);
   mask_reg_3_2_inst : DLH_X1 port map( G => n605, D => n711, Q => 
                           mask_3_2_port);
   mask_reg_3_1_inst : DLH_X1 port map( G => n605, D => n710, Q => 
                           mask_3_1_port);
   mask_reg_3_0_inst : DLH_X1 port map( G => n605, D => n709, Q => 
                           mask_3_0_port);
   U437 : AOI21_X2 port map( B1 => conf(1), B2 => conf(0), A => n398, ZN => 
                           n442);
   U564 : NAND3_X1 port map( A1 => data_in(31), A2 => n690, A3 => conf(0), ZN 
                           => n443);
   U3 : INV_X1 port map( A => n442, ZN => n708);
   U4 : BUF_X1 port map( A => n531, Z => n595);
   U5 : AND2_X1 port map( A1 => n398, A2 => n718, ZN => n526);
   U6 : AND2_X1 port map( A1 => R(4), A2 => n716, ZN => n527);
   U7 : OR2_X1 port map( A1 => n717, A2 => R(2), ZN => n528);
   U8 : OR2_X1 port map( A1 => R(1), A2 => R(2), ZN => n529);
   U9 : AND2_X1 port map( A1 => R(3), A2 => R(4), ZN => n530);
   U10 : BUF_X1 port map( A => n626, Z => n621);
   U11 : BUF_X1 port map( A => n626, Z => n620);
   U12 : BUF_X1 port map( A => n625, Z => n624);
   U13 : BUF_X1 port map( A => n625, Z => n623);
   U14 : BUF_X1 port map( A => n625, Z => n622);
   U15 : BUF_X1 port map( A => n528, Z => n584);
   U16 : BUF_X1 port map( A => n532, Z => n592);
   U17 : BUF_X1 port map( A => n533, Z => n588);
   U18 : BUF_X1 port map( A => n529, Z => n550);
   U19 : AND2_X1 port map( A1 => n544, A2 => n718, ZN => n531);
   U20 : BUF_X1 port map( A => n604, Z => n625);
   U21 : BUF_X1 port map( A => n532, Z => n591);
   U22 : BUF_X1 port map( A => n533, Z => n587);
   U23 : BUF_X1 port map( A => n528, Z => n583);
   U24 : BUF_X1 port map( A => n534, Z => n597);
   U25 : BUF_X1 port map( A => n529, Z => n549);
   U26 : BUF_X1 port map( A => n568, Z => n566);
   U27 : BUF_X1 port map( A => n561, Z => n559);
   U28 : BUF_X1 port map( A => n527, Z => n575);
   U29 : BUF_X1 port map( A => n530, Z => n569);
   U30 : AND2_X1 port map( A1 => R(2), A2 => n717, ZN => n532);
   U31 : BUF_X1 port map( A => n535, Z => n553);
   U32 : BUF_X1 port map( A => n691, Z => n539);
   U33 : BUF_X1 port map( A => n603, Z => n601);
   U34 : BUF_X1 port map( A => n603, Z => n602);
   U35 : BUF_X1 port map( A => n624, Z => n605);
   U36 : BUF_X1 port map( A => n624, Z => n606);
   U37 : BUF_X1 port map( A => n624, Z => n607);
   U38 : BUF_X1 port map( A => n623, Z => n608);
   U39 : BUF_X1 port map( A => n623, Z => n609);
   U40 : BUF_X1 port map( A => n623, Z => n610);
   U41 : BUF_X1 port map( A => n622, Z => n611);
   U42 : BUF_X1 port map( A => n622, Z => n612);
   U43 : BUF_X1 port map( A => n622, Z => n613);
   U44 : BUF_X1 port map( A => n621, Z => n614);
   U45 : BUF_X1 port map( A => n621, Z => n615);
   U46 : BUF_X1 port map( A => n621, Z => n616);
   U47 : BUF_X1 port map( A => n620, Z => n617);
   U48 : BUF_X1 port map( A => n620, Z => n618);
   U49 : BUF_X1 port map( A => n620, Z => n619);
   U50 : BUF_X1 port map( A => n575, Z => n577);
   U51 : BUF_X1 port map( A => n575, Z => n578);
   U52 : BUF_X1 port map( A => n566, Z => n563);
   U53 : BUF_X1 port map( A => n575, Z => n579);
   U54 : BUF_X1 port map( A => n566, Z => n564);
   U55 : BUF_X1 port map( A => n569, Z => n571);
   U56 : BUF_X1 port map( A => n569, Z => n572);
   U57 : BUF_X1 port map( A => n559, Z => n556);
   U58 : BUF_X1 port map( A => n569, Z => n573);
   U59 : BUF_X1 port map( A => n559, Z => n557);
   U60 : INV_X1 port map( A => n550, ZN => n547);
   U61 : INV_X1 port map( A => n550, ZN => n546);
   U62 : INV_X1 port map( A => n592, ZN => n589);
   U63 : INV_X1 port map( A => n588, ZN => n585);
   U64 : INV_X1 port map( A => n583, ZN => n582);
   U65 : INV_X1 port map( A => n549, ZN => n548);
   U66 : INV_X1 port map( A => n587, ZN => n586);
   U67 : INV_X1 port map( A => n591, ZN => n590);
   U68 : INV_X1 port map( A => n584, ZN => n581);
   U69 : INV_X1 port map( A => n595, ZN => n594);
   U70 : INV_X1 port map( A => n597, ZN => n596);
   U71 : BUF_X1 port map( A => n566, Z => n565);
   U72 : BUF_X1 port map( A => n559, Z => n558);
   U73 : OAI21_X1 port map( B1 => n541, B2 => n719, A => n600, ZN => n473);
   U74 : BUF_X1 port map( A => n604, Z => n626);
   U75 : BUF_X1 port map( A => n539, Z => n541);
   U76 : BUF_X1 port map( A => n539, Z => n543);
   U77 : BUF_X1 port map( A => n539, Z => n542);
   U78 : BUF_X1 port map( A => n567, Z => n562);
   U79 : BUF_X1 port map( A => n568, Z => n567);
   U80 : BUF_X1 port map( A => n560, Z => n555);
   U81 : BUF_X1 port map( A => n561, Z => n560);
   U82 : INV_X1 port map( A => n553, ZN => n552);
   U83 : INV_X1 port map( A => n553, ZN => n551);
   U84 : BUF_X1 port map( A => n534, Z => n598);
   U85 : BUF_X1 port map( A => n576, Z => n580);
   U86 : BUF_X1 port map( A => n527, Z => n576);
   U87 : BUF_X1 port map( A => n570, Z => n574);
   U88 : BUF_X1 port map( A => n530, Z => n570);
   U89 : BUF_X1 port map( A => n532, Z => n593);
   U90 : AOI221_X1 port map( B1 => n554, B2 => n680, C1 => n598, C2 => n376, A 
                           => n382, ZN => n381);
   U91 : OAI22_X1 port map( A1 => n374, A2 => n545, B1 => n383, B2 => n594, ZN 
                           => n382);
   U92 : AOI221_X1 port map( B1 => n554, B2 => n205, C1 => n598, C2 => n199, A 
                           => n206, ZN => n204);
   U93 : OAI22_X1 port map( A1 => n197, A2 => n545, B1 => n207, B2 => n594, ZN 
                           => n206);
   U94 : AOI221_X1 port map( B1 => n554, B2 => n160, C1 => n598, C2 => n152, A 
                           => n161, ZN => n159);
   U95 : OAI22_X1 port map( A1 => n149, A2 => n545, B1 => n163, B2 => n594, ZN 
                           => n161);
   U96 : NOR2_X1 port map( A1 => n708, A2 => n727, ZN => n483);
   U97 : NOR2_X1 port map( A1 => n734, A2 => n708, ZN => N45);
   U98 : NOR2_X1 port map( A1 => n733, A2 => n708, ZN => N46);
   U99 : NOR2_X1 port map( A1 => n732, A2 => n708, ZN => N47);
   U100 : NOR2_X1 port map( A1 => n731, A2 => n708, ZN => N48);
   U101 : NOR2_X1 port map( A1 => n730, A2 => n708, ZN => N49);
   U102 : NOR2_X1 port map( A1 => n729, A2 => n708, ZN => N50);
   U103 : NOR2_X1 port map( A1 => n728, A2 => n708, ZN => N51);
   U104 : AOI22_X1 port map( A1 => n680, A2 => n526, B1 => n684, B2 => n595, ZN
                           => n390);
   U105 : AOI22_X1 port map( A1 => n367, A2 => n526, B1 => n376, B2 => n595, ZN
                           => n375);
   U106 : AOI22_X1 port map( A1 => n367, A2 => n554, B1 => n359, B2 => n598, ZN
                           => n366);
   U107 : AOI22_X1 port map( A1 => n674, A2 => n526, B1 => n359, B2 => n595, ZN
                           => n358);
   U108 : INV_X1 port map( A => n349, ZN => n674);
   U109 : AOI22_X1 port map( A1 => n205, A2 => n526, B1 => n643, B2 => n595, ZN
                           => n215);
   U110 : INV_X1 port map( A => n216, ZN => n643);
   U111 : AOI22_X1 port map( A1 => n190, A2 => n526, B1 => n199, B2 => n595, ZN
                           => n198);
   U112 : AOI22_X1 port map( A1 => n190, A2 => n554, B1 => n182, B2 => n598, ZN
                           => n189);
   U113 : AOI22_X1 port map( A1 => n631, A2 => n526, B1 => n182, B2 => n595, ZN
                           => n181);
   U114 : INV_X1 port map( A => n172, ZN => n631);
   U115 : AOI22_X1 port map( A1 => n160, A2 => n526, B1 => n634, B2 => n595, ZN
                           => n173);
   U116 : INV_X1 port map( A => n174, ZN => n634);
   U117 : AOI22_X1 port map( A1 => n526, A2 => n132, B1 => n152, B2 => n595, ZN
                           => n151);
   U118 : OAI221_X1 port map( B1 => n552, B2 => n357, C1 => n596, C2 => n351, A
                           => n358, ZN => data_out(5));
   U119 : OAI221_X1 port map( B1 => n552, B2 => n349, C1 => n596, C2 => n343, A
                           => n672, ZN => data_out(6));
   U120 : OAI221_X1 port map( B1 => n552, B2 => n341, C1 => n596, C2 => n335, A
                           => n670, ZN => data_out(7));
   U121 : OAI221_X1 port map( B1 => n552, B2 => n325, C1 => n596, C2 => n319, A
                           => n666, ZN => data_out(9));
   U122 : OAI221_X1 port map( B1 => n552, B2 => n317, C1 => n596, C2 => n311, A
                           => n664, ZN => data_out(10));
   U123 : OAI221_X1 port map( B1 => n552, B2 => n309, C1 => n596, C2 => n303, A
                           => n662, ZN => data_out(11));
   U124 : OAI221_X1 port map( B1 => n552, B2 => n293, C1 => n596, C2 => n287, A
                           => n658, ZN => data_out(13));
   U125 : OAI221_X1 port map( B1 => n551, B2 => n285, C1 => n596, C2 => n279, A
                           => n656, ZN => data_out(14));
   U126 : OAI221_X1 port map( B1 => n551, B2 => n277, C1 => n596, C2 => n271, A
                           => n654, ZN => data_out(15));
   U127 : OAI221_X1 port map( B1 => n551, B2 => n261, C1 => n596, C2 => n255, A
                           => n650, ZN => data_out(17));
   U128 : OAI221_X1 port map( B1 => n551, B2 => n253, C1 => n596, C2 => n247, A
                           => n648, ZN => data_out(18));
   U129 : OAI221_X1 port map( B1 => n551, B2 => n245, C1 => n596, C2 => n239, A
                           => n646, ZN => data_out(19));
   U130 : OAI221_X1 port map( B1 => n552, B2 => n229, C1 => n596, C2 => n223, A
                           => n641, ZN => data_out(21));
   U131 : OAI221_X1 port map( B1 => n551, B2 => n221, C1 => n596, C2 => n216, A
                           => n639, ZN => data_out(22));
   U132 : OAI221_X1 port map( B1 => n551, B2 => n214, C1 => n596, C2 => n207, A
                           => n215, ZN => data_out(23));
   U133 : OAI221_X1 port map( B1 => n551, B2 => n197, C1 => n596, C2 => n188, A
                           => n198, ZN => data_out(25));
   U134 : OAI221_X1 port map( B1 => n545, B2 => n180, C1 => n594, C2 => n188, A
                           => n189, ZN => data_out(26));
   U135 : OAI221_X1 port map( B1 => n551, B2 => n180, C1 => n596, C2 => n174, A
                           => n181, ZN => data_out(27));
   U136 : INV_X1 port map( A => n159, ZN => data_out(29));
   U137 : OAI221_X1 port map( B1 => n149, B2 => n552, C1 => n596, C2 => n129, A
                           => n151, ZN => data_out(30));
   U138 : OAI222_X1 port map( A1 => n627, A2 => n596, B1 => n128, B2 => n544, 
                           C1 => n129, C2 => n594, ZN => data_out(31));
   U139 : NOR2_X1 port map( A1 => n742, A2 => n708, ZN => n498);
   U140 : NOR2_X1 port map( A1 => n741, A2 => n708, ZN => n497);
   U141 : NOR2_X1 port map( A1 => n740, A2 => n708, ZN => n496);
   U142 : NOR2_X1 port map( A1 => n739, A2 => n708, ZN => n495);
   U143 : NOR2_X1 port map( A1 => n738, A2 => n708, ZN => n494);
   U144 : NOR2_X1 port map( A1 => n737, A2 => n708, ZN => n493);
   U145 : NOR2_X1 port map( A1 => n736, A2 => n708, ZN => n492);
   U146 : NOR2_X1 port map( A1 => n735, A2 => n708, ZN => N68);
   U147 : INV_X1 port map( A => R(0), ZN => n718);
   U148 : OAI21_X1 port map( B1 => n543, B2 => n742, A => n600, ZN => N53);
   U149 : OAI21_X1 port map( B1 => n543, B2 => n741, A => n600, ZN => N54);
   U150 : OAI21_X1 port map( B1 => n543, B2 => n740, A => n600, ZN => N55);
   U151 : OAI21_X1 port map( B1 => n543, B2 => n739, A => n600, ZN => N56);
   U152 : OAI21_X1 port map( B1 => n543, B2 => n738, A => n600, ZN => N57);
   U153 : OAI21_X1 port map( B1 => n543, B2 => n737, A => n600, ZN => N58);
   U154 : OAI21_X1 port map( B1 => n543, B2 => n736, A => n600, ZN => N59);
   U155 : OAI21_X1 port map( B1 => n542, B2 => n735, A => n600, ZN => N60);
   U156 : AND2_X1 port map( A1 => R(2), A2 => R(1), ZN => n533);
   U157 : OAI21_X1 port map( B1 => n543, B2 => n734, A => n434, ZN => N109);
   U158 : OAI21_X1 port map( B1 => n544, B2 => n733, A => n433, ZN => N110);
   U159 : OAI21_X1 port map( B1 => n544, B2 => n732, A => n432, ZN => N111);
   U160 : OAI21_X1 port map( B1 => n543, B2 => n731, A => n431, ZN => N112);
   U161 : OAI21_X1 port map( B1 => n543, B2 => n730, A => n430, ZN => N113);
   U162 : OAI21_X1 port map( B1 => n543, B2 => n729, A => n429, ZN => N114);
   U163 : OAI21_X1 port map( B1 => n543, B2 => n728, A => n428, ZN => N115);
   U164 : AND2_X1 port map( A1 => R(0), A2 => n541, ZN => n534);
   U165 : OAI21_X1 port map( B1 => n542, B2 => n734, A => n600, ZN => N77);
   U166 : OAI21_X1 port map( B1 => n542, B2 => n733, A => n600, ZN => N78);
   U167 : OAI21_X1 port map( B1 => n542, B2 => n732, A => n600, ZN => N79);
   U168 : OAI21_X1 port map( B1 => n542, B2 => n731, A => n599, ZN => N80);
   U169 : OAI21_X1 port map( B1 => n542, B2 => n730, A => n599, ZN => N81);
   U170 : OAI21_X1 port map( B1 => n542, B2 => n729, A => n599, ZN => N82);
   U171 : OAI21_X1 port map( B1 => n542, B2 => n728, A => n599, ZN => N83);
   U172 : OAI21_X1 port map( B1 => n541, B2 => n727, A => n599, ZN => n475);
   U173 : OAI21_X1 port map( B1 => n542, B2 => n742, A => n706, ZN => n490);
   U174 : INV_X1 port map( A => N45, ZN => n706);
   U175 : OAI21_X1 port map( B1 => n542, B2 => n741, A => n705, ZN => n489);
   U176 : INV_X1 port map( A => N46, ZN => n705);
   U177 : OAI21_X1 port map( B1 => n542, B2 => n740, A => n704, ZN => n488);
   U178 : INV_X1 port map( A => N47, ZN => n704);
   U179 : OAI21_X1 port map( B1 => n542, B2 => n739, A => n703, ZN => n487);
   U180 : INV_X1 port map( A => N48, ZN => n703);
   U181 : OAI21_X1 port map( B1 => n541, B2 => n738, A => n702, ZN => n486);
   U182 : INV_X1 port map( A => N49, ZN => n702);
   U183 : OAI21_X1 port map( B1 => n541, B2 => n737, A => n701, ZN => n485);
   U184 : INV_X1 port map( A => N50, ZN => n701);
   U185 : OAI21_X1 port map( B1 => n541, B2 => n736, A => n700, ZN => n484);
   U186 : INV_X1 port map( A => N51, ZN => n700);
   U187 : OAI21_X1 port map( B1 => n541, B2 => n735, A => n707, ZN => N108);
   U188 : INV_X1 port map( A => n483, ZN => n707);
   U189 : OAI21_X1 port map( B1 => n543, B2 => n727, A => n689, ZN => N116);
   U190 : OAI21_X1 port map( B1 => n541, B2 => n726, A => n599, ZN => n476);
   U191 : INV_X1 port map( A => data_in(24), ZN => n726);
   U192 : OAI21_X1 port map( B1 => n541, B2 => n725, A => n599, ZN => n477);
   U193 : INV_X1 port map( A => data_in(25), ZN => n725);
   U194 : OAI21_X1 port map( B1 => n541, B2 => n724, A => n599, ZN => n478);
   U195 : INV_X1 port map( A => data_in(26), ZN => n724);
   U196 : OAI21_X1 port map( B1 => n541, B2 => n723, A => n599, ZN => n479);
   U197 : INV_X1 port map( A => data_in(27), ZN => n723);
   U198 : OAI21_X1 port map( B1 => n541, B2 => n722, A => n599, ZN => n480);
   U199 : INV_X1 port map( A => data_in(28), ZN => n722);
   U200 : OAI21_X1 port map( B1 => n542, B2 => n721, A => n599, ZN => n481);
   U201 : INV_X1 port map( A => data_in(29), ZN => n721);
   U202 : OAI21_X1 port map( B1 => n541, B2 => n720, A => n599, ZN => n482);
   U203 : INV_X1 port map( A => data_in(30), ZN => n720);
   U204 : NAND2_X1 port map( A1 => n434, A2 => n441, ZN => N69);
   U205 : NAND2_X1 port map( A1 => n433, A2 => n440, ZN => N70);
   U206 : NAND2_X1 port map( A1 => n432, A2 => n439, ZN => N71);
   U207 : NAND2_X1 port map( A1 => n431, A2 => n438, ZN => N72);
   U208 : NAND2_X1 port map( A1 => n430, A2 => n437, ZN => N73);
   U209 : NAND2_X1 port map( A1 => n429, A2 => n436, ZN => N74);
   U210 : NAND2_X1 port map( A1 => n428, A2 => n435, ZN => N75);
   U211 : INV_X1 port map( A => R(1), ZN => n717);
   U212 : INV_X1 port map( A => n434, ZN => n709);
   U213 : INV_X1 port map( A => n433, ZN => n710);
   U214 : INV_X1 port map( A => n432, ZN => n711);
   U215 : INV_X1 port map( A => n431, ZN => n712);
   U216 : INV_X1 port map( A => n430, ZN => n713);
   U217 : INV_X1 port map( A => n429, ZN => n714);
   U218 : INV_X1 port map( A => n428, ZN => n715);
   U219 : INV_X1 port map( A => data_in(31), ZN => n719);
   U220 : NAND2_X1 port map( A1 => n599, A2 => n441, ZN => N37);
   U221 : NAND2_X1 port map( A1 => n600, A2 => n440, ZN => N38);
   U222 : NAND2_X1 port map( A1 => n599, A2 => n439, ZN => N39);
   U223 : NAND2_X1 port map( A1 => n600, A2 => n438, ZN => N40);
   U224 : NAND2_X1 port map( A1 => n599, A2 => n437, ZN => N41);
   U225 : NAND2_X1 port map( A1 => n600, A2 => n436, ZN => N42);
   U226 : NAND2_X1 port map( A1 => n599, A2 => n435, ZN => N43);
   U227 : NAND2_X1 port map( A1 => n600, A2 => n427, ZN => n474);
   U228 : INV_X1 port map( A => R(3), ZN => n716);
   U229 : BUF_X1 port map( A => n143, Z => n568);
   U230 : NOR2_X1 port map( A1 => R(3), A2 => R(4), ZN => n143);
   U231 : BUF_X1 port map( A => n144, Z => n561);
   U232 : NOR2_X1 port map( A1 => n716, A2 => R(4), ZN => n144);
   U233 : NAND2_X1 port map( A1 => n698, A2 => n441, ZN => N93);
   U234 : INV_X1 port map( A => n498, ZN => n698);
   U235 : NAND2_X1 port map( A1 => n697, A2 => n440, ZN => N94);
   U236 : INV_X1 port map( A => n497, ZN => n697);
   U237 : NAND2_X1 port map( A1 => n696, A2 => n439, ZN => N95);
   U238 : INV_X1 port map( A => n496, ZN => n696);
   U239 : NAND2_X1 port map( A1 => n695, A2 => n438, ZN => N96);
   U240 : INV_X1 port map( A => n495, ZN => n695);
   U241 : NAND2_X1 port map( A1 => n694, A2 => n437, ZN => N97);
   U242 : INV_X1 port map( A => n494, ZN => n694);
   U243 : NAND2_X1 port map( A1 => n693, A2 => n436, ZN => N98);
   U244 : INV_X1 port map( A => n493, ZN => n693);
   U245 : NAND2_X1 port map( A1 => n692, A2 => n435, ZN => N99);
   U246 : INV_X1 port map( A => n492, ZN => n692);
   U247 : NAND2_X1 port map( A1 => n699, A2 => n427, ZN => n491);
   U248 : INV_X1 port map( A => N68, ZN => n699);
   U249 : INV_X1 port map( A => n270, ZN => n652);
   U250 : OAI22_X1 port map( A1 => n261, A2 => n545, B1 => n271, B2 => n594, ZN
                           => n270);
   U251 : INV_X1 port map( A => n350, ZN => n672);
   U252 : OAI22_X1 port map( A1 => n341, A2 => n545, B1 => n351, B2 => n594, ZN
                           => n350);
   U253 : INV_X1 port map( A => n342, ZN => n670);
   U254 : OAI22_X1 port map( A1 => n333, A2 => n545, B1 => n343, B2 => n594, ZN
                           => n342);
   U255 : INV_X1 port map( A => n334, ZN => n668);
   U256 : OAI22_X1 port map( A1 => n325, A2 => n545, B1 => n335, B2 => n594, ZN
                           => n334);
   U257 : INV_X1 port map( A => n326, ZN => n666);
   U258 : OAI22_X1 port map( A1 => n317, A2 => n545, B1 => n327, B2 => n594, ZN
                           => n326);
   U259 : INV_X1 port map( A => n318, ZN => n664);
   U260 : OAI22_X1 port map( A1 => n309, A2 => n545, B1 => n319, B2 => n594, ZN
                           => n318);
   U261 : INV_X1 port map( A => n310, ZN => n662);
   U262 : OAI22_X1 port map( A1 => n301, A2 => n545, B1 => n311, B2 => n594, ZN
                           => n310);
   U263 : INV_X1 port map( A => n302, ZN => n660);
   U264 : OAI22_X1 port map( A1 => n293, A2 => n545, B1 => n303, B2 => n594, ZN
                           => n302);
   U265 : INV_X1 port map( A => n294, ZN => n658);
   U266 : OAI22_X1 port map( A1 => n285, A2 => n545, B1 => n295, B2 => n594, ZN
                           => n294);
   U267 : INV_X1 port map( A => n286, ZN => n656);
   U268 : OAI22_X1 port map( A1 => n277, A2 => n545, B1 => n287, B2 => n594, ZN
                           => n286);
   U269 : INV_X1 port map( A => n278, ZN => n654);
   U270 : OAI22_X1 port map( A1 => n269, A2 => n545, B1 => n279, B2 => n594, ZN
                           => n278);
   U271 : INV_X1 port map( A => n262, ZN => n650);
   U272 : OAI22_X1 port map( A1 => n253, A2 => n545, B1 => n263, B2 => n594, ZN
                           => n262);
   U273 : INV_X1 port map( A => n254, ZN => n648);
   U274 : OAI22_X1 port map( A1 => n245, A2 => n545, B1 => n255, B2 => n594, ZN
                           => n254);
   U275 : INV_X1 port map( A => n246, ZN => n646);
   U276 : OAI22_X1 port map( A1 => n237, A2 => n545, B1 => n247, B2 => n594, ZN
                           => n246);
   U277 : INV_X1 port map( A => n238, ZN => n644);
   U278 : OAI22_X1 port map( A1 => n229, A2 => n545, B1 => n239, B2 => n594, ZN
                           => n238);
   U279 : INV_X1 port map( A => n230, ZN => n641);
   U280 : OAI22_X1 port map( A1 => n221, A2 => n545, B1 => n231, B2 => n594, ZN
                           => n230);
   U281 : INV_X1 port map( A => n222, ZN => n639);
   U282 : OAI22_X1 port map( A1 => n214, A2 => n545, B1 => n223, B2 => n594, ZN
                           => n222);
   U283 : NAND2_X1 port map( A1 => n427, A2 => n689, ZN => N76);
   U284 : BUF_X1 port map( A => N28, Z => n604);
   U285 : NAND2_X1 port map( A1 => n544, A2 => n708, ZN => N28);
   U286 : INV_X1 port map( A => n526, ZN => n545);
   U287 : INV_X1 port map( A => n601, ZN => n599);
   U288 : INV_X1 port map( A => n601, ZN => n600);
   U289 : BUF_X1 port map( A => n535, Z => n554);
   U290 : BUF_X1 port map( A => n540, Z => n544);
   U291 : BUF_X1 port map( A => n691, Z => n540);
   U292 : BUF_X1 port map( A => n602, Z => n537);
   U293 : BUF_X1 port map( A => n602, Z => n536);
   U294 : BUF_X1 port map( A => n602, Z => n538);
   U295 : AOI221_X1 port map( B1 => n592, B2 => n633, C1 => n588, C2 => n637, A
                           => n153, ZN => n132);
   U296 : OAI22_X1 port map( A1 => n148, A2 => n550, B1 => n147, B2 => n584, ZN
                           => n153);
   U297 : AOI221_X1 port map( B1 => n588, B2 => n681, C1 => n581, C2 => n686, A
                           => n387, ZN => n376);
   U298 : OAI22_X1 port map( A1 => n388, A2 => n550, B1 => n360, B2 => n590, ZN
                           => n387);
   U299 : AOI221_X1 port map( B1 => n588, B2 => n638, C1 => n592, C2 => n642, A
                           => n212, ZN => n199);
   U300 : OAI22_X1 port map( A1 => n192, A2 => n584, B1 => n213, B2 => n550, ZN
                           => n212);
   U301 : AOI221_X1 port map( B1 => n588, B2 => n630, C1 => n593, C2 => n633, A
                           => n169, ZN => n152);
   U302 : INV_X1 port map( A => n147, ZN => n630);
   U303 : OAI22_X1 port map( A1 => n170, A2 => n584, B1 => n171, B2 => n550, ZN
                           => n169);
   U304 : AOI221_X1 port map( B1 => n588, B2 => n686, C1 => n592, C2 => n683, A
                           => n377, ZN => n367);
   U305 : OAI22_X1 port map( A1 => n328, A2 => n550, B1 => n344, B2 => n584, ZN
                           => n377);
   U306 : AOI221_X1 port map( B1 => n592, B2 => n642, C1 => n588, C2 => n647, A
                           => n200, ZN => n190);
   U307 : OAI22_X1 port map( A1 => n164, A2 => n550, B1 => n165, B2 => n584, ZN
                           => n200);
   U308 : AOI221_X1 port map( B1 => n592, B2 => n647, C1 => n533, C2 => n651, A
                           => n217, ZN => n205);
   U309 : OAI22_X1 port map( A1 => n165, A2 => n550, B1 => n183, B2 => n584, ZN
                           => n217);
   U310 : AOI221_X1 port map( B1 => n592, B2 => n637, C1 => n588, C2 => n640, A
                           => n175, ZN => n160);
   U311 : OAI22_X1 port map( A1 => n147, A2 => n550, B1 => n176, B2 => n584, ZN
                           => n175);
   U312 : AOI221_X1 port map( B1 => n588, B2 => n677, C1 => n592, C2 => n681, A
                           => n368, ZN => n359);
   U313 : OAI22_X1 port map( A1 => n369, A2 => n550, B1 => n360, B2 => n584, ZN
                           => n368);
   U314 : AOI221_X1 port map( B1 => n588, B2 => n635, C1 => n592, C2 => n638, A
                           => n191, ZN => n182);
   U315 : OAI22_X1 port map( A1 => n183, A2 => n584, B1 => n192, B2 => n550, ZN
                           => n191);
   U316 : OAI221_X1 port map( B1 => n590, B2 => n164, C1 => n586, C2 => n165, A
                           => n166, ZN => n149);
   U317 : AOI22_X1 port map( A1 => n629, A2 => n546, B1 => n632, B2 => n582, ZN
                           => n166);
   U318 : INV_X1 port map( A => n137, ZN => n629);
   U319 : OAI221_X1 port map( B1 => n585, B2 => n137, C1 => n590, C2 => n156, A
                           => n157, ZN => n129);
   U320 : AOI22_X1 port map( A1 => n635, A2 => n581, B1 => n638, B2 => n548, ZN
                           => n157);
   U321 : OAI221_X1 port map( B1 => n585, B2 => n183, C1 => n589, C2 => n192, A
                           => n228, ZN => n216);
   U322 : AOI22_X1 port map( A1 => n651, A2 => n582, B1 => n655, B2 => n546, ZN
                           => n228);
   U323 : OAI221_X1 port map( B1 => n586, B2 => n176, C1 => n590, C2 => n170, A
                           => n187, ZN => n174);
   U324 : AOI22_X1 port map( A1 => n640, A2 => n581, B1 => n645, B2 => n547, ZN
                           => n187);
   U325 : OAI221_X1 port map( B1 => n589, B2 => n352, C1 => n584, C2 => n370, A
                           => n380, ZN => n365);
   U326 : AOI22_X1 port map( A1 => n679, A2 => n588, B1 => n687, B2 => n546, ZN
                           => n380);
   U327 : OAI221_X1 port map( B1 => n585, B2 => n170, C1 => n589, C2 => n171, A
                           => n203, ZN => n188);
   U328 : AOI22_X1 port map( A1 => n645, A2 => n581, B1 => n649, B2 => n548, ZN
                           => n203);
   U329 : OAI221_X1 port map( B1 => n590, B2 => n165, C1 => n586, C2 => n183, A
                           => n184, ZN => n172);
   U330 : AOI22_X1 port map( A1 => n632, A2 => n546, B1 => n635, B2 => n582, ZN
                           => n184);
   U331 : OAI221_X1 port map( B1 => n589, B2 => n344, C1 => n585, C2 => n360, A
                           => n361, ZN => n349);
   U332 : AOI22_X1 port map( A1 => n675, A2 => n546, B1 => n677, B2 => n582, ZN
                           => n361);
   U333 : OAI221_X1 port map( B1 => n585, B2 => n232, C1 => n590, C2 => n248, A
                           => n276, ZN => n263);
   U334 : AOI22_X1 port map( A1 => n663, A2 => n581, B1 => n667, B2 => n548, ZN
                           => n276);
   U335 : OAI221_X1 port map( B1 => n585, B2 => n320, C1 => n590, C2 => n336, A
                           => n364, ZN => n351);
   U336 : AOI22_X1 port map( A1 => n682, A2 => n581, B1 => n685, B2 => n548, ZN
                           => n364);
   U337 : OAI221_X1 port map( B1 => n586, B2 => n312, C1 => n589, C2 => n328, A
                           => n356, ZN => n343);
   U338 : AOI22_X1 port map( A1 => n681, A2 => n581, B1 => n683, B2 => n548, ZN
                           => n356);
   U339 : OAI221_X1 port map( B1 => n585, B2 => n304, C1 => n590, C2 => n320, A
                           => n348, ZN => n335);
   U340 : AOI22_X1 port map( A1 => n679, A2 => n581, B1 => n682, B2 => n548, ZN
                           => n348);
   U341 : OAI221_X1 port map( B1 => n586, B2 => n296, C1 => n589, C2 => n312, A
                           => n340, ZN => n327);
   U342 : AOI22_X1 port map( A1 => n677, A2 => n581, B1 => n681, B2 => n548, ZN
                           => n340);
   U343 : OAI221_X1 port map( B1 => n585, B2 => n288, C1 => n590, C2 => n304, A
                           => n332, ZN => n319);
   U344 : AOI22_X1 port map( A1 => n676, A2 => n581, B1 => n679, B2 => n548, ZN
                           => n332);
   U345 : OAI221_X1 port map( B1 => n586, B2 => n280, C1 => n589, C2 => n296, A
                           => n324, ZN => n311);
   U346 : AOI22_X1 port map( A1 => n675, A2 => n582, B1 => n677, B2 => n548, ZN
                           => n324);
   U347 : OAI221_X1 port map( B1 => n585, B2 => n272, C1 => n590, C2 => n288, A
                           => n316, ZN => n303);
   U348 : AOI22_X1 port map( A1 => n673, A2 => n581, B1 => n676, B2 => n548, ZN
                           => n316);
   U349 : OAI221_X1 port map( B1 => n585, B2 => n264, C1 => n590, C2 => n280, A
                           => n308, ZN => n295);
   U350 : AOI22_X1 port map( A1 => n671, A2 => n582, B1 => n675, B2 => n548, ZN
                           => n308);
   U351 : OAI221_X1 port map( B1 => n585, B2 => n256, C1 => n590, C2 => n272, A
                           => n300, ZN => n287);
   U352 : AOI22_X1 port map( A1 => n669, A2 => n582, B1 => n673, B2 => n548, ZN
                           => n300);
   U353 : OAI221_X1 port map( B1 => n585, B2 => n248, C1 => n590, C2 => n264, A
                           => n292, ZN => n279);
   U354 : AOI22_X1 port map( A1 => n667, A2 => n582, B1 => n671, B2 => n548, ZN
                           => n292);
   U355 : OAI221_X1 port map( B1 => n585, B2 => n240, C1 => n590, C2 => n256, A
                           => n284, ZN => n271);
   U356 : AOI22_X1 port map( A1 => n665, A2 => n582, B1 => n669, B2 => n548, ZN
                           => n284);
   U357 : OAI221_X1 port map( B1 => n585, B2 => n224, C1 => n590, C2 => n240, A
                           => n268, ZN => n255);
   U358 : AOI22_X1 port map( A1 => n661, A2 => n582, B1 => n665, B2 => n546, ZN
                           => n268);
   U359 : OAI221_X1 port map( B1 => n585, B2 => n213, C1 => n590, C2 => n232, A
                           => n260, ZN => n247);
   U360 : AOI22_X1 port map( A1 => n659, A2 => n582, B1 => n663, B2 => n547, ZN
                           => n260);
   U361 : OAI221_X1 port map( B1 => n585, B2 => n208, C1 => n590, C2 => n224, A
                           => n252, ZN => n239);
   U362 : AOI22_X1 port map( A1 => n657, A2 => n582, B1 => n661, B2 => n548, ZN
                           => n252);
   U363 : OAI221_X1 port map( B1 => n586, B2 => n192, C1 => n590, C2 => n213, A
                           => n244, ZN => n231);
   U364 : AOI22_X1 port map( A1 => n655, A2 => n582, B1 => n659, B2 => n546, ZN
                           => n244);
   U365 : OAI221_X1 port map( B1 => n585, B2 => n193, C1 => n590, C2 => n208, A
                           => n236, ZN => n223);
   U366 : AOI22_X1 port map( A1 => n653, A2 => n582, B1 => n657, B2 => n547, ZN
                           => n236);
   U367 : OAI221_X1 port map( B1 => n585, B2 => n171, C1 => n589, C2 => n193, A
                           => n220, ZN => n207);
   U368 : AOI22_X1 port map( A1 => n649, A2 => n581, B1 => n653, B2 => n548, ZN
                           => n220);
   U369 : OAI221_X1 port map( B1 => n584, B2 => n395, C1 => n589, C2 => n370, A
                           => n396, ZN => n383);
   U370 : AOI22_X1 port map( A1 => n682, A2 => n588, B1 => n688, B2 => n547, ZN
                           => n396);
   U371 : OAI221_X1 port map( B1 => n586, B2 => n156, C1 => n590, C2 => n164, A
                           => n179, ZN => n163);
   U372 : AOI22_X1 port map( A1 => n638, A2 => n581, B1 => n642, B2 => n546, ZN
                           => n179);
   U373 : OAI221_X1 port map( B1 => n590, B2 => n370, C1 => n584, C2 => n352, A
                           => n384, ZN => n374);
   U374 : AOI22_X1 port map( A1 => n679, A2 => n546, B1 => n687, B2 => n588, ZN
                           => n384);
   U375 : OAI221_X1 port map( B1 => n589, B2 => n264, C1 => n586, C2 => n280, A
                           => n281, ZN => n269);
   U376 : AOI22_X1 port map( A1 => n655, A2 => n547, B1 => n659, B2 => n582, ZN
                           => n281);
   U377 : OAI221_X1 port map( B1 => n589, B2 => n328, C1 => n585, C2 => n344, A
                           => n345, ZN => n333);
   U378 : AOI22_X1 port map( A1 => n671, A2 => n546, B1 => n675, B2 => n581, ZN
                           => n345);
   U379 : OAI221_X1 port map( B1 => n589, B2 => n320, C1 => n585, C2 => n336, A
                           => n337, ZN => n325);
   U380 : AOI22_X1 port map( A1 => n669, A2 => n546, B1 => n673, B2 => n582, ZN
                           => n337);
   U381 : OAI221_X1 port map( B1 => n589, B2 => n312, C1 => n586, C2 => n328, A
                           => n329, ZN => n317);
   U382 : AOI22_X1 port map( A1 => n667, A2 => n547, B1 => n671, B2 => n581, ZN
                           => n329);
   U383 : OAI221_X1 port map( B1 => n589, B2 => n304, C1 => n585, C2 => n320, A
                           => n321, ZN => n309);
   U384 : AOI22_X1 port map( A1 => n665, A2 => n547, B1 => n669, B2 => n582, ZN
                           => n321);
   U385 : OAI221_X1 port map( B1 => n589, B2 => n296, C1 => n586, C2 => n312, A
                           => n313, ZN => n301);
   U386 : AOI22_X1 port map( A1 => n663, A2 => n547, B1 => n667, B2 => n581, ZN
                           => n313);
   U387 : OAI221_X1 port map( B1 => n589, B2 => n288, C1 => n586, C2 => n304, A
                           => n305, ZN => n293);
   U388 : AOI22_X1 port map( A1 => n661, A2 => n547, B1 => n665, B2 => n581, ZN
                           => n305);
   U389 : OAI221_X1 port map( B1 => n589, B2 => n280, C1 => n585, C2 => n296, A
                           => n297, ZN => n285);
   U390 : AOI22_X1 port map( A1 => n659, A2 => n547, B1 => n663, B2 => n582, ZN
                           => n297);
   U391 : OAI221_X1 port map( B1 => n589, B2 => n272, C1 => n585, C2 => n288, A
                           => n289, ZN => n277);
   U392 : AOI22_X1 port map( A1 => n657, A2 => n547, B1 => n661, B2 => n581, ZN
                           => n289);
   U393 : OAI221_X1 port map( B1 => n590, B2 => n256, C1 => n586, C2 => n272, A
                           => n273, ZN => n261);
   U394 : AOI22_X1 port map( A1 => n653, A2 => n547, B1 => n657, B2 => n581, ZN
                           => n273);
   U395 : OAI221_X1 port map( B1 => n589, B2 => n248, C1 => n585, C2 => n264, A
                           => n265, ZN => n253);
   U396 : AOI22_X1 port map( A1 => n651, A2 => n547, B1 => n655, B2 => n582, ZN
                           => n265);
   U397 : OAI221_X1 port map( B1 => n590, B2 => n240, C1 => n586, C2 => n256, A
                           => n257, ZN => n245);
   U398 : AOI22_X1 port map( A1 => n649, A2 => n547, B1 => n653, B2 => n581, ZN
                           => n257);
   U399 : OAI221_X1 port map( B1 => n590, B2 => n232, C1 => n586, C2 => n248, A
                           => n249, ZN => n237);
   U400 : AOI22_X1 port map( A1 => n647, A2 => n547, B1 => n651, B2 => n582, ZN
                           => n249);
   U401 : OAI221_X1 port map( B1 => n589, B2 => n224, C1 => n586, C2 => n240, A
                           => n241, ZN => n229);
   U402 : AOI22_X1 port map( A1 => n645, A2 => n547, B1 => n649, B2 => n582, ZN
                           => n241);
   U403 : OAI221_X1 port map( B1 => n589, B2 => n208, C1 => n586, C2 => n224, A
                           => n225, ZN => n214);
   U404 : AOI22_X1 port map( A1 => n640, A2 => n547, B1 => n645, B2 => n581, ZN
                           => n225);
   U405 : OAI221_X1 port map( B1 => n590, B2 => n193, C1 => n586, C2 => n208, A
                           => n209, ZN => n197);
   U406 : AOI22_X1 port map( A1 => n637, A2 => n546, B1 => n640, B2 => n581, ZN
                           => n209);
   U407 : OAI221_X1 port map( B1 => n589, B2 => n336, C1 => n586, C2 => n352, A
                           => n353, ZN => n341);
   U408 : AOI22_X1 port map( A1 => n673, A2 => n546, B1 => n676, B2 => n582, ZN
                           => n353);
   U409 : OAI221_X1 port map( B1 => n589, B2 => n213, C1 => n586, C2 => n232, A
                           => n233, ZN => n221);
   U410 : AOI22_X1 port map( A1 => n642, A2 => n546, B1 => n647, B2 => n582, ZN
                           => n233);
   U411 : OAI221_X1 port map( B1 => n589, B2 => n352, C1 => n585, C2 => n370, A
                           => n371, ZN => n357);
   U412 : AOI22_X1 port map( A1 => n676, A2 => n546, B1 => n679, B2 => n581, ZN
                           => n371);
   U413 : OAI221_X1 port map( B1 => n589, B2 => n171, C1 => n586, C2 => n193, A
                           => n194, ZN => n180);
   U414 : AOI22_X1 port map( A1 => n633, A2 => n546, B1 => n637, B2 => n581, ZN
                           => n194);
   U415 : OAI221_X1 port map( B1 => n585, B2 => n400, C1 => n584, C2 => n370, A
                           => n401, ZN => n389);
   U416 : AOI22_X1 port map( A1 => n687, A2 => n592, B1 => n682, B2 => n546, ZN
                           => n401);
   U417 : AOI221_X1 port map( B1 => n592, B2 => n388, C1 => n548, C2 => n360, A
                           => n418, ZN => n397);
   U418 : OAI22_X1 port map( A1 => n407, A2 => n586, B1 => n686, B2 => n584, ZN
                           => n418);
   U419 : NAND2_X1 port map( A1 => n442, A2 => data_in(24), ZN => n434);
   U420 : NAND2_X1 port map( A1 => n442, A2 => data_in(25), ZN => n433);
   U421 : NAND2_X1 port map( A1 => n442, A2 => data_in(26), ZN => n432);
   U422 : NAND2_X1 port map( A1 => n442, A2 => data_in(27), ZN => n431);
   U423 : NAND2_X1 port map( A1 => n442, A2 => data_in(28), ZN => n430);
   U424 : NAND2_X1 port map( A1 => n442, A2 => data_in(29), ZN => n429);
   U425 : NAND2_X1 port map( A1 => n442, A2 => data_in(30), ZN => n428);
   U426 : OAI221_X1 port map( B1 => n551, B2 => n269, C1 => n596, C2 => n263, A
                           => n652, ZN => data_out(16));
   U427 : OAI222_X1 port map( A1 => n397, A2 => n551, B1 => n398, B2 => n399, 
                           C1 => n545, C2 => n389, ZN => data_out(0));
   U428 : OAI221_X1 port map( B1 => n552, B2 => n389, C1 => n596, C2 => n383, A
                           => n390, ZN => data_out(1));
   U429 : INV_X1 port map( A => n381, ZN => data_out(2));
   U430 : OAI221_X1 port map( B1 => n552, B2 => n374, C1 => n596, C2 => n365, A
                           => n375, ZN => data_out(3));
   U431 : OAI221_X1 port map( B1 => n545, B2 => n357, C1 => n594, C2 => n365, A
                           => n366, ZN => data_out(4));
   U432 : OAI221_X1 port map( B1 => n552, B2 => n333, C1 => n596, C2 => n327, A
                           => n668, ZN => data_out(8));
   U433 : OAI221_X1 port map( B1 => n552, B2 => n301, C1 => n596, C2 => n295, A
                           => n660, ZN => data_out(12));
   U434 : OAI221_X1 port map( B1 => n551, B2 => n237, C1 => n596, C2 => n231, A
                           => n644, ZN => data_out(20));
   U435 : INV_X1 port map( A => n204, ZN => data_out(24));
   U436 : OAI221_X1 port map( B1 => n551, B2 => n172, C1 => n596, C2 => n163, A
                           => n173, ZN => data_out(28));
   U438 : AOI22_X1 port map( A1 => n131, A2 => n718, B1 => R(0), B2 => n132, ZN
                           => n128);
   U439 : OAI221_X1 port map( B1 => n632, B2 => n590, C1 => n635, C2 => n586, A
                           => n135, ZN => n131);
   U440 : AOI21_X1 port map( B1 => n582, B2 => n137, A => n138, ZN => n135);
   U441 : AOI21_X1 port map( B1 => n139, B2 => n140, A => n550, ZN => n138);
   U442 : AOI22_X1 port map( A1 => n404, A2 => n718, B1 => n684, B2 => R(0), ZN
                           => n399);
   U443 : OAI221_X1 port map( B1 => n685, B2 => n586, C1 => n688, C2 => n584, A
                           => n408, ZN => n404);
   U444 : AOI21_X1 port map( B1 => n593, B2 => n395, A => n409, ZN => n408);
   U445 : AOI21_X1 port map( B1 => n410, B2 => n411, A => n550, ZN => n409);
   U446 : INV_X1 port map( A => n170, ZN => n637);
   U447 : INV_X1 port map( A => n369, ZN => n686);
   U448 : INV_X1 port map( A => n344, ZN => n681);
   U449 : INV_X1 port map( A => n336, ZN => n679);
   U450 : INV_X1 port map( A => n213, ZN => n651);
   U451 : INV_X1 port map( A => n171, ZN => n640);
   U452 : INV_X1 port map( A => n192, ZN => n647);
   U453 : INV_X1 port map( A => n183, ZN => n642);
   U454 : INV_X1 port map( A => n165, ZN => n638);
   U455 : NAND2_X1 port map( A1 => data_in(0), A2 => n398, ZN => n441);
   U456 : NAND2_X1 port map( A1 => data_in(1), A2 => n398, ZN => n440);
   U457 : NAND2_X1 port map( A1 => data_in(2), A2 => n398, ZN => n439);
   U458 : NAND2_X1 port map( A1 => data_in(3), A2 => n398, ZN => n438);
   U459 : NAND2_X1 port map( A1 => data_in(4), A2 => n398, ZN => n437);
   U460 : NAND2_X1 port map( A1 => data_in(5), A2 => n398, ZN => n436);
   U461 : NAND2_X1 port map( A1 => data_in(6), A2 => n398, ZN => n435);
   U462 : INV_X1 port map( A => n176, ZN => n633);
   U463 : INV_X1 port map( A => n352, ZN => n682);
   U464 : INV_X1 port map( A => n320, ZN => n676);
   U465 : INV_X1 port map( A => n312, ZN => n675);
   U466 : INV_X1 port map( A => n304, ZN => n673);
   U467 : INV_X1 port map( A => n296, ZN => n671);
   U468 : INV_X1 port map( A => n280, ZN => n667);
   U469 : INV_X1 port map( A => n288, ZN => n669);
   U470 : INV_X1 port map( A => n272, ZN => n665);
   U471 : INV_X1 port map( A => n264, ZN => n663);
   U472 : INV_X1 port map( A => n256, ZN => n661);
   U473 : INV_X1 port map( A => n248, ZN => n659);
   U474 : INV_X1 port map( A => n240, ZN => n657);
   U475 : INV_X1 port map( A => n232, ZN => n655);
   U476 : INV_X1 port map( A => n224, ZN => n653);
   U477 : INV_X1 port map( A => n208, ZN => n649);
   U478 : INV_X1 port map( A => n193, ZN => n645);
   U479 : INV_X1 port map( A => n328, ZN => n677);
   U480 : NAND2_X1 port map( A1 => data_in(7), A2 => n398, ZN => n427);
   U481 : INV_X1 port map( A => n164, ZN => n635);
   U482 : INV_X1 port map( A => data_in(23), ZN => n727);
   U483 : INV_X1 port map( A => data_in(8), ZN => n742);
   U484 : INV_X1 port map( A => data_in(9), ZN => n741);
   U485 : INV_X1 port map( A => data_in(10), ZN => n740);
   U486 : INV_X1 port map( A => data_in(11), ZN => n739);
   U487 : INV_X1 port map( A => data_in(12), ZN => n738);
   U488 : INV_X1 port map( A => data_in(13), ZN => n737);
   U489 : INV_X1 port map( A => data_in(14), ZN => n736);
   U490 : INV_X1 port map( A => data_in(15), ZN => n735);
   U491 : INV_X1 port map( A => data_in(16), ZN => n734);
   U492 : INV_X1 port map( A => data_in(17), ZN => n733);
   U493 : INV_X1 port map( A => data_in(18), ZN => n732);
   U494 : INV_X1 port map( A => data_in(19), ZN => n731);
   U495 : INV_X1 port map( A => data_in(20), ZN => n730);
   U496 : INV_X1 port map( A => data_in(21), ZN => n729);
   U497 : INV_X1 port map( A => data_in(22), ZN => n728);
   U498 : INV_X1 port map( A => n156, ZN => n632);
   U499 : AND2_X1 port map( A1 => n398, A2 => R(0), ZN => n535);
   U500 : INV_X1 port map( A => n395, ZN => n687);
   U501 : INV_X1 port map( A => n360, ZN => n683);
   U502 : INV_X1 port map( A => n370, ZN => n685);
   U503 : INV_X1 port map( A => n391, ZN => n680);
   U504 : OAI221_X1 port map( B1 => n586, B2 => n388, C1 => n584, C2 => n360, A
                           => n392, ZN => n391);
   U505 : AOI22_X1 port map( A1 => n681, A2 => n546, B1 => n686, B2 => n592, ZN
                           => n392);
   U506 : INV_X1 port map( A => n405, ZN => n684);
   U507 : OAI221_X1 port map( B1 => n584, B2 => n388, C1 => n586, C2 => n360, A
                           => n406, ZN => n405);
   U508 : AOI22_X1 port map( A1 => n686, A2 => n592, B1 => n407, B2 => n548, ZN
                           => n406);
   U509 : INV_X1 port map( A => N35, ZN => n689);
   U510 : INV_X1 port map( A => n400, ZN => n688);
   U511 : AND2_X1 port map( A1 => n442, A2 => data_in(0), ZN => N85);
   U512 : AND2_X1 port map( A1 => n442, A2 => data_in(1), ZN => N86);
   U513 : AND2_X1 port map( A1 => n442, A2 => data_in(2), ZN => N87);
   U514 : AND2_X1 port map( A1 => n442, A2 => data_in(3), ZN => N88);
   U515 : AND2_X1 port map( A1 => n442, A2 => data_in(4), ZN => N89);
   U516 : AND2_X1 port map( A1 => n442, A2 => data_in(5), ZN => N90);
   U517 : AND2_X1 port map( A1 => n442, A2 => data_in(6), ZN => N91);
   U518 : INV_X1 port map( A => n145, ZN => n627);
   U519 : OAI221_X1 port map( B1 => n584, B2 => n633, C1 => n550, C2 => n637, A
                           => n146, ZN => n145);
   U520 : AOI22_X1 port map( A1 => n147, A2 => n592, B1 => n148, B2 => n588, ZN
                           => n146);
   U521 : AND2_X1 port map( A1 => data_in(7), A2 => n442, ZN => N92);
   U522 : INV_X1 port map( A => n398, ZN => n691);
   U523 : NOR2_X2 port map( A1 => conf(1), A2 => conf(0), ZN => n398);
   U524 : NAND2_X1 port map( A1 => n423, A2 => n424, ZN => n360);
   U525 : AOI22_X1 port map( A1 => mask_0_7_port, A2 => n562, B1 => 
                           mask_1_7_port, B2 => n555, ZN => n423);
   U526 : AOI22_X1 port map( A1 => mask_2_7_port, A2 => n577, B1 => 
                           mask_3_7_port, B2 => n571, ZN => n424);
   U527 : NAND2_X1 port map( A1 => n416, A2 => n417, ZN => n370);
   U528 : AOI22_X1 port map( A1 => mask_0_6_port, A2 => n562, B1 => 
                           mask_1_6_port, B2 => n555, ZN => n416);
   U529 : AOI22_X1 port map( A1 => mask_2_6_port, A2 => n577, B1 => 
                           mask_3_6_port, B2 => n571, ZN => n417);
   U530 : NAND2_X1 port map( A1 => n378, A2 => n379, ZN => n328);
   U531 : AOI22_X1 port map( A1 => mask_0_11_port, A2 => n562, B1 => 
                           mask_1_11_port, B2 => n555, ZN => n378);
   U532 : AOI22_X1 port map( A1 => mask_2_11_port, A2 => n577, B1 => 
                           mask_3_11_port, B2 => n571, ZN => n379);
   U533 : NAND2_X1 port map( A1 => n402, A2 => n403, ZN => n352);
   U534 : AOI22_X1 port map( A1 => mask_0_8_port, A2 => n562, B1 => 
                           mask_1_8_port, B2 => n555, ZN => n402);
   U535 : AOI22_X1 port map( A1 => mask_2_8_port, A2 => n577, B1 => 
                           mask_3_8_port, B2 => n571, ZN => n403);
   U536 : NAND2_X1 port map( A1 => n372, A2 => n373, ZN => n320);
   U537 : AOI22_X1 port map( A1 => mask_0_12_port, A2 => n563, B1 => 
                           mask_1_12_port, B2 => n556, ZN => n372);
   U538 : AOI22_X1 port map( A1 => mask_2_12_port, A2 => n578, B1 => 
                           mask_3_12_port, B2 => n572, ZN => n373);
   U539 : NAND2_X1 port map( A1 => n362, A2 => n363, ZN => n312);
   U540 : AOI22_X1 port map( A1 => mask_0_13_port, A2 => n563, B1 => 
                           mask_1_13_port, B2 => n556, ZN => n362);
   U541 : AOI22_X1 port map( A1 => mask_2_13_port, A2 => n578, B1 => 
                           mask_3_13_port, B2 => n572, ZN => n363);
   U542 : NAND2_X1 port map( A1 => n354, A2 => n355, ZN => n304);
   U543 : AOI22_X1 port map( A1 => mask_0_14_port, A2 => n563, B1 => 
                           mask_1_14_port, B2 => n556, ZN => n354);
   U544 : AOI22_X1 port map( A1 => mask_2_14_port, A2 => n578, B1 => 
                           mask_3_14_port, B2 => n572, ZN => n355);
   U545 : NAND2_X1 port map( A1 => n346, A2 => n347, ZN => n296);
   U546 : AOI22_X1 port map( A1 => mask_0_15_port, A2 => n563, B1 => 
                           mask_1_15_port, B2 => n556, ZN => n346);
   U547 : AOI22_X1 port map( A1 => mask_2_15_port, A2 => n578, B1 => 
                           mask_3_15_port, B2 => n572, ZN => n347);
   U548 : NAND2_X1 port map( A1 => n330, A2 => n331, ZN => n280);
   U549 : AOI22_X1 port map( A1 => mask_0_17_port, A2 => n563, B1 => 
                           mask_1_17_port, B2 => n556, ZN => n330);
   U550 : AOI22_X1 port map( A1 => mask_2_17_port, A2 => n578, B1 => 
                           mask_3_17_port, B2 => n572, ZN => n331);
   U551 : NAND2_X1 port map( A1 => n338, A2 => n339, ZN => n288);
   U552 : AOI22_X1 port map( A1 => mask_0_16_port, A2 => n563, B1 => 
                           mask_1_16_port, B2 => n556, ZN => n338);
   U553 : AOI22_X1 port map( A1 => mask_2_16_port, A2 => n578, B1 => 
                           mask_3_16_port, B2 => n572, ZN => n339);
   U554 : NAND2_X1 port map( A1 => n322, A2 => n323, ZN => n272);
   U555 : AOI22_X1 port map( A1 => mask_0_18_port, A2 => n563, B1 => 
                           mask_1_18_port, B2 => n556, ZN => n322);
   U556 : AOI22_X1 port map( A1 => mask_2_18_port, A2 => n578, B1 => 
                           mask_3_18_port, B2 => n572, ZN => n323);
   U557 : NAND2_X1 port map( A1 => n314, A2 => n315, ZN => n264);
   U558 : AOI22_X1 port map( A1 => mask_0_19_port, A2 => n563, B1 => 
                           mask_1_19_port, B2 => n556, ZN => n314);
   U559 : AOI22_X1 port map( A1 => mask_2_19_port, A2 => n578, B1 => 
                           mask_3_19_port, B2 => n572, ZN => n315);
   U560 : NAND2_X1 port map( A1 => n306, A2 => n307, ZN => n256);
   U561 : AOI22_X1 port map( A1 => mask_0_20_port, A2 => n563, B1 => 
                           mask_1_20_port, B2 => n556, ZN => n306);
   U562 : AOI22_X1 port map( A1 => mask_2_20_port, A2 => n578, B1 => 
                           mask_3_20_port, B2 => n572, ZN => n307);
   U563 : NAND2_X1 port map( A1 => n298, A2 => n299, ZN => n248);
   U565 : AOI22_X1 port map( A1 => mask_0_21_port, A2 => n563, B1 => 
                           mask_1_21_port, B2 => n556, ZN => n298);
   U566 : AOI22_X1 port map( A1 => mask_2_21_port, A2 => n578, B1 => 
                           mask_3_21_port, B2 => n572, ZN => n299);
   U567 : NAND2_X1 port map( A1 => n290, A2 => n291, ZN => n240);
   U568 : AOI22_X1 port map( A1 => mask_0_22_port, A2 => n563, B1 => 
                           mask_1_22_port, B2 => n556, ZN => n290);
   U569 : AOI22_X1 port map( A1 => mask_2_22_port, A2 => n578, B1 => 
                           mask_3_22_port, B2 => n572, ZN => n291);
   U570 : NAND2_X1 port map( A1 => n282, A2 => n283, ZN => n232);
   U571 : AOI22_X1 port map( A1 => mask_0_23_port, A2 => n563, B1 => 
                           mask_1_23_port, B2 => n556, ZN => n282);
   U572 : AOI22_X1 port map( A1 => mask_2_23_port, A2 => n578, B1 => 
                           mask_3_23_port, B2 => n572, ZN => n283);
   U573 : NAND2_X1 port map( A1 => n274, A2 => n275, ZN => n224);
   U574 : AOI22_X1 port map( A1 => mask_0_24_port, A2 => n564, B1 => 
                           mask_1_24_port, B2 => n557, ZN => n274);
   U575 : AOI22_X1 port map( A1 => mask_2_24_port, A2 => n579, B1 => 
                           mask_3_24_port, B2 => n573, ZN => n275);
   U576 : NAND2_X1 port map( A1 => n258, A2 => n259, ZN => n208);
   U577 : AOI22_X1 port map( A1 => mask_0_26_port, A2 => n564, B1 => 
                           mask_1_26_port, B2 => n557, ZN => n258);
   U578 : AOI22_X1 port map( A1 => mask_2_26_port, A2 => n579, B1 => 
                           mask_3_26_port, B2 => n573, ZN => n259);
   U579 : NAND2_X1 port map( A1 => n242, A2 => n243, ZN => n193);
   U580 : AOI22_X1 port map( A1 => mask_0_28_port, A2 => n564, B1 => 
                           mask_1_28_port, B2 => n557, ZN => n242);
   U581 : AOI22_X1 port map( A1 => mask_2_28_port, A2 => n579, B1 => 
                           mask_3_28_port, B2 => n573, ZN => n243);
   U582 : NAND2_X1 port map( A1 => n250, A2 => n251, ZN => n192);
   U583 : AOI22_X1 port map( A1 => mask_0_27_port, A2 => n564, B1 => 
                           mask_1_27_port, B2 => n557, ZN => n250);
   U584 : AOI22_X1 port map( A1 => mask_2_27_port, A2 => n579, B1 => 
                           mask_3_27_port, B2 => n573, ZN => n251);
   U585 : NAND2_X1 port map( A1 => n234, A2 => n235, ZN => n183);
   U586 : AOI22_X1 port map( A1 => mask_0_29_port, A2 => n564, B1 => 
                           mask_1_29_port, B2 => n557, ZN => n234);
   U587 : AOI22_X1 port map( A1 => mask_2_29_port, A2 => n579, B1 => 
                           mask_3_29_port, B2 => n573, ZN => n235);
   U588 : NAND2_X1 port map( A1 => n218, A2 => n219, ZN => n165);
   U589 : AOI22_X1 port map( A1 => mask_0_31_port, A2 => n564, B1 => 
                           mask_1_31_port, B2 => n557, ZN => n218);
   U590 : AOI22_X1 port map( A1 => mask_2_31_port, A2 => n579, B1 => 
                           mask_3_31_port, B2 => n573, ZN => n219);
   U591 : NAND2_X1 port map( A1 => n266, A2 => n267, ZN => n213);
   U592 : AOI22_X1 port map( A1 => mask_0_25_port, A2 => n564, B1 => 
                           mask_1_25_port, B2 => n557, ZN => n266);
   U593 : AOI22_X1 port map( A1 => mask_2_25_port, A2 => n579, B1 => 
                           mask_3_25_port, B2 => n573, ZN => n267);
   U594 : NAND2_X1 port map( A1 => n226, A2 => n227, ZN => n171);
   U595 : AOI22_X1 port map( A1 => mask_0_30_port, A2 => n564, B1 => 
                           mask_1_30_port, B2 => n557, ZN => n226);
   U596 : AOI22_X1 port map( A1 => mask_2_30_port, A2 => n579, B1 => 
                           mask_3_30_port, B2 => n573, ZN => n227);
   U597 : AOI22_X1 port map( A1 => mask_2_0_port, A2 => n577, B1 => 
                           mask_3_0_port, B2 => n571, ZN => n411);
   U598 : AOI22_X1 port map( A1 => mask_2_39_port, A2 => n580, B1 => 
                           mask_3_39_port, B2 => n574, ZN => n140);
   U599 : AOI22_X1 port map( A1 => mask_0_0_port, A2 => n562, B1 => 
                           mask_1_0_port, B2 => n555, ZN => n410);
   U600 : AOI22_X1 port map( A1 => mask_0_39_port, A2 => n565, B1 => 
                           mask_1_39_port, B2 => n558, ZN => n139);
   U601 : NAND2_X1 port map( A1 => n385, A2 => n386, ZN => n336);
   U602 : AOI22_X1 port map( A1 => mask_0_10_port, A2 => n562, B1 => 
                           mask_1_10_port, B2 => n555, ZN => n385);
   U603 : AOI22_X1 port map( A1 => mask_2_10_port, A2 => n577, B1 => 
                           mask_3_10_port, B2 => n571, ZN => n386);
   U604 : NAND2_X1 port map( A1 => n393, A2 => n394, ZN => n344);
   U605 : AOI22_X1 port map( A1 => mask_0_9_port, A2 => n562, B1 => 
                           mask_1_9_port, B2 => n555, ZN => n393);
   U606 : AOI22_X1 port map( A1 => mask_2_9_port, A2 => n577, B1 => 
                           mask_3_9_port, B2 => n571, ZN => n394);
   U607 : NAND2_X1 port map( A1 => n201, A2 => n202, ZN => n164);
   U608 : AOI22_X1 port map( A1 => mask_0_33_port, A2 => n564, B1 => 
                           mask_1_33_port, B2 => n557, ZN => n201);
   U609 : AOI22_X1 port map( A1 => mask_2_33_port, A2 => n579, B1 => 
                           mask_3_33_port, B2 => n573, ZN => n202);
   U610 : NAND2_X1 port map( A1 => n210, A2 => n211, ZN => n170);
   U611 : AOI22_X1 port map( A1 => mask_0_32_port, A2 => n564, B1 => 
                           mask_1_32_port, B2 => n557, ZN => n210);
   U612 : AOI22_X1 port map( A1 => mask_2_32_port, A2 => n579, B1 => 
                           mask_3_32_port, B2 => n573, ZN => n211);
   U613 : NAND2_X1 port map( A1 => n177, A2 => n178, ZN => n147);
   U614 : AOI22_X1 port map( A1 => mask_0_36_port, A2 => n565, B1 => 
                           mask_1_36_port, B2 => n558, ZN => n177);
   U615 : AOI22_X1 port map( A1 => mask_2_36_port, A2 => n580, B1 => 
                           mask_3_36_port, B2 => n574, ZN => n178);
   U616 : NAND2_X1 port map( A1 => n425, A2 => n426, ZN => n388);
   U617 : AOI22_X1 port map( A1 => mask_0_3_port, A2 => n562, B1 => 
                           mask_1_3_port, B2 => n555, ZN => n425);
   U618 : AOI22_X1 port map( A1 => mask_2_3_port, A2 => n577, B1 => 
                           mask_3_3_port, B2 => n571, ZN => n426);
   U619 : NAND2_X1 port map( A1 => n412, A2 => n413, ZN => n395);
   U620 : AOI22_X1 port map( A1 => mask_0_4_port, A2 => n562, B1 => 
                           mask_1_4_port, B2 => n555, ZN => n412);
   U621 : AOI22_X1 port map( A1 => mask_2_4_port, A2 => n577, B1 => 
                           mask_3_4_port, B2 => n571, ZN => n413);
   U622 : NAND2_X1 port map( A1 => n167, A2 => n168, ZN => n137);
   U623 : AOI22_X1 port map( A1 => mask_0_37_port, A2 => n565, B1 => 
                           mask_1_37_port, B2 => n558, ZN => n167);
   U624 : AOI22_X1 port map( A1 => mask_2_37_port, A2 => n580, B1 => 
                           mask_3_37_port, B2 => n574, ZN => n168);
   U625 : NAND2_X1 port map( A1 => n185, A2 => n186, ZN => n156);
   U626 : AOI22_X1 port map( A1 => mask_0_35_port, A2 => n564, B1 => 
                           mask_1_35_port, B2 => n557, ZN => n185);
   U627 : AOI22_X1 port map( A1 => mask_2_35_port, A2 => n579, B1 => 
                           mask_3_35_port, B2 => n573, ZN => n186);
   U628 : NAND2_X1 port map( A1 => n195, A2 => n196, ZN => n176);
   U629 : AOI22_X1 port map( A1 => mask_0_34_port, A2 => n564, B1 => 
                           mask_1_34_port, B2 => n557, ZN => n195);
   U630 : AOI22_X1 port map( A1 => mask_2_34_port, A2 => n579, B1 => 
                           mask_3_34_port, B2 => n573, ZN => n196);
   U631 : NAND2_X1 port map( A1 => n419, A2 => n420, ZN => n369);
   U632 : AOI22_X1 port map( A1 => mask_0_5_port, A2 => n562, B1 => 
                           mask_1_5_port, B2 => n555, ZN => n419);
   U633 : AOI22_X1 port map( A1 => mask_2_5_port, A2 => n577, B1 => 
                           mask_3_5_port, B2 => n571, ZN => n420);
   U634 : NAND2_X1 port map( A1 => n414, A2 => n415, ZN => n400);
   U635 : AOI22_X1 port map( A1 => mask_0_2_port, A2 => n562, B1 => 
                           mask_1_2_port, B2 => n555, ZN => n414);
   U636 : AOI22_X1 port map( A1 => mask_2_2_port, A2 => n577, B1 => 
                           mask_3_2_port, B2 => n571, ZN => n415);
   U637 : NAND2_X1 port map( A1 => n154, A2 => n155, ZN => n148);
   U638 : AOI22_X1 port map( A1 => mask_0_38_port, A2 => n565, B1 => 
                           mask_3_38_port, B2 => n574, ZN => n154);
   U639 : AOI22_X1 port map( A1 => mask_2_38_port, A2 => n580, B1 => 
                           mask_1_38_port, B2 => n558, ZN => n155);
   U640 : NAND2_X1 port map( A1 => n599, A2 => n443, ZN => N35);
   U641 : AND2_X1 port map( A1 => n421, A2 => n422, ZN => n407);
   U642 : AOI22_X1 port map( A1 => mask_0_1_port, A2 => n562, B1 => 
                           mask_3_1_port, B2 => n571, ZN => n421);
   U643 : AOI22_X1 port map( A1 => mask_2_1_port, A2 => n577, B1 => 
                           mask_1_1_port, B2 => n555, ZN => n422);
   U644 : INV_X1 port map( A => conf(1), ZN => n690);
   U645 : BUF_X1 port map( A => n9, Z => n603);
   U646 : NOR3_X1 port map( A1 => n719, A2 => conf(0), A3 => n690, ZN => n9);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_4_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3, n4, n8, n12, n13, n14 : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(1), B => n14, Z => n4);
   U6 : XOR2_X1 port map( A => B(5), B => n14, Z => n3);
   U7 : XOR2_X1 port map( A => B(2), B => n14, Z => n2);
   U8 : XOR2_X1 port map( A => B(3), B => n14, Z => n1);
   U9 : XOR2_X1 port map( A => B(9), B => n14, Z => B_in_9_port);
   U10 : XOR2_X1 port map( A => B(8), B => n14, Z => B_in_8_port);
   U11 : XOR2_X1 port map( A => B(7), B => n14, Z => B_in_7_port);
   U12 : XOR2_X1 port map( A => B(6), B => n13, Z => B_in_6_port);
   U13 : XOR2_X1 port map( A => B(4), B => n13, Z => B_in_4_port);
   U14 : XOR2_X1 port map( A => B(31), B => n13, Z => B_in_31_port);
   U15 : XOR2_X1 port map( A => B(30), B => n13, Z => B_in_30_port);
   U16 : XOR2_X1 port map( A => B(29), B => n13, Z => B_in_29_port);
   U17 : XOR2_X1 port map( A => B(28), B => n13, Z => B_in_28_port);
   U18 : XOR2_X1 port map( A => B(27), B => n13, Z => B_in_27_port);
   U19 : XOR2_X1 port map( A => B(26), B => n13, Z => B_in_26_port);
   U20 : XOR2_X1 port map( A => B(25), B => n13, Z => B_in_25_port);
   U21 : XOR2_X1 port map( A => B(24), B => n13, Z => B_in_24_port);
   U22 : XOR2_X1 port map( A => B(23), B => n13, Z => B_in_23_port);
   U23 : XOR2_X1 port map( A => B(22), B => n12, Z => B_in_22_port);
   U24 : XOR2_X1 port map( A => B(21), B => n12, Z => B_in_21_port);
   U25 : XOR2_X1 port map( A => B(20), B => n12, Z => B_in_20_port);
   U26 : XOR2_X1 port map( A => B(19), B => n12, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => n12, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => n13, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => n12, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => n12, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => n12, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => n12, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => n12, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => n12, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => n12, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => n14, B => B(0), Z => n8);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => n3, B(4) 
                           => B_in_4_port, B(3) => n1, B(2) => n2, B(1) => n4, 
                           B(0) => n8, Cin => C_internal, Co(8) => Cout, Co(7) 
                           => carry_7_port, Co(6) => carry_6_port, Co(5) => 
                           carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => n3, B(4) => B_in_4_port, B(3) 
                           => n1, B(2) => n2, B(1) => n4, B(0) => n8, Ci(7) => 
                           carry_7_port, Ci(6) => carry_6_port, Ci(5) => 
                           carry_5_port, Ci(4) => carry_4_port, Ci(3) => 
                           carry_3_port, Ci(2) => carry_2_port, Ci(1) => 
                           carry_1_port, Ci(0) => carry_0_port, S(31) => S(31),
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U4 : BUF_X1 port map( A => ADD_SUB, Z => n12);
   U37 : BUF_X1 port map( A => ADD_SUB, Z => n13);
   U38 : BUF_X1 port map( A => ADD_SUB, Z => n14);
   U39 : OR2_X1 port map( A1 => n14, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_41;

architecture SYN_Behavioral of AND2_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_0;

architecture SYN_Behavioral of AND2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_1_DW01_add_0_DW01_add_128 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_adder_1_DW01_add_0_DW01_add_128;

architecture SYN_rpl of PC_adder_1_DW01_add_0_DW01_add_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1530 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1530, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_0_DW01_add_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_adder_0_DW01_add_2;

architecture SYN_cla of PC_adder_0_DW01_add_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n29, n31, n32, n33, n34
      , n36, n37, n40, n41, n42, n43, n44, n45, n46, n48, n49, n51, n52, n53, 
      n54, n55, n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69
      , n70, n71, n73, n74, n76, n77, n78, n79, n80, n81, n82, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98, n99, n101, n102, 
      n103, n104, n105, n106, n107, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n120, n121, n122, n124, n125, n126, n128, n129, n130, 
      n131, n132, n133, n134, n135, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n149, n150, n152, n153, n154, n155, n157, n159, n160, 
      n162, n163, n164, n165, n167, n168, n169, n170, n171, n172, n173, n174, 
      n176, n177, n180, n181, n184, n185, n186, n188, n189, n191, n193, n194, 
      n197, n198, n200, n201, n202, n204, n208, n209, n210, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => n51, B => n60, Z => SUM(29));
   U124 : XOR2_X1 port map( A => B(31), B => A(31), Z => n5);
   U205 : NAND3_X1 port map( A1 => n73, A2 => n79, A3 => n78, ZN => n67);
   U209 : NAND3_X1 port map( A1 => n98, A2 => n104, A3 => n103, ZN => n92);
   U216 : NAND3_X1 port map( A1 => n125, A2 => n124, A3 => n130, ZN => n117);
   U2 : AND2_X1 port map( A1 => n133, A2 => n208, ZN => SUM(0));
   U3 : INV_X1 port map( A => n169, ZN => n224);
   U4 : OAI21_X1 port map( B1 => n229, B2 => n169, A => n222, ZN => n13);
   U5 : OR2_X1 port map( A1 => n165, A2 => n215, ZN => n180);
   U6 : AND2_X1 port map( A1 => n4, A2 => n13, ZN => n215);
   U7 : INV_X1 port map( A => n138, ZN => n218);
   U8 : INV_X1 port map( A => n197, ZN => n219);
   U9 : INV_X1 port map( A => n41, ZN => n242);
   U10 : NOR2_X1 port map( A1 => n244, A2 => n120, ZN => n118);
   U11 : INV_X1 port map( A => n131, ZN => n244);
   U12 : NOR2_X1 port map( A1 => n6, A2 => n94, ZN => n93);
   U13 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n238, ZN => n94);
   U14 : NOR2_X1 port map( A1 => n7, A2 => n69, ZN => n68);
   U15 : AOI21_X1 port map( B1 => n70, B2 => n71, A => n235, ZN => n69);
   U16 : OAI21_X1 port map( B1 => n209, B2 => n230, A => n43, ZN => n168);
   U17 : INV_X1 port map( A => n42, ZN => n230);
   U18 : INV_X1 port map( A => n40, ZN => n233);
   U19 : XNOR2_X1 port map( A => n2, B => n49, ZN => SUM(30));
   U20 : NAND2_X1 port map( A1 => n48, A2 => n46, ZN => n49);
   U21 : OAI21_X1 port map( B1 => n241, B2 => n133, A => n56, ZN => n210);
   U22 : INV_X1 port map( A => n57, ZN => n241);
   U23 : AND2_X1 port map( A1 => n61, A2 => n62, ZN => n51);
   U24 : NOR2_X1 port map( A1 => n235, A2 => n7, ZN => n81);
   U25 : AOI21_X1 port map( B1 => n73, B2 => n82, A => n236, ZN => n80);
   U26 : INV_X1 port map( A => n71, ZN => n236);
   U27 : NAND2_X1 port map( A1 => n66, A2 => n76, ZN => n86);
   U28 : NAND2_X1 port map( A1 => n85, A2 => n77, ZN => n82);
   U29 : NAND2_X1 port map( A1 => n78, A2 => n86, ZN => n85);
   U30 : NAND4_X1 port map( A1 => n32, A2 => n33, A3 => n20, A4 => n22, ZN => 
                           n169);
   U31 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n60);
   U32 : XNOR2_X1 port map( A => n82, B => n84, ZN => SUM(26));
   U33 : NAND2_X1 port map( A1 => n71, A2 => n73, ZN => n84);
   U34 : OAI21_X1 port map( B1 => n216, B2 => n250, A => n160, ZN => n173);
   U35 : INV_X1 port map( A => n176, ZN => n216);
   U36 : OAI21_X1 port map( B1 => n251, B2 => n217, A => n159, ZN => n176);
   U37 : INV_X1 port map( A => n162, ZN => n251);
   U38 : INV_X1 port map( A => n180, ZN => n217);
   U39 : XNOR2_X1 port map( A => n170, B => n171, ZN => SUM(15));
   U41 : NAND2_X1 port map( A1 => n152, A2 => n153, ZN => n170);
   U42 : NAND2_X1 port map( A1 => n172, A2 => n157, ZN => n171);
   U43 : NAND2_X1 port map( A1 => n154, A2 => n173, ZN => n172);
   U44 : XNOR2_X1 port map( A => n105, B => n106, ZN => SUM(23));
   U45 : NOR2_X1 port map( A1 => n238, A2 => n6, ZN => n106);
   U46 : AOI21_X1 port map( B1 => n98, B2 => n107, A => n239, ZN => n105);
   U47 : INV_X1 port map( A => n96, ZN => n239);
   U48 : NAND2_X1 port map( A1 => n110, A2 => n102, ZN => n107);
   U49 : NAND2_X1 port map( A1 => n103, A2 => n111, ZN => n110);
   U50 : AND4_X1 port map( A1 => n184, A2 => n185, A3 => n10, A4 => n15, ZN => 
                           n4);
   U51 : NAND2_X1 port map( A1 => n62, A2 => n64, ZN => n65);
   U52 : XNOR2_X1 port map( A => n87, B => n86, ZN => SUM(25));
   U53 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n87);
   U54 : XNOR2_X1 port map( A => n174, B => n173, ZN => SUM(14));
   U55 : NAND2_X1 port map( A1 => n157, A2 => n154, ZN => n174);
   U56 : XNOR2_X1 port map( A => n107, B => n109, ZN => SUM(22));
   U57 : NAND2_X1 port map( A1 => n96, A2 => n98, ZN => n109);
   U58 : XNOR2_X1 port map( A => n134, B => n135, ZN => SUM(19));
   U59 : NAND2_X1 port map( A1 => n131, A2 => n124, ZN => n134);
   U60 : OAI21_X1 port map( B1 => n218, B2 => n245, A => n122, ZN => n135);
   U61 : INV_X1 port map( A => n125, ZN => n245);
   U62 : NAND2_X1 port map( A1 => n140, A2 => n129, ZN => n138);
   U63 : NAND2_X1 port map( A1 => n130, A2 => n141, ZN => n140);
   U64 : OAI21_X1 port map( B1 => n220, B2 => n221, A => n11, ZN => n197);
   U65 : INV_X1 port map( A => n9, ZN => n221);
   U66 : XNOR2_X1 port map( A => n193, B => n194, ZN => SUM(11));
   U67 : NAND2_X1 port map( A1 => n188, A2 => n184, ZN => n193);
   U68 : OAI21_X1 port map( B1 => n219, B2 => n253, A => n191, ZN => n194);
   U69 : INV_X1 port map( A => n185, ZN => n253);
   U70 : NAND2_X1 port map( A1 => n200, A2 => n14, ZN => n9);
   U71 : NAND2_X1 port map( A1 => n13, A2 => n15, ZN => n200);
   U72 : NAND4_X1 port map( A1 => n162, A2 => n163, A3 => n154, A4 => n153, ZN 
                           => n147);
   U73 : NAND2_X1 port map( A1 => n76, A2 => n89, ZN => n90);
   U74 : XNOR2_X1 port map( A => n112, B => n111, ZN => SUM(21));
   U75 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => n112);
   U76 : XNOR2_X1 port map( A => n177, B => n176, ZN => SUM(13));
   U77 : NAND2_X1 port map( A1 => n160, A2 => n163, ZN => n177);
   U78 : XNOR2_X1 port map( A => n198, B => n197, ZN => SUM(10));
   U79 : NAND2_X1 port map( A1 => n191, A2 => n185, ZN => n198);
   U80 : XNOR2_X1 port map( A => n139, B => n138, ZN => SUM(18));
   U81 : NAND2_X1 port map( A1 => n122, A2 => n125, ZN => n139);
   U82 : OAI21_X1 port map( B1 => n227, B2 => n226, A => n27, ZN => n21);
   U83 : INV_X1 port map( A => n28, ZN => n227);
   U84 : OAI21_X1 port map( B1 => n228, B2 => n229, A => n31, ZN => n28);
   U85 : INV_X1 port map( A => n32, ZN => n228);
   U86 : XNOR2_X1 port map( A => n16, B => n17, ZN => SUM(7));
   U87 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n16);
   U88 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n17);
   U89 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n18);
   U90 : NAND2_X1 port map( A1 => n101, A2 => n114, ZN => n115);
   U91 : XNOR2_X1 port map( A => n142, B => n141, ZN => SUM(17));
   U92 : NAND2_X1 port map( A1 => n129, A2 => n130, ZN => n142);
   U93 : XNOR2_X1 port map( A => n24, B => n21, ZN => SUM(6));
   U94 : NAND2_X1 port map( A1 => n20, A2 => n19, ZN => n24);
   U95 : XNOR2_X1 port map( A => n181, B => n180, ZN => SUM(12));
   U96 : NAND2_X1 port map( A1 => n159, A2 => n162, ZN => n181);
   U97 : XNOR2_X1 port map( A => n8, B => n9, ZN => SUM(9));
   U98 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => n8);
   U99 : XNOR2_X1 port map( A => n145, B => n1, ZN => SUM(16));
   U100 : NAND2_X1 port map( A1 => n128, A2 => n144, ZN => n145);
   U101 : XNOR2_X1 port map( A => n12, B => n13, ZN => SUM(8));
   U102 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n12);
   U103 : XNOR2_X1 port map( A => n29, B => n28, ZN => SUM(5));
   U104 : NAND2_X1 port map( A1 => n33, A2 => n27, ZN => n29);
   U105 : XNOR2_X1 port map( A => n36, B => n37, ZN => SUM(3));
   U106 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => n36);
   U107 : OAI21_X1 port map( B1 => n242, B2 => n232, A => n40, ZN => n37);
   U108 : INV_X1 port map( A => n59, ZN => n232);
   U109 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n41);
   U110 : NAND2_X1 port map( A1 => n57, A2 => n255, ZN => n55);
   U111 : INV_X1 port map( A => n133, ZN => n255);
   U112 : INV_X1 port map( A => n163, ZN => n250);
   U113 : INV_X1 port map( A => n33, ZN => n226);
   U114 : INV_X1 port map( A => n10, ZN => n220);
   U115 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => n34);
   U116 : XNOR2_X1 port map( A => n54, B => n41, ZN => SUM(2));
   U117 : NAND2_X1 port map( A1 => n59, A2 => n40, ZN => n54);
   U118 : INV_X1 port map( A => n53, ZN => n234);
   U119 : INV_X1 port map( A => n104, ZN => n238);
   U120 : INV_X1 port map( A => n79, ZN => n235);
   U121 : XNOR2_X1 port map( A => n132, B => n255, ZN => SUM(1));
   U122 : NAND2_X1 port map( A1 => n57, A2 => n56, ZN => n132);
   U123 : OAI21_X1 port map( B1 => n186, B2 => n252, A => n188, ZN => n165);
   U125 : INV_X1 port map( A => n184, ZN => n252);
   U126 : AOI21_X1 port map( B1 => n185, B2 => n189, A => n254, ZN => n186);
   U127 : INV_X1 port map( A => n191, ZN => n254);
   U128 : AOI21_X1 port map( B1 => n121, B2 => n122, A => n243, ZN => n120);
   U129 : INV_X1 port map( A => n124, ZN => n243);
   U130 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n121);
   U131 : OAI21_X1 port map( B1 => n246, B2 => n128, A => n129, ZN => n126);
   U132 : OAI21_X1 port map( B1 => n226, B2 => n31, A => n27, ZN => n204);
   U133 : OAI21_X1 port map( B1 => n220, B2 => n14, A => n11, ZN => n189);
   U134 : OAI21_X1 port map( B1 => n250, B2 => n159, A => n160, ZN => n155);
   U135 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => n70);
   U136 : OAI21_X1 port map( B1 => n237, B2 => n76, A => n77, ZN => n74);
   U137 : INV_X1 port map( A => n78, ZN => n237);
   U138 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => n95);
   U139 : OAI21_X1 port map( B1 => n240, B2 => n101, A => n102, ZN => n99);
   U140 : INV_X1 port map( A => n103, ZN => n240);
   U141 : INV_X1 port map( A => n201, ZN => n222);
   U142 : OAI21_X1 port map( B1 => n202, B2 => n223, A => n23, ZN => n201);
   U143 : INV_X1 port map( A => n22, ZN => n223);
   U144 : AOI21_X1 port map( B1 => n20, B2 => n204, A => n225, ZN => n202);
   U145 : INV_X1 port map( A => n130, ZN => n246);
   U146 : INV_X1 port map( A => n149, ZN => n247);
   U147 : OAI21_X1 port map( B1 => n150, B2 => n248, A => n152, ZN => n149);
   U148 : INV_X1 port map( A => n153, ZN => n248);
   U149 : AOI21_X1 port map( B1 => n154, B2 => n155, A => n249, ZN => n150);
   U150 : INV_X1 port map( A => n19, ZN => n225);
   U151 : INV_X1 port map( A => n157, ZN => n249);
   U152 : OR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n57);
   U153 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n133);
   U154 : INV_X1 port map( A => n48, ZN => n231);
   U155 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n22);
   U156 : OR2_X1 port map( A1 => B(5), A2 => A(5), ZN => n33);
   U157 : OR2_X1 port map( A1 => B(6), A2 => A(6), ZN => n20);
   U158 : OR2_X1 port map( A1 => B(3), A2 => A(3), ZN => n42);
   U159 : OR2_X1 port map( A1 => B(4), A2 => A(4), ZN => n32);
   U160 : OR2_X1 port map( A1 => B(2), A2 => A(2), ZN => n59);
   U161 : OR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n185);
   U162 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U163 : OR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n10);
   U164 : OR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n184);
   U165 : OR2_X1 port map( A1 => B(14), A2 => A(14), ZN => n154);
   U166 : OR2_X1 port map( A1 => B(15), A2 => A(15), ZN => n153);
   U167 : OR2_X1 port map( A1 => B(13), A2 => A(13), ZN => n163);
   U168 : OR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n162);
   U169 : OR2_X1 port map( A1 => B(17), A2 => A(17), ZN => n130);
   U170 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n125);
   U171 : OR2_X1 port map( A1 => B(19), A2 => A(19), ZN => n124);
   U172 : OR2_X1 port map( A1 => B(16), A2 => A(16), ZN => n144);
   U173 : OR2_X1 port map( A1 => B(21), A2 => A(21), ZN => n103);
   U174 : OR2_X1 port map( A1 => B(22), A2 => A(22), ZN => n98);
   U175 : OR2_X1 port map( A1 => B(23), A2 => A(23), ZN => n104);
   U176 : OR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n114);
   U177 : OR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n78);
   U178 : OR2_X1 port map( A1 => B(26), A2 => A(26), ZN => n73);
   U179 : OR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n89);
   U180 : OR2_X1 port map( A1 => B(27), A2 => A(27), ZN => n79);
   U181 : OR2_X1 port map( A1 => B(28), A2 => A(28), ZN => n64);
   U182 : OR2_X1 port map( A1 => B(29), A2 => A(29), ZN => n53);
   U183 : OR2_X1 port map( A1 => B(30), A2 => A(30), ZN => n46);
   U184 : OR2_X1 port map( A1 => B(0), A2 => A(0), ZN => n208);
   U185 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n19);
   U186 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n56);
   U187 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n40);
   U188 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n76);
   U189 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U190 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n27);
   U191 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U192 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n96);
   U193 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => n71);
   U194 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n157);
   U195 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n122);
   U196 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n102);
   U197 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n77);
   U198 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n129);
   U199 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n31);
   U200 : NAND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n159);
   U201 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n191);
   U202 : NAND2_X1 port map( A1 => B(13), A2 => A(13), ZN => n160);
   U203 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n128);
   U204 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n101);
   U206 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n52);
   U207 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n43);
   U208 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n23);
   U210 : NAND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n48);
   U211 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n131);
   U212 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n188);
   U213 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n152);
   U214 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n6);
   U215 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => n7);
   U217 : NAND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n62);
   U218 : NAND2_X1 port map( A1 => n116, A2 => n128, ZN => n141);
   U219 : NAND2_X1 port map( A1 => n143, A2 => n144, ZN => n116);
   U220 : OAI21_X1 port map( B1 => n116, B2 => n117, A => n118, ZN => n113);
   U221 : NAND2_X1 port map( A1 => n91, A2 => n101, ZN => n111);
   U222 : OAI21_X1 port map( B1 => n234, B2 => n51, A => n52, ZN => n2);
   U223 : NAND2_X1 port map( A1 => n222, A2 => n167, ZN => n164);
   U224 : AOI21_X1 port map( B1 => n59, B2 => n210, A => n233, ZN => n209);
   U225 : XNOR2_X1 port map( A => n80, B => n81, ZN => SUM(27));
   U226 : OAI21_X1 port map( B1 => n234, B2 => n51, A => n52, ZN => n45);
   U227 : XNOR2_X1 port map( A => n88, B => n90, ZN => SUM(24));
   U228 : XNOR2_X1 port map( A => n63, B => n65, ZN => SUM(28));
   U229 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => n61);
   U230 : AOI21_X1 port map( B1 => n4, B2 => n164, A => n165, ZN => n146);
   U231 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n63);
   U232 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => n66);
   U233 : OAI21_X1 port map( B1 => n91, B2 => n92, A => n93, ZN => n88);
   U234 : AOI21_X1 port map( B1 => n45, B2 => n46, A => n231, ZN => n44);
   U235 : XNOR2_X1 port map( A => n115, B => n113, ZN => SUM(20));
   U236 : XNOR2_X1 port map( A => n34, B => n168, ZN => SUM(4));
   U237 : XNOR2_X1 port map( A => n44, B => n5, ZN => SUM(31));
   U238 : OAI21_X1 port map( B1 => n146, B2 => n147, A => n247, ZN => n1);
   U239 : NAND2_X1 port map( A1 => n113, A2 => n114, ZN => n91);
   U240 : INV_X1 port map( A => n168, ZN => n229);
   U241 : OAI21_X1 port map( B1 => n146, B2 => n147, A => n247, ZN => n143);
   U242 : NAND2_X1 port map( A1 => n224, A2 => n168, ZN => n167);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_NBIT32_NREG32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_NBIT32_NREG32;

architecture SYN_BEHAVIORAL of RF_NBIT32_NREG32 is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N128, N129, N130, N131, N132, 
      N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, 
      N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, 
      N157, N158, N159, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
      N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, 
      N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N291, 
      N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, 
      N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, 
      N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, 
      N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, 
      N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, 
      N352, N353, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n934, n935, n936, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
      n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1449, n1450, n1451, 
      n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, 
      n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, 
      n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
      n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
      n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, 
      n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, 
      n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, 
      n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
      n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, 
      n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, 
      n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, 
      n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, 
      n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
      n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
      n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, 
      n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
      n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, 
      n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, 
      n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, 
      n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
      n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
      n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, 
      n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, 
      n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
      n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, 
      n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
      n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
      n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, 
      n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, 
      n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, 
      n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, 
      n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, 
      n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
      n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
      n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, 
      n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, 
      n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, 
      n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, 
      n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, 
      n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
      n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, 
      n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, 
      n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
      n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
      n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, 
      n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, 
      n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
      n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, 
      n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, 
      n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, 
      n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
      n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
      n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
      n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, 
      n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, 
      n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
      n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, 
      n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, 
      n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, 
      n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, 
      n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, 
      n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
      n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, 
      n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
      n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, 
      n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
      n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, 
      n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
      n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, 
      n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
      n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
      n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, 
      n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
      n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
      n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, 
      n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, 
      n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, 
      n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
      n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, 
      n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
      n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, 
      n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, 
      n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, 
      n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
      n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, 
      n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, 
      n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
      n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
      n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, 
      n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, 
      n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, 
      n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
      n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, 
      n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
      n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, 
      n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, 
      n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
      n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
      n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, 
      n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, 
      n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, 
      n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, 
      n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, 
      n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
      n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
      n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
      n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
      n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, 
      n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, 
      n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
      n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
      n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
      n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
      n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
      n3214, n3215, n3216, n3217, n3218, n3219, n3220 : std_logic;

begin
   
   OUT1_reg_31_inst : DLH_X1 port map( G => CLK, D => N256, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => CLK, D => N255, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => CLK, D => N254, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => CLK, D => N253, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => CLK, D => N252, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => CLK, D => N251, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => CLK, D => N250, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => CLK, D => N249, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => CLK, D => N248, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => CLK, D => N247, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => CLK, D => N246, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => CLK, D => N245, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => CLK, D => N244, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => CLK, D => N243, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => CLK, D => N242, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => CLK, D => N241, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => CLK, D => N240, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => CLK, D => N239, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => CLK, D => N238, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => CLK, D => N237, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => CLK, D => N236, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => CLK, D => N235, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => CLK, D => N234, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => CLK, D => N233, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => CLK, D => N232, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => CLK, D => N231, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => CLK, D => N230, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => CLK, D => N229, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => CLK, D => N228, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => CLK, D => N227, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => CLK, D => N226, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => CLK, D => N225, Q => OUT1(0));
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => N353, D => n2208, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => N353, D => n2212, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => N353, D => n2216, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => N353, D => n2220, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => N353, D => n2224, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N353, D => n2228, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => N353, D => n2232, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => N353, D => n2236, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => N353, D => n2240, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => N353, D => n2244, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => N353, D => n2248, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => N353, D => n2252, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => N353, D => n2256, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => N353, D => n2260, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => N353, D => n2264, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => N353, D => n2268, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N353, D => n2272, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => N353, D => n2276, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N353, D => n2280, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N353, D => n2284, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => N353, D => n2288, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => N353, D => n2292, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => N353, D => n2296, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => N353, D => n2300, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => N353, D => n2304, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => N353, D => n2308, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => N353, D => n2312, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => N353, D => n2316, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => N353, D => n2320, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => N353, D => n2324, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => N353, D => n2328, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => N353, D => n2332, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => N352, D => n2208, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => N352, D => n2212, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => N352, D => n2216, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => N352, D => n2220, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => N352, D => n2224, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => N352, D => n2228, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => N352, D => n2232, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => N352, D => n2236, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => N352, D => n2240, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => N352, D => n2244, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => N352, D => n2248, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => N352, D => n2252, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => N352, D => n2256, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => N352, D => n2260, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => N352, D => n2264, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N352, D => n2268, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => N352, D => n2272, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N352, D => n2276, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N352, D => n2280, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N352, D => n2284, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => N352, D => n2288, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => N352, D => n2292, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => N352, D => n2296, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => N352, D => n2300, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => N352, D => n2304, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => N352, D => n2308, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => N352, D => n2312, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => N352, D => n2316, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => N352, D => n2320, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => N352, D => n2324, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => N352, D => n2328, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => N352, D => n2332, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => N351, D => n2208, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => N351, D => n2212, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => N351, D => n2216, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => N351, D => n2220, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => N351, D => n2224, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => N351, D => n2228, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => N351, D => n2232, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => N351, D => n2236, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => N351, D => n2240, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => N351, D => n2244, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => N351, D => n2248, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => N351, D => n2252, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => N351, D => n2256, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => N351, D => n2260, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => N351, D => n2264, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N351, D => n2268, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => N351, D => n2272, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N351, D => n2276, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N351, D => n2280, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N351, D => n2284, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => N351, D => n2288, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => N351, D => n2292, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => N351, D => n2296, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => N351, D => n2300, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => N351, D => n2304, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => N351, D => n2308, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => N351, D => n2312, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => N351, D => n2316, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => N351, D => n2320, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => N351, D => n2324, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => N351, D => n2328, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => N351, D => n2332, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => N350, D => n2208, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => N350, D => n2212, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => N350, D => n2216, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => N350, D => n2220, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => N350, D => n2224, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => N350, D => n2228, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => N350, D => n2232, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => N350, D => n2236, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => N350, D => n2240, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => N350, D => n2244, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => N350, D => n2248, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => N350, D => n2252, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => N350, D => n2256, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => N350, D => n2260, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => N350, D => n2264, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N350, D => n2268, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => N350, D => n2272, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N350, D => n2276, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N350, D => n2280, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N350, D => n2284, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => N350, D => n2288, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => N350, D => n2292, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => N350, D => n2296, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => N350, D => n2300, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => N350, D => n2304, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => N350, D => n2308, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => N350, D => n2312, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => N350, D => n2316, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => N350, D => n2320, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => N350, D => n2324, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => N350, D => n2328, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => N350, D => n2332, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => N349, D => n2208, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => N349, D => n2212, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => N349, D => n2216, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => N349, D => n2220, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => N349, D => n2224, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => N349, D => n2228, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => N349, D => n2232, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => N349, D => n2236, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => N349, D => n2240, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => N349, D => n2244, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => N349, D => n2248, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => N349, D => n2252, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => N349, D => n2256, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => N349, D => n2260, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => N349, D => n2264, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N349, D => n2268, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => N349, D => n2272, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N349, D => n2276, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N349, D => n2280, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N349, D => n2284, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => N349, D => n2288, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => N349, D => n2292, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => N349, D => n2296, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => N349, D => n2300, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => N349, D => n2304, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => N349, D => n2308, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => N349, D => n2312, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => N349, D => n2316, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => N349, D => n2320, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => N349, D => n2324, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => N349, D => n2328, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => N349, D => n2332, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => N348, D => n2208, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => N348, D => n2212, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => N348, D => n2216, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => N348, D => n2220, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => N348, D => n2224, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => N348, D => n2228, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => N348, D => n2232, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => N348, D => n2236, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => N348, D => n2240, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => N348, D => n2244, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => N348, D => n2248, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => N348, D => n2252, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => N348, D => n2256, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => N348, D => n2260, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => N348, D => n2264, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N348, D => n2268, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => N348, D => n2272, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N348, D => n2276, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N348, D => n2280, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N348, D => n2284, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => N348, D => n2288, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => N348, D => n2292, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => N348, D => n2296, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => N348, D => n2300, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => N348, D => n2304, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => N348, D => n2308, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => N348, D => n2312, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => N348, D => n2316, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => N348, D => n2320, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => N348, D => n2324, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => N348, D => n2328, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => N348, D => n2332, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => N347, D => n2208, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => N347, D => n2212, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => N347, D => n2216, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => N347, D => n2220, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => N347, D => n2224, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => N347, D => n2228, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => N347, D => n2232, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => N347, D => n2236, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => N347, D => n2240, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => N347, D => n2244, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => N347, D => n2248, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => N347, D => n2252, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => N347, D => n2256, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => N347, D => n2260, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => N347, D => n2264, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N347, D => n2268, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => N347, D => n2272, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N347, D => n2276, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N347, D => n2280, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N347, D => n2284, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => N347, D => n2288, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => N347, D => n2292, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => N347, D => n2296, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => N347, D => n2300, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => N347, D => n2304, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => N347, D => n2308, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => N347, D => n2312, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => N347, D => n2316, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => N347, D => n2320, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => N347, D => n2324, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => N347, D => n2328, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => N347, D => n2332, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => N346, D => n2208, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => N346, D => n2212, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => N346, D => n2216, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => N346, D => n2220, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => N346, D => n2224, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => N346, D => n2228, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => N346, D => n2232, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => N346, D => n2236, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => N346, D => n2240, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => N346, D => n2244, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => N346, D => n2248, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => N346, D => n2252, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => N346, D => n2256, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => N346, D => n2260, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => N346, D => n2264, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => N346, D => n2268, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => N346, D => n2272, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N346, D => n2276, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N346, D => n2280, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N346, D => n2284, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => N346, D => n2288, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => N346, D => n2292, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => N346, D => n2296, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => N346, D => n2300, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => N346, D => n2304, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => N346, D => n2308, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => N346, D => n2312, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => N346, D => n2316, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => N346, D => n2320, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => N346, D => n2324, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => N346, D => n2328, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N346, D => n2332, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => N345, D => n2208, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => N345, D => n2212, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => N345, D => n2216, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => N345, D => n2220, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => N345, D => n2224, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => N345, D => n2228, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => N345, D => n2232, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => N345, D => n2236, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => N345, D => n2240, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => N345, D => n2244, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => N345, D => n2248, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => N345, D => n2252, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => N345, D => n2256, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => N345, D => n2260, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => N345, D => n2264, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N345, D => n2268, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => N345, D => n2272, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N345, D => n2276, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N345, D => n2280, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N345, D => n2284, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => N345, D => n2288, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => N345, D => n2292, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => N345, D => n2296, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => N345, D => n2300, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => N345, D => n2304, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => N345, D => n2308, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => N345, D => n2312, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => N345, D => n2316, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => N345, D => n2320, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => N345, D => n2324, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => N345, D => n2328, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => N345, D => n2332, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => N344, D => n2208, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => N344, D => n2212, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => N344, D => n2216, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => N344, D => n2220, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => N344, D => n2224, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => N344, D => n2228, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => N344, D => n2232, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => N344, D => n2236, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => N344, D => n2240, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => N344, D => n2244, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => N344, D => n2248, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => N344, D => n2252, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => N344, D => n2256, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => N344, D => n2260, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N344, D => n2264, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => N344, D => n2268, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N344, D => n2272, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => N344, D => n2276, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => N344, D => n2280, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N344, D => n2284, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => N344, D => n2288, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => N344, D => n2292, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => N344, D => n2296, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => N344, D => n2300, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => N344, D => n2304, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => N344, D => n2308, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => N344, D => n2312, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => N344, D => n2316, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => N344, D => n2320, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => N344, D => n2324, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => N344, D => n2328, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N344, D => n2332, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => N343, D => n2208, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => N343, D => n2212, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => N343, D => n2216, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => N343, D => n2220, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => N343, D => n2224, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => N343, D => n2228, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => N343, D => n2232, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => N343, D => n2236, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => N343, D => n2240, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => N343, D => n2244, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => N343, D => n2248, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => N343, D => n2252, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => N343, D => n2256, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => N343, D => n2260, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => N343, D => n2264, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N343, D => n2268, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => N343, D => n2272, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N343, D => n2276, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N343, D => n2280, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N343, D => n2284, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => N343, D => n2288, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => N343, D => n2292, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => N343, D => n2296, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => N343, D => n2300, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => N343, D => n2304, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => N343, D => n2308, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => N343, D => n2312, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => N343, D => n2316, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => N343, D => n2320, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => N343, D => n2324, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => N343, D => n2328, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => N343, D => n2332, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => N342, D => n2209, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => N342, D => n2213, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => N342, D => n2217, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => N342, D => n2221, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => N342, D => n2225, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => N342, D => n2229, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => N342, D => n2233, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => N342, D => n2237, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => N342, D => n2241, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => N342, D => n2245, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => N342, D => n2249, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => N342, D => n2253, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => N342, D => n2257, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => N342, D => n2261, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => N342, D => n2265, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N342, D => n2269, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => N342, D => n2273, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N342, D => n2277, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N342, D => n2281, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N342, D => n2285, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => N342, D => n2289, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => N342, D => n2293, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => N342, D => n2297, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => N342, D => n2301, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => N342, D => n2305, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => N342, D => n2309, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => N342, D => n2313, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => N342, D => n2317, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => N342, D => n2321, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => N342, D => n2325, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => N342, D => n2329, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => N342, D => n2333, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => N341, D => n2209, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => N341, D => n2213, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => N341, D => n2217, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => N341, D => n2221, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => N341, D => n2225, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => N341, D => n2229, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => N341, D => n2233, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => N341, D => n2237, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => N341, D => n2241, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => N341, D => n2245, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => N341, D => n2249, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => N341, D => n2253, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => N341, D => n2257, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => N341, D => n2261, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => N341, D => n2265, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N341, D => n2269, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => N341, D => n2273, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N341, D => n2277, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N341, D => n2281, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N341, D => n2285, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => N341, D => n2289, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => N341, D => n2293, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => N341, D => n2297, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => N341, D => n2301, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => N341, D => n2305, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => N341, D => n2309, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => N341, D => n2313, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => N341, D => n2317, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => N341, D => n2321, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => N341, D => n2325, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => N341, D => n2329, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => N341, D => n2333, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => N340, D => n2209, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => N340, D => n2213, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => N340, D => n2217, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => N340, D => n2221, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => N340, D => n2225, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => N340, D => n2229, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => N340, D => n2233, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => N340, D => n2237, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => N340, D => n2241, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => N340, D => n2245, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => N340, D => n2249, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => N340, D => n2253, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => N340, D => n2257, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => N340, D => n2261, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => N340, D => n2265, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N340, D => n2269, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => N340, D => n2273, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N340, D => n2277, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N340, D => n2281, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N340, D => n2285, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => N340, D => n2289, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => N340, D => n2293, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => N340, D => n2297, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => N340, D => n2301, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => N340, D => n2305, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => N340, D => n2309, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => N340, D => n2313, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => N340, D => n2317, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => N340, D => n2321, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => N340, D => n2325, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => N340, D => n2329, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => N340, D => n2333, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => N339, D => n2209, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => N339, D => n2213, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => N339, D => n2217, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => N339, D => n2221, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => N339, D => n2225, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => N339, D => n2229, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => N339, D => n2233, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => N339, D => n2237, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => N339, D => n2241, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => N339, D => n2245, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => N339, D => n2249, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => N339, D => n2253, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => N339, D => n2257, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => N339, D => n2261, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => N339, D => n2265, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N339, D => n2269, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => N339, D => n2273, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N339, D => n2277, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N339, D => n2281, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N339, D => n2285, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => N339, D => n2289, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => N339, D => n2293, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => N339, D => n2297, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => N339, D => n2301, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => N339, D => n2305, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => N339, D => n2309, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => N339, D => n2313, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => N339, D => n2317, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => N339, D => n2321, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => N339, D => n2325, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => N339, D => n2329, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => N339, D => n2333, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => N338, D => n2209, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => N338, D => n2213, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => N338, D => n2217, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => N338, D => n2221, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => N338, D => n2225, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => N338, D => n2229, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => N338, D => n2233, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => N338, D => n2237, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => N338, D => n2241, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => N338, D => n2245, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => N338, D => n2249, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => N338, D => n2253, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => N338, D => n2257, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => N338, D => n2261, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => N338, D => n2265, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N338, D => n2269, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => N338, D => n2273, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N338, D => n2277, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N338, D => n2281, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N338, D => n2285, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => N338, D => n2289, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => N338, D => n2293, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => N338, D => n2297, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => N338, D => n2301, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => N338, D => n2305, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => N338, D => n2309, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => N338, D => n2313, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => N338, D => n2317, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => N338, D => n2321, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => N338, D => n2325, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => N338, D => n2329, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => N338, D => n2333, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => N337, D => n2209, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => N337, D => n2213, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => N337, D => n2217, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => N337, D => n2221, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => N337, D => n2225, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => N337, D => n2229, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => N337, D => n2233, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => N337, D => n2237, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => N337, D => n2241, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => N337, D => n2245, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => N337, D => n2249, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => N337, D => n2253, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => N337, D => n2257, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => N337, D => n2261, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => N337, D => n2265, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N337, D => n2269, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => N337, D => n2273, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N337, D => n2277, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N337, D => n2281, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N337, D => n2285, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => N337, D => n2289, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => N337, D => n2293, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => N337, D => n2297, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => N337, D => n2301, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => N337, D => n2305, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => N337, D => n2309, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => N337, D => n2313, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => N337, D => n2317, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => N337, D => n2321, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => N337, D => n2325, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => N337, D => n2329, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => N337, D => n2333, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => N336, D => n2209, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => N336, D => n2213, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => N336, D => n2217, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => N336, D => n2221, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => N336, D => n2225, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => N336, D => n2229, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => N336, D => n2233, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => N336, D => n2237, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => N336, D => n2241, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => N336, D => n2245, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => N336, D => n2249, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => N336, D => n2253, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => N336, D => n2257, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => N336, D => n2261, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => N336, D => n2265, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N336, D => n2269, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => N336, D => n2273, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N336, D => n2277, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N336, D => n2281, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N336, D => n2285, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => N336, D => n2289, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => N336, D => n2293, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => N336, D => n2297, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => N336, D => n2301, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => N336, D => n2305, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => N336, D => n2309, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => N336, D => n2313, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => N336, D => n2317, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => N336, D => n2321, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => N336, D => n2325, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => N336, D => n2329, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => N336, D => n2333, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => N335, D => n2209, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => N335, D => n2213, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => N335, D => n2217, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => N335, D => n2221, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => N335, D => n2225, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => N335, D => n2229, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => N335, D => n2233, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => N335, D => n2237, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => N335, D => n2241, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => N335, D => n2245, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => N335, D => n2249, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => N335, D => n2253, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => N335, D => n2257, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => N335, D => n2261, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => N335, D => n2265, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N335, D => n2269, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => N335, D => n2273, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N335, D => n2277, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N335, D => n2281, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N335, D => n2285, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => N335, D => n2289, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => N335, D => n2293, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => N335, D => n2297, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => N335, D => n2301, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => N335, D => n2305, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => N335, D => n2309, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => N335, D => n2313, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => N335, D => n2317, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => N335, D => n2321, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => N335, D => n2325, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => N335, D => n2329, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => N335, D => n2333, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => N334, D => n2209, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => N334, D => n2213, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => N334, D => n2217, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => N334, D => n2221, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => N334, D => n2225, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => N334, D => n2229, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => N334, D => n2233, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => N334, D => n2237, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => N334, D => n2241, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => N334, D => n2245, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => N334, D => n2249, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => N334, D => n2253, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => N334, D => n2257, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => N334, D => n2261, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => N334, D => n2265, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N334, D => n2269, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => N334, D => n2273, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N334, D => n2277, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N334, D => n2281, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N334, D => n2285, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => N334, D => n2289, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => N334, D => n2293, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => N334, D => n2297, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => N334, D => n2301, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => N334, D => n2305, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => N334, D => n2309, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => N334, D => n2313, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => N334, D => n2317, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => N334, D => n2321, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => N334, D => n2325, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => N334, D => n2329, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => N334, D => n2333, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => N333, D => n2209, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => N333, D => n2213, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => N333, D => n2217, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => N333, D => n2221, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => N333, D => n2225, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => N333, D => n2229, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => N333, D => n2233, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => N333, D => n2237, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => N333, D => n2241, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => N333, D => n2245, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => N333, D => n2249, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => N333, D => n2253, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => N333, D => n2257, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => N333, D => n2261, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => N333, D => n2265, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N333, D => n2269, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => N333, D => n2273, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N333, D => n2277, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N333, D => n2281, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N333, D => n2285, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => N333, D => n2289, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => N333, D => n2293, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => N333, D => n2297, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => N333, D => n2301, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => N333, D => n2305, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => N333, D => n2309, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => N333, D => n2313, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => N333, D => n2317, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => N333, D => n2321, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => N333, D => n2325, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => N333, D => n2329, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => N333, D => n2333, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => N332, D => n2209, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => N332, D => n2213, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => N332, D => n2217, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => N332, D => n2221, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => N332, D => n2225, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => N332, D => n2229, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => N332, D => n2233, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => N332, D => n2237, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => N332, D => n2241, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => N332, D => n2245, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => N332, D => n2249, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => N332, D => n2253, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => N332, D => n2257, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => N332, D => n2261, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => N332, D => n2265, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N332, D => n2269, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => N332, D => n2273, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N332, D => n2277, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N332, D => n2281, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N332, D => n2285, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => N332, D => n2289, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => N332, D => n2293, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => N332, D => n2297, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => N332, D => n2301, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => N332, D => n2305, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => N332, D => n2309, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => N332, D => n2313, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => N332, D => n2317, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => N332, D => n2321, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => N332, D => n2325, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => N332, D => n2329, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => N332, D => n2333, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => N331, D => n2210, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => N331, D => n2214, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => N331, D => n2218, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => N331, D => n2222, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => N331, D => n2226, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => N331, D => n2230, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => N331, D => n2234, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => N331, D => n2238, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => N331, D => n2242, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => N331, D => n2246, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => N331, D => n2250, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => N331, D => n2254, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => N331, D => n2258, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => N331, D => n2262, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => N331, D => n2266, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N331, D => n2270, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => N331, D => n2274, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N331, D => n2278, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N331, D => n2282, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N331, D => n2286, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => N331, D => n2290, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => N331, D => n2294, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => N331, D => n2298, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => N331, D => n2302, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => N331, D => n2306, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => N331, D => n2310, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => N331, D => n2314, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => N331, D => n2318, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => N331, D => n2322, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => N331, D => n2326, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => N331, D => n2330, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => N331, D => n2334, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => N330, D => n2210, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => N330, D => n2214, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => N330, D => n2218, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => N330, D => n2222, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => N330, D => n2226, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => N330, D => n2230, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => N330, D => n2234, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => N330, D => n2238, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => N330, D => n2242, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => N330, D => n2246, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => N330, D => n2250, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => N330, D => n2254, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => N330, D => n2258, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => N330, D => n2262, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N330, D => n2266, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N330, D => n2270, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => N330, D => n2274, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N330, D => n2278, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N330, D => n2282, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => N330, D => n2286, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => N330, D => n2290, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => N330, D => n2294, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => N330, D => n2298, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => N330, D => n2302, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => N330, D => n2306, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => N330, D => n2310, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => N330, D => n2314, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => N330, D => n2318, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => N330, D => n2322, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => N330, D => n2326, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => N330, D => n2330, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => N330, D => n2334, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => N329, D => n2210, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => N329, D => n2214, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => N329, D => n2218, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => N329, D => n2222, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => N329, D => n2226, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => N329, D => n2230, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => N329, D => n2234, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => N329, D => n2238, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => N329, D => n2242, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => N329, D => n2246, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => N329, D => n2250, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => N329, D => n2254, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => N329, D => n2258, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => N329, D => n2262, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => N329, D => n2266, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N329, D => n2270, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => N329, D => n2274, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N329, D => n2278, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N329, D => n2282, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N329, D => n2286, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => N329, D => n2290, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => N329, D => n2294, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => N329, D => n2298, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => N329, D => n2302, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => N329, D => n2306, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => N329, D => n2310, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => N329, D => n2314, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => N329, D => n2318, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => N329, D => n2322, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => N329, D => n2326, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => N329, D => n2330, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => N329, D => n2334, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => N328, D => n2210, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => N328, D => n2214, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => N328, D => n2218, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => N328, D => n2222, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => N328, D => n2226, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => N328, D => n2230, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => N328, D => n2234, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => N328, D => n2238, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => N328, D => n2242, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => N328, D => n2246, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => N328, D => n2250, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => N328, D => n2254, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => N328, D => n2258, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => N328, D => n2262, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => N328, D => n2266, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N328, D => n2270, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => N328, D => n2274, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N328, D => n2278, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N328, D => n2282, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N328, D => n2286, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => N328, D => n2290, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => N328, D => n2294, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => N328, D => n2298, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => N328, D => n2302, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => N328, D => n2306, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => N328, D => n2310, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => N328, D => n2314, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => N328, D => n2318, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => N328, D => n2322, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => N328, D => n2326, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => N328, D => n2330, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => N328, D => n2334, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => N327, D => n2210, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => N327, D => n2214, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => N327, D => n2218, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => N327, D => n2222, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => N327, D => n2226, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => N327, D => n2230, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => N327, D => n2234, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => N327, D => n2238, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => N327, D => n2242, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => N327, D => n2246, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => N327, D => n2250, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => N327, D => n2254, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => N327, D => n2258, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => N327, D => n2262, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => N327, D => n2266, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N327, D => n2270, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => N327, D => n2274, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N327, D => n2278, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N327, D => n2282, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N327, D => n2286, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => N327, D => n2290, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => N327, D => n2294, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => N327, D => n2298, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => N327, D => n2302, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => N327, D => n2306, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => N327, D => n2310, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => N327, D => n2314, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => N327, D => n2318, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => N327, D => n2322, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => N327, D => n2326, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => N327, D => n2330, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => N327, D => n2334, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => N326, D => n2210, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => N326, D => n2214, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => N326, D => n2218, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => N326, D => n2222, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => N326, D => n2226, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => N326, D => n2230, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => N326, D => n2234, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => N326, D => n2238, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => N326, D => n2242, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => N326, D => n2246, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => N326, D => n2250, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => N326, D => n2254, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => N326, D => n2258, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => N326, D => n2262, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => N326, D => n2266, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N326, D => n2270, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => N326, D => n2274, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N326, D => n2278, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N326, D => n2282, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N326, D => n2286, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => N326, D => n2290, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => N326, D => n2294, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => N326, D => n2298, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => N326, D => n2302, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => N326, D => n2306, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => N326, D => n2310, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => N326, D => n2314, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => N326, D => n2318, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => N326, D => n2322, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => N326, D => n2326, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => N326, D => n2330, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => N326, D => n2334, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => N325, D => n2210, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => N325, D => n2214, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => N325, D => n2218, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => N325, D => n2222, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => N325, D => n2226, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => N325, D => n2230, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => N325, D => n2234, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => N325, D => n2238, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => N325, D => n2242, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => N325, D => n2246, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => N325, D => n2250, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => N325, D => n2254, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => N325, D => n2258, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => N325, D => n2262, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => N325, D => n2266, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N325, D => n2270, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => N325, D => n2274, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N325, D => n2278, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N325, D => n2282, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N325, D => n2286, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => N325, D => n2290, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => N325, D => n2294, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => N325, D => n2298, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => N325, D => n2302, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => N325, D => n2306, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => N325, D => n2310, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => N325, D => n2314, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => N325, D => n2318, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => N325, D => n2322, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => N325, D => n2326, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => N325, D => n2330, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => N325, D => n2334, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => N324, D => n2210, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => N324, D => n2214, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => N324, D => n2218, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => N324, D => n2222, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => N324, D => n2226, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => N324, D => n2230, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => N324, D => n2234, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => N324, D => n2238, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => N324, D => n2242, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => N324, D => n2246, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => N324, D => n2250, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => N324, D => n2254, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => N324, D => n2258, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => N324, D => n2262, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => N324, D => n2266, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N324, D => n2270, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => N324, D => n2274, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N324, D => n2278, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N324, D => n2282, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N324, D => n2286, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => N324, D => n2290, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => N324, D => n2294, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => N324, D => n2298, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => N324, D => n2302, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => N324, D => n2306, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => N324, D => n2310, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => N324, D => n2314, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => N324, D => n2318, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => N324, D => n2322, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => N324, D => n2326, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => N324, D => n2330, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => N324, D => n2334, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => N323, D => n2210, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => N323, D => n2214, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => N323, D => n2218, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => N323, D => n2222, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => N323, D => n2226, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => N323, D => n2230, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => N323, D => n2234, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => N323, D => n2238, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => N323, D => n2242, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => N323, D => n2246, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => N323, D => n2250, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => N323, D => n2254, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => N323, D => n2258, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => N323, D => n2262, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => N323, D => n2266, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N323, D => n2270, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => N323, D => n2274, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N323, D => n2278, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N323, D => n2282, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N323, D => n2286, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => N323, D => n2290, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => N323, D => n2294, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => N323, D => n2298, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => N323, D => n2302, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => N323, D => n2306, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => N323, D => n2310, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => N323, D => n2314, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => N323, D => n2318, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => N323, D => n2322, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => N323, D => n2326, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => N323, D => n2330, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => N323, D => n2334, Q => 
                           REGISTERS_31_0_port);
   OUT2_reg_31_inst : DLH_X1 port map( G => CLK, D => N322, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => CLK, D => N321, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => CLK, D => N320, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => CLK, D => N319, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => CLK, D => N318, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => CLK, D => N317, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => CLK, D => N316, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => CLK, D => N315, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => CLK, D => N314, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => CLK, D => N313, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => CLK, D => N312, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => CLK, D => N311, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => CLK, D => N310, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => CLK, D => N309, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => CLK, D => N308, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => CLK, D => N307, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => CLK, D => N306, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => CLK, D => N305, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => CLK, D => N304, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => CLK, D => N303, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => CLK, D => N302, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => CLK, D => N301, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => CLK, D => N300, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => CLK, D => N299, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => CLK, D => N298, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => CLK, D => N297, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => CLK, D => N296, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => CLK, D => N295, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => CLK, D => N294, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => CLK, D => N293, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => CLK, D => N292, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => CLK, D => N291, Q => OUT2(0));
   U3 : OAI21_X2 port map( B1 => n890, B2 => n891, A => n2207, ZN => N353);
   U4 : OAI21_X2 port map( B1 => n890, B2 => n893, A => n2207, ZN => N352);
   U5 : OAI21_X2 port map( B1 => n890, B2 => n894, A => n2207, ZN => N351);
   U6 : OAI21_X2 port map( B1 => n890, B2 => n895, A => n2207, ZN => N350);
   U7 : OAI21_X2 port map( B1 => n890, B2 => n896, A => n2207, ZN => N349);
   U8 : OAI21_X2 port map( B1 => n890, B2 => n897, A => n2207, ZN => N348);
   U9 : OAI21_X2 port map( B1 => n890, B2 => n898, A => n2207, ZN => N347);
   U10 : OAI21_X2 port map( B1 => n900, B2 => n901, A => n2206, ZN => N346);
   U11 : OAI21_X2 port map( B1 => n891, B2 => n900, A => n2206, ZN => N345);
   U12 : OAI21_X2 port map( B1 => n893, B2 => n900, A => n2206, ZN => N344);
   U13 : OAI21_X2 port map( B1 => n894, B2 => n900, A => n2206, ZN => N343);
   U14 : OAI21_X2 port map( B1 => n895, B2 => n900, A => n2206, ZN => N342);
   U15 : OAI21_X2 port map( B1 => n896, B2 => n900, A => n2206, ZN => N341);
   U16 : OAI21_X2 port map( B1 => n897, B2 => n900, A => n2206, ZN => N340);
   U17 : OAI21_X2 port map( B1 => n898, B2 => n900, A => n2206, ZN => N339);
   U18 : OAI21_X2 port map( B1 => n901, B2 => n902, A => n2206, ZN => N338);
   U19 : OAI21_X2 port map( B1 => n891, B2 => n902, A => n2206, ZN => N337);
   U20 : OAI21_X2 port map( B1 => n893, B2 => n902, A => n2206, ZN => N336);
   U21 : OAI21_X2 port map( B1 => n894, B2 => n902, A => n2206, ZN => N335);
   U22 : OAI21_X2 port map( B1 => n895, B2 => n902, A => n2205, ZN => N334);
   U23 : OAI21_X2 port map( B1 => n896, B2 => n902, A => n2205, ZN => N333);
   U24 : OAI21_X2 port map( B1 => n897, B2 => n902, A => n2205, ZN => N332);
   U25 : OAI21_X2 port map( B1 => n898, B2 => n902, A => n2205, ZN => N331);
   U26 : OAI21_X2 port map( B1 => n901, B2 => n903, A => n2205, ZN => N330);
   U27 : OAI21_X2 port map( B1 => n891, B2 => n903, A => n2205, ZN => N329);
   U28 : OAI21_X2 port map( B1 => n893, B2 => n903, A => n2205, ZN => N328);
   U29 : OAI21_X2 port map( B1 => n894, B2 => n903, A => n2205, ZN => N327);
   U30 : OAI21_X2 port map( B1 => n895, B2 => n903, A => n2205, ZN => N326);
   U31 : OAI21_X2 port map( B1 => n896, B2 => n903, A => n2205, ZN => N325);
   U32 : OAI21_X2 port map( B1 => n897, B2 => n903, A => n2205, ZN => N324);
   U33 : OAI21_X2 port map( B1 => n898, B2 => n903, A => n2205, ZN => N323);
   U2043 : NAND3_X1 port map( A1 => n3208, A2 => n3207, A3 => n899, ZN => n890)
                           ;
   U2044 : NAND3_X1 port map( A1 => n899, A2 => n3207, A3 => ADD_WR(3), ZN => 
                           n900);
   U2045 : NAND3_X1 port map( A1 => n899, A2 => n3208, A3 => ADD_WR(4), ZN => 
                           n902);
   U2046 : NAND3_X1 port map( A1 => n3210, A2 => n3209, A3 => n3211, ZN => n901
                           );
   U2047 : NAND3_X1 port map( A1 => n3210, A2 => n3209, A3 => ADD_WR(0), ZN => 
                           n891);
   U2048 : NAND3_X1 port map( A1 => n3211, A2 => n3209, A3 => ADD_WR(1), ZN => 
                           n893);
   U2049 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n3209, A3 => ADD_WR(1), ZN
                           => n894);
   U2050 : NAND3_X1 port map( A1 => n3211, A2 => n3210, A3 => ADD_WR(2), ZN => 
                           n895);
   U2051 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n3210, A3 => ADD_WR(2), ZN
                           => n896);
   U2052 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n3211, A3 => ADD_WR(2), ZN
                           => n897);
   U2053 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n899, A3 => ADD_WR(4), ZN 
                           => n903);
   U2054 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n898);
   U34 : NOR2_X1 port map( A1 => n3216, A2 => n3217, ZN => n1408);
   U35 : NOR2_X1 port map( A1 => n3212, A2 => n3213, ZN => n1923);
   U36 : NOR2_X1 port map( A1 => n3212, A2 => ADD_RD1(3), ZN => n1933);
   U37 : BUF_X1 port map( A => n2336, Z => n2340);
   U38 : BUF_X1 port map( A => n1934, Z => n2122);
   U39 : BUF_X1 port map( A => n1425, Z => n2072);
   U40 : BUF_X1 port map( A => n1436, Z => n2028);
   U41 : BUF_X1 port map( A => n1434, Z => n2036);
   U42 : BUF_X1 port map( A => n919, Z => n2164);
   U43 : BUF_X1 port map( A => n910, Z => n2200);
   U44 : BUF_X1 port map( A => n915, Z => n2180);
   U45 : BUF_X1 port map( A => n921, Z => n2156);
   U46 : BUF_X1 port map( A => n1430, Z => n2052);
   U47 : BUF_X1 port map( A => n914, Z => n2184);
   U48 : BUF_X1 port map( A => n916, Z => n2176);
   U49 : BUF_X1 port map( A => n950, Z => n2076);
   U50 : BUF_X1 port map( A => n949, Z => n2080);
   U51 : BUF_X1 port map( A => n1429, Z => n2056);
   U52 : BUF_X1 port map( A => n1431, Z => n2048);
   U53 : BUF_X1 port map( A => n1465, Z => n1948);
   U54 : BUF_X1 port map( A => n1464, Z => n1952);
   U55 : BUF_X1 port map( A => N128, Z => n2335);
   U56 : BUF_X1 port map( A => N129, Z => n2331);
   U57 : BUF_X1 port map( A => N130, Z => n2327);
   U58 : BUF_X1 port map( A => N131, Z => n2323);
   U59 : BUF_X1 port map( A => N132, Z => n2319);
   U60 : BUF_X1 port map( A => N133, Z => n2315);
   U61 : BUF_X1 port map( A => N134, Z => n2311);
   U62 : BUF_X1 port map( A => N135, Z => n2307);
   U63 : BUF_X1 port map( A => N136, Z => n2303);
   U64 : BUF_X1 port map( A => N137, Z => n2299);
   U65 : BUF_X1 port map( A => N138, Z => n2295);
   U66 : BUF_X1 port map( A => N139, Z => n2291);
   U67 : BUF_X1 port map( A => N140, Z => n2287);
   U68 : BUF_X1 port map( A => N141, Z => n2283);
   U69 : BUF_X1 port map( A => N142, Z => n2279);
   U70 : BUF_X1 port map( A => N143, Z => n2275);
   U71 : BUF_X1 port map( A => N144, Z => n2271);
   U72 : BUF_X1 port map( A => N145, Z => n2267);
   U73 : BUF_X1 port map( A => N146, Z => n2263);
   U74 : BUF_X1 port map( A => N147, Z => n2259);
   U75 : BUF_X1 port map( A => N148, Z => n2255);
   U76 : BUF_X1 port map( A => N149, Z => n2251);
   U77 : BUF_X1 port map( A => N150, Z => n2247);
   U78 : BUF_X1 port map( A => N151, Z => n2243);
   U79 : BUF_X1 port map( A => N159, Z => n2211);
   U80 : BUF_X1 port map( A => N152, Z => n2239);
   U81 : BUF_X1 port map( A => N153, Z => n2235);
   U82 : BUF_X1 port map( A => N154, Z => n2231);
   U83 : BUF_X1 port map( A => N155, Z => n2227);
   U84 : BUF_X1 port map( A => N156, Z => n2223);
   U85 : BUF_X1 port map( A => N157, Z => n2219);
   U86 : BUF_X1 port map( A => N158, Z => n2215);
   U87 : BUF_X1 port map( A => n935, Z => n2135);
   U88 : BUF_X1 port map( A => n1940, Z => n2142);
   U89 : BUF_X1 port map( A => n1941, Z => n2138);
   U90 : BUF_X1 port map( A => n1939, Z => n2126);
   U91 : BUF_X1 port map( A => n1935, Z => n2010);
   U92 : BUF_X1 port map( A => n1936, Z => n2014);
   U93 : BUF_X1 port map( A => n1937, Z => n1994);
   U94 : BUF_X1 port map( A => n1938, Z => n1998);
   U95 : BUF_X1 port map( A => n1427, Z => n2064);
   U96 : BUF_X1 port map( A => n1426, Z => n2068);
   U97 : BUF_X1 port map( A => n1428, Z => n2060);
   U98 : BUF_X1 port map( A => n1433, Z => n2040);
   U99 : BUF_X1 port map( A => n1432, Z => n2044);
   U100 : BUF_X1 port map( A => n1435, Z => n2032);
   U101 : BUF_X1 port map( A => n1463, Z => n1956);
   U102 : BUF_X1 port map( A => n944, Z => n2100);
   U103 : BUF_X1 port map( A => n945, Z => n2096);
   U104 : BUF_X1 port map( A => n1459, Z => n1972);
   U105 : BUF_X1 port map( A => n1457, Z => n1980);
   U106 : BUF_X1 port map( A => n1461, Z => n1964);
   U107 : BUF_X1 port map( A => n1460, Z => n1968);
   U108 : BUF_X1 port map( A => n912, Z => n2192);
   U109 : BUF_X1 port map( A => n911, Z => n2196);
   U110 : BUF_X1 port map( A => n913, Z => n2188);
   U111 : BUF_X1 port map( A => n918, Z => n2168);
   U112 : BUF_X1 port map( A => n917, Z => n2172);
   U113 : BUF_X1 port map( A => n920, Z => n2160);
   U114 : BUF_X1 port map( A => n942, Z => n2108);
   U115 : BUF_X1 port map( A => n946, Z => n2092);
   U116 : BUF_X1 port map( A => n948, Z => n2084);
   U117 : BUF_X1 port map( A => n943, Z => n2104);
   U118 : BUF_X1 port map( A => n947, Z => n2088);
   U119 : BUF_X1 port map( A => n926, Z => n2152);
   U120 : BUF_X1 port map( A => n927, Z => n2148);
   U121 : BUF_X1 port map( A => n1458, Z => n1976);
   U122 : BUF_X1 port map( A => n1462, Z => n1960);
   U123 : BUF_X1 port map( A => n1442, Z => n2020);
   U124 : BUF_X1 port map( A => n1441, Z => n2024);
   U125 : BUF_X1 port map( A => n892, Z => n2204);
   U126 : BUF_X1 port map( A => n1451, Z => n2003);
   U127 : BUF_X1 port map( A => n1455, Z => n1991);
   U128 : BUF_X1 port map( A => n1456, Z => n1987);
   U129 : BUF_X1 port map( A => n936, Z => n2131);
   U130 : BUF_X1 port map( A => n941, Z => n2115);
   U131 : BUF_X1 port map( A => n940, Z => n2119);
   U132 : BUF_X1 port map( A => n1446, Z => n2019);
   U133 : BUF_X1 port map( A => n931, Z => n2147);
   U134 : BUF_X1 port map( A => n1450, Z => n2007);
   U135 : INV_X1 port map( A => n2340, ZN => n2337);
   U136 : INV_X1 port map( A => n2340, ZN => n2338);
   U137 : INV_X1 port map( A => n2340, ZN => n2339);
   U138 : BUF_X1 port map( A => n2180, Z => n2181);
   U139 : BUF_X1 port map( A => n2156, Z => n2157);
   U140 : BUF_X1 port map( A => n2076, Z => n2077);
   U141 : BUF_X1 port map( A => n2180, Z => n2182);
   U142 : BUF_X1 port map( A => n2156, Z => n2158);
   U143 : BUF_X1 port map( A => n2076, Z => n2078);
   U144 : BUF_X1 port map( A => n2184, Z => n2185);
   U145 : BUF_X1 port map( A => n2080, Z => n2081);
   U146 : BUF_X1 port map( A => n2184, Z => n2186);
   U147 : BUF_X1 port map( A => n2080, Z => n2082);
   U148 : BUF_X1 port map( A => n2200, Z => n2201);
   U149 : BUF_X1 port map( A => n2176, Z => n2177);
   U150 : BUF_X1 port map( A => n2164, Z => n2165);
   U151 : BUF_X1 port map( A => n2200, Z => n2202);
   U152 : BUF_X1 port map( A => n2176, Z => n2178);
   U153 : BUF_X1 port map( A => n2164, Z => n2166);
   U154 : BUF_X1 port map( A => n2052, Z => n2053);
   U155 : BUF_X1 port map( A => n2028, Z => n2029);
   U156 : BUF_X1 port map( A => n1948, Z => n1949);
   U157 : BUF_X1 port map( A => n2052, Z => n2054);
   U158 : BUF_X1 port map( A => n2028, Z => n2030);
   U159 : BUF_X1 port map( A => n1948, Z => n1950);
   U160 : BUF_X1 port map( A => n2056, Z => n2057);
   U161 : BUF_X1 port map( A => n1952, Z => n1953);
   U162 : BUF_X1 port map( A => n2056, Z => n2058);
   U163 : BUF_X1 port map( A => n1952, Z => n1954);
   U164 : BUF_X1 port map( A => n2072, Z => n2073);
   U165 : BUF_X1 port map( A => n2048, Z => n2049);
   U166 : BUF_X1 port map( A => n2036, Z => n2037);
   U167 : BUF_X1 port map( A => n2072, Z => n2074);
   U168 : BUF_X1 port map( A => n2048, Z => n2050);
   U169 : BUF_X1 port map( A => n2036, Z => n2038);
   U170 : INV_X1 port map( A => n2122, ZN => n2120);
   U171 : INV_X1 port map( A => n2122, ZN => n2121);
   U172 : BUF_X1 port map( A => n2180, Z => n2183);
   U173 : BUF_X1 port map( A => n2156, Z => n2159);
   U174 : BUF_X1 port map( A => n2076, Z => n2079);
   U175 : BUF_X1 port map( A => n2184, Z => n2187);
   U176 : BUF_X1 port map( A => n2080, Z => n2083);
   U177 : BUF_X1 port map( A => n2200, Z => n2203);
   U178 : BUF_X1 port map( A => n2176, Z => n2179);
   U179 : BUF_X1 port map( A => n2164, Z => n2167);
   U180 : BUF_X1 port map( A => n2052, Z => n2055);
   U181 : BUF_X1 port map( A => n2028, Z => n2031);
   U182 : BUF_X1 port map( A => n1948, Z => n1951);
   U183 : BUF_X1 port map( A => n2056, Z => n2059);
   U184 : BUF_X1 port map( A => n1952, Z => n1955);
   U185 : BUF_X1 port map( A => n2072, Z => n2075);
   U186 : BUF_X1 port map( A => n2048, Z => n2051);
   U187 : BUF_X1 port map( A => n2036, Z => n2039);
   U188 : BUF_X1 port map( A => n2335, Z => n2333);
   U189 : BUF_X1 port map( A => n2331, Z => n2329);
   U190 : BUF_X1 port map( A => n2327, Z => n2325);
   U191 : BUF_X1 port map( A => n2323, Z => n2321);
   U192 : BUF_X1 port map( A => n2319, Z => n2317);
   U193 : BUF_X1 port map( A => n2315, Z => n2313);
   U194 : BUF_X1 port map( A => n2311, Z => n2309);
   U195 : BUF_X1 port map( A => n2307, Z => n2305);
   U196 : BUF_X1 port map( A => n2303, Z => n2301);
   U197 : BUF_X1 port map( A => n2299, Z => n2297);
   U198 : BUF_X1 port map( A => n2295, Z => n2293);
   U199 : BUF_X1 port map( A => n2291, Z => n2289);
   U200 : BUF_X1 port map( A => n2287, Z => n2285);
   U201 : BUF_X1 port map( A => n2283, Z => n2281);
   U202 : BUF_X1 port map( A => n2279, Z => n2277);
   U203 : BUF_X1 port map( A => n2275, Z => n2273);
   U204 : BUF_X1 port map( A => n2271, Z => n2269);
   U205 : BUF_X1 port map( A => n2267, Z => n2265);
   U206 : BUF_X1 port map( A => n2263, Z => n2261);
   U207 : BUF_X1 port map( A => n2259, Z => n2257);
   U208 : BUF_X1 port map( A => n2255, Z => n2253);
   U209 : BUF_X1 port map( A => n2251, Z => n2249);
   U210 : BUF_X1 port map( A => n2247, Z => n2245);
   U211 : BUF_X1 port map( A => n2243, Z => n2241);
   U212 : BUF_X1 port map( A => n2239, Z => n2237);
   U213 : BUF_X1 port map( A => n2235, Z => n2233);
   U214 : BUF_X1 port map( A => n2231, Z => n2229);
   U215 : BUF_X1 port map( A => n2227, Z => n2225);
   U216 : BUF_X1 port map( A => n2223, Z => n2221);
   U217 : BUF_X1 port map( A => n2219, Z => n2217);
   U218 : BUF_X1 port map( A => n2215, Z => n2213);
   U219 : BUF_X1 port map( A => n2335, Z => n2332);
   U220 : BUF_X1 port map( A => n2331, Z => n2328);
   U221 : BUF_X1 port map( A => n2327, Z => n2324);
   U222 : BUF_X1 port map( A => n2323, Z => n2320);
   U223 : BUF_X1 port map( A => n2319, Z => n2316);
   U224 : BUF_X1 port map( A => n2315, Z => n2312);
   U225 : BUF_X1 port map( A => n2311, Z => n2308);
   U226 : BUF_X1 port map( A => n2307, Z => n2304);
   U227 : BUF_X1 port map( A => n2303, Z => n2300);
   U228 : BUF_X1 port map( A => n2299, Z => n2296);
   U229 : BUF_X1 port map( A => n2295, Z => n2292);
   U230 : BUF_X1 port map( A => n2291, Z => n2288);
   U231 : BUF_X1 port map( A => n2287, Z => n2284);
   U232 : BUF_X1 port map( A => n2283, Z => n2280);
   U233 : BUF_X1 port map( A => n2279, Z => n2276);
   U234 : BUF_X1 port map( A => n2275, Z => n2272);
   U235 : BUF_X1 port map( A => n2271, Z => n2268);
   U236 : BUF_X1 port map( A => n2267, Z => n2264);
   U237 : BUF_X1 port map( A => n2263, Z => n2260);
   U238 : BUF_X1 port map( A => n2259, Z => n2256);
   U239 : BUF_X1 port map( A => n2255, Z => n2252);
   U240 : BUF_X1 port map( A => n2251, Z => n2248);
   U241 : BUF_X1 port map( A => n2247, Z => n2244);
   U242 : BUF_X1 port map( A => n2243, Z => n2240);
   U243 : BUF_X1 port map( A => n2239, Z => n2236);
   U244 : BUF_X1 port map( A => n2235, Z => n2232);
   U245 : BUF_X1 port map( A => n2231, Z => n2228);
   U246 : BUF_X1 port map( A => n2227, Z => n2224);
   U247 : BUF_X1 port map( A => n2223, Z => n2220);
   U248 : BUF_X1 port map( A => n2219, Z => n2216);
   U249 : BUF_X1 port map( A => n2215, Z => n2212);
   U250 : BUF_X1 port map( A => n2211, Z => n2209);
   U251 : BUF_X1 port map( A => n2211, Z => n2208);
   U252 : BUF_X1 port map( A => n2335, Z => n2334);
   U253 : BUF_X1 port map( A => n2331, Z => n2330);
   U254 : BUF_X1 port map( A => n2327, Z => n2326);
   U255 : BUF_X1 port map( A => n2323, Z => n2322);
   U256 : BUF_X1 port map( A => n2319, Z => n2318);
   U257 : BUF_X1 port map( A => n2315, Z => n2314);
   U258 : BUF_X1 port map( A => n2311, Z => n2310);
   U259 : BUF_X1 port map( A => n2307, Z => n2306);
   U260 : BUF_X1 port map( A => n2303, Z => n2302);
   U261 : BUF_X1 port map( A => n2299, Z => n2298);
   U262 : BUF_X1 port map( A => n2295, Z => n2294);
   U263 : BUF_X1 port map( A => n2291, Z => n2290);
   U264 : BUF_X1 port map( A => n2287, Z => n2286);
   U265 : BUF_X1 port map( A => n2283, Z => n2282);
   U266 : BUF_X1 port map( A => n2279, Z => n2278);
   U267 : BUF_X1 port map( A => n2275, Z => n2274);
   U268 : BUF_X1 port map( A => n2271, Z => n2270);
   U269 : BUF_X1 port map( A => n2267, Z => n2266);
   U270 : BUF_X1 port map( A => n2263, Z => n2262);
   U271 : BUF_X1 port map( A => n2259, Z => n2258);
   U272 : BUF_X1 port map( A => n2255, Z => n2254);
   U273 : BUF_X1 port map( A => n2251, Z => n2250);
   U274 : BUF_X1 port map( A => n2247, Z => n2246);
   U275 : BUF_X1 port map( A => n2243, Z => n2242);
   U276 : BUF_X1 port map( A => n2239, Z => n2238);
   U277 : BUF_X1 port map( A => n2235, Z => n2234);
   U278 : BUF_X1 port map( A => n2231, Z => n2230);
   U279 : BUF_X1 port map( A => n2227, Z => n2226);
   U280 : BUF_X1 port map( A => n2223, Z => n2222);
   U281 : BUF_X1 port map( A => n2219, Z => n2218);
   U282 : BUF_X1 port map( A => n2215, Z => n2214);
   U283 : BUF_X1 port map( A => n2211, Z => n2210);
   U284 : NAND2_X1 port map( A1 => n2130, A2 => n1408, ZN => n910);
   U285 : NAND2_X1 port map( A1 => n2134, A2 => n1408, ZN => n915);
   U286 : NAND2_X1 port map( A1 => n2123, A2 => n1408, ZN => n914);
   U287 : NAND2_X1 port map( A1 => n2127, A2 => n1408, ZN => n916);
   U288 : NAND2_X1 port map( A1 => n2114, A2 => n1408, ZN => n921);
   U289 : NAND2_X1 port map( A1 => n1408, A2 => n2118, ZN => n919);
   U290 : NAND2_X1 port map( A1 => n2139, A2 => n1408, ZN => n950);
   U291 : NAND2_X1 port map( A1 => n2143, A2 => n1408, ZN => n949);
   U292 : NAND2_X1 port map( A1 => n2000, A2 => n1923, ZN => n1425);
   U293 : NAND2_X1 port map( A1 => n2006, A2 => n1923, ZN => n1430);
   U294 : NAND2_X1 port map( A1 => n1995, A2 => n1923, ZN => n1429);
   U295 : NAND2_X1 port map( A1 => n1999, A2 => n1923, ZN => n1431);
   U296 : NAND2_X1 port map( A1 => n1984, A2 => n1923, ZN => n1436);
   U297 : NAND2_X1 port map( A1 => n1923, A2 => n1988, ZN => n1434);
   U298 : NAND2_X1 port map( A1 => n2011, A2 => n1923, ZN => n1465);
   U299 : NAND2_X1 port map( A1 => n2015, A2 => n1923, ZN => n1464);
   U300 : BUF_X1 port map( A => RESET, Z => n2336);
   U301 : BUF_X1 port map( A => n2135, Z => n2132);
   U302 : BUF_X1 port map( A => n2135, Z => n2133);
   U303 : BUF_X1 port map( A => n2152, Z => n2153);
   U304 : BUF_X1 port map( A => n2152, Z => n2154);
   U305 : BUF_X1 port map( A => n2192, Z => n2193);
   U306 : BUF_X1 port map( A => n2168, Z => n2169);
   U307 : BUF_X1 port map( A => n2100, Z => n2101);
   U308 : BUF_X1 port map( A => n2088, Z => n2089);
   U309 : BUF_X1 port map( A => n2192, Z => n2194);
   U310 : BUF_X1 port map( A => n2168, Z => n2170);
   U311 : BUF_X1 port map( A => n2100, Z => n2102);
   U312 : BUF_X1 port map( A => n2088, Z => n2090);
   U313 : BUF_X1 port map( A => n2196, Z => n2197);
   U314 : BUF_X1 port map( A => n2172, Z => n2173);
   U315 : BUF_X1 port map( A => n2160, Z => n2161);
   U316 : BUF_X1 port map( A => n2104, Z => n2105);
   U317 : BUF_X1 port map( A => n2092, Z => n2093);
   U318 : BUF_X1 port map( A => n2196, Z => n2198);
   U319 : BUF_X1 port map( A => n2172, Z => n2174);
   U320 : BUF_X1 port map( A => n2160, Z => n2162);
   U321 : BUF_X1 port map( A => n2104, Z => n2106);
   U322 : BUF_X1 port map( A => n2092, Z => n2094);
   U323 : BUF_X1 port map( A => n2188, Z => n2189);
   U324 : BUF_X1 port map( A => n2108, Z => n2109);
   U325 : BUF_X1 port map( A => n2096, Z => n2097);
   U326 : BUF_X1 port map( A => n2084, Z => n2085);
   U327 : BUF_X1 port map( A => n2188, Z => n2190);
   U328 : BUF_X1 port map( A => n2108, Z => n2110);
   U329 : BUF_X1 port map( A => n2096, Z => n2098);
   U330 : BUF_X1 port map( A => n2084, Z => n2086);
   U331 : BUF_X1 port map( A => n2020, Z => n2021);
   U332 : BUF_X1 port map( A => n2020, Z => n2022);
   U333 : BUF_X1 port map( A => n2204, Z => n2205);
   U334 : BUF_X1 port map( A => n2204, Z => n2206);
   U335 : BUF_X1 port map( A => n2135, Z => n2134);
   U336 : BUF_X1 port map( A => n3205, Z => n1942);
   U337 : BUF_X1 port map( A => n3205, Z => n1943);
   U338 : BUF_X1 port map( A => n3206, Z => n1945);
   U339 : BUF_X1 port map( A => n3206, Z => n1946);
   U340 : BUF_X1 port map( A => n2024, Z => n2025);
   U341 : BUF_X1 port map( A => n2024, Z => n2026);
   U342 : INV_X1 port map( A => n2142, ZN => n2140);
   U343 : INV_X1 port map( A => n2126, ZN => n2124);
   U344 : BUF_X1 port map( A => n2064, Z => n2065);
   U345 : BUF_X1 port map( A => n2040, Z => n2041);
   U346 : BUF_X1 port map( A => n1972, Z => n1973);
   U347 : BUF_X1 port map( A => n1960, Z => n1961);
   U348 : BUF_X1 port map( A => n2064, Z => n2066);
   U349 : BUF_X1 port map( A => n2040, Z => n2042);
   U350 : BUF_X1 port map( A => n1972, Z => n1974);
   U351 : BUF_X1 port map( A => n1960, Z => n1962);
   U352 : BUF_X1 port map( A => n2068, Z => n2069);
   U353 : BUF_X1 port map( A => n2044, Z => n2045);
   U354 : BUF_X1 port map( A => n2032, Z => n2033);
   U355 : BUF_X1 port map( A => n1976, Z => n1977);
   U356 : BUF_X1 port map( A => n1964, Z => n1965);
   U357 : BUF_X1 port map( A => n2068, Z => n2070);
   U358 : BUF_X1 port map( A => n2044, Z => n2046);
   U359 : BUF_X1 port map( A => n2032, Z => n2034);
   U360 : BUF_X1 port map( A => n1976, Z => n1978);
   U361 : BUF_X1 port map( A => n1964, Z => n1966);
   U362 : BUF_X1 port map( A => n2148, Z => n2149);
   U363 : BUF_X1 port map( A => n2148, Z => n2150);
   U364 : BUF_X1 port map( A => n2060, Z => n2061);
   U365 : BUF_X1 port map( A => n1980, Z => n1981);
   U366 : BUF_X1 port map( A => n1968, Z => n1969);
   U367 : BUF_X1 port map( A => n1956, Z => n1957);
   U368 : BUF_X1 port map( A => n2060, Z => n2062);
   U369 : BUF_X1 port map( A => n1980, Z => n1982);
   U370 : BUF_X1 port map( A => n1968, Z => n1970);
   U371 : BUF_X1 port map( A => n1956, Z => n1958);
   U372 : INV_X1 port map( A => n2010, ZN => n2008);
   U373 : INV_X1 port map( A => n1994, ZN => n1992);
   U374 : INV_X1 port map( A => n2010, ZN => n2009);
   U375 : INV_X1 port map( A => n1994, ZN => n1993);
   U376 : INV_X1 port map( A => n2014, ZN => n2012);
   U377 : INV_X1 port map( A => n1998, ZN => n1996);
   U378 : INV_X1 port map( A => n2138, ZN => n2136);
   U379 : INV_X1 port map( A => n2138, ZN => n2137);
   U380 : BUF_X1 port map( A => n2152, Z => n2155);
   U381 : BUF_X1 port map( A => n2192, Z => n2195);
   U382 : BUF_X1 port map( A => n2168, Z => n2171);
   U383 : BUF_X1 port map( A => n2100, Z => n2103);
   U384 : BUF_X1 port map( A => n2088, Z => n2091);
   U385 : BUF_X1 port map( A => n2196, Z => n2199);
   U386 : BUF_X1 port map( A => n2172, Z => n2175);
   U387 : BUF_X1 port map( A => n2160, Z => n2163);
   U388 : BUF_X1 port map( A => n2104, Z => n2107);
   U389 : BUF_X1 port map( A => n2092, Z => n2095);
   U390 : BUF_X1 port map( A => n2188, Z => n2191);
   U391 : BUF_X1 port map( A => n2108, Z => n2111);
   U392 : BUF_X1 port map( A => n2096, Z => n2099);
   U393 : BUF_X1 port map( A => n2084, Z => n2087);
   U394 : BUF_X1 port map( A => n2020, Z => n2023);
   U395 : BUF_X1 port map( A => n3205, Z => n1944);
   U396 : BUF_X1 port map( A => n3206, Z => n1947);
   U397 : BUF_X1 port map( A => n2024, Z => n2027);
   U398 : BUF_X1 port map( A => n2064, Z => n2067);
   U399 : BUF_X1 port map( A => n2040, Z => n2043);
   U400 : BUF_X1 port map( A => n1972, Z => n1975);
   U401 : BUF_X1 port map( A => n1960, Z => n1963);
   U402 : BUF_X1 port map( A => n2068, Z => n2071);
   U403 : BUF_X1 port map( A => n2044, Z => n2047);
   U404 : BUF_X1 port map( A => n2032, Z => n2035);
   U405 : BUF_X1 port map( A => n1976, Z => n1979);
   U406 : BUF_X1 port map( A => n1964, Z => n1967);
   U407 : BUF_X1 port map( A => n2148, Z => n2151);
   U408 : BUF_X1 port map( A => n2060, Z => n2063);
   U409 : BUF_X1 port map( A => n1980, Z => n1983);
   U410 : BUF_X1 port map( A => n1968, Z => n1971);
   U411 : BUF_X1 port map( A => n1956, Z => n1959);
   U412 : INV_X1 port map( A => n2142, ZN => n2141);
   U413 : INV_X1 port map( A => n2126, ZN => n2125);
   U414 : BUF_X1 port map( A => n2204, Z => n2207);
   U415 : INV_X1 port map( A => n2014, ZN => n2013);
   U416 : INV_X1 port map( A => n1998, ZN => n1997);
   U417 : BUF_X1 port map( A => n1934, Z => n2123);
   U418 : AND2_X1 port map( A1 => DATAIN(0), A2 => n2337, ZN => N128);
   U419 : AND2_X1 port map( A1 => DATAIN(1), A2 => n2337, ZN => N129);
   U420 : AND2_X1 port map( A1 => DATAIN(2), A2 => n2337, ZN => N130);
   U421 : AND2_X1 port map( A1 => DATAIN(3), A2 => n2337, ZN => N131);
   U422 : AND2_X1 port map( A1 => DATAIN(4), A2 => n2337, ZN => N132);
   U423 : AND2_X1 port map( A1 => DATAIN(5), A2 => n2337, ZN => N133);
   U424 : AND2_X1 port map( A1 => DATAIN(6), A2 => n2337, ZN => N134);
   U425 : AND2_X1 port map( A1 => DATAIN(7), A2 => n2337, ZN => N135);
   U426 : AND2_X1 port map( A1 => DATAIN(8), A2 => n2337, ZN => N136);
   U427 : AND2_X1 port map( A1 => DATAIN(9), A2 => n2337, ZN => N137);
   U428 : AND2_X1 port map( A1 => DATAIN(10), A2 => n2337, ZN => N138);
   U429 : AND2_X1 port map( A1 => DATAIN(11), A2 => n2337, ZN => N139);
   U430 : AND2_X1 port map( A1 => DATAIN(12), A2 => n2338, ZN => N140);
   U431 : AND2_X1 port map( A1 => DATAIN(13), A2 => n2338, ZN => N141);
   U432 : AND2_X1 port map( A1 => DATAIN(14), A2 => n2338, ZN => N142);
   U433 : AND2_X1 port map( A1 => DATAIN(15), A2 => n2338, ZN => N143);
   U434 : AND2_X1 port map( A1 => DATAIN(16), A2 => n2338, ZN => N144);
   U435 : AND2_X1 port map( A1 => DATAIN(17), A2 => n2338, ZN => N145);
   U436 : AND2_X1 port map( A1 => DATAIN(18), A2 => n2338, ZN => N146);
   U437 : AND2_X1 port map( A1 => DATAIN(19), A2 => n2338, ZN => N147);
   U438 : AND2_X1 port map( A1 => DATAIN(20), A2 => n2338, ZN => N148);
   U439 : AND2_X1 port map( A1 => DATAIN(21), A2 => n2338, ZN => N149);
   U440 : AND2_X1 port map( A1 => DATAIN(22), A2 => n2338, ZN => N150);
   U441 : AND2_X1 port map( A1 => DATAIN(23), A2 => n2338, ZN => N151);
   U442 : AND2_X1 port map( A1 => DATAIN(24), A2 => n2339, ZN => N152);
   U443 : AND2_X1 port map( A1 => DATAIN(25), A2 => n2339, ZN => N153);
   U444 : AND2_X1 port map( A1 => DATAIN(26), A2 => n2339, ZN => N154);
   U445 : AND2_X1 port map( A1 => DATAIN(27), A2 => n2339, ZN => N155);
   U446 : AND2_X1 port map( A1 => DATAIN(28), A2 => n2339, ZN => N156);
   U447 : AND2_X1 port map( A1 => DATAIN(29), A2 => n2339, ZN => N157);
   U448 : AND2_X1 port map( A1 => DATAIN(30), A2 => n2339, ZN => N158);
   U449 : AND2_X1 port map( A1 => DATAIN(31), A2 => n2339, ZN => N159);
   U450 : OAI222_X1 port map( A1 => n2201, A2 => n3012, B1 => n2197, B2 => 
                           n2372, C1 => n2193, C2 => n2564, ZN => n1406);
   U451 : OAI222_X1 port map( A1 => n2201, A2 => n3011, B1 => n2197, B2 => 
                           n2371, C1 => n2193, C2 => n2563, ZN => n1391);
   U452 : OAI222_X1 port map( A1 => n2201, A2 => n3010, B1 => n2197, B2 => 
                           n2370, C1 => n2193, C2 => n2562, ZN => n1376);
   U453 : OAI222_X1 port map( A1 => n2201, A2 => n3009, B1 => n2197, B2 => 
                           n2369, C1 => n2193, C2 => n2561, ZN => n1361);
   U454 : OAI222_X1 port map( A1 => n2201, A2 => n3008, B1 => n2197, B2 => 
                           n2368, C1 => n2193, C2 => n2560, ZN => n1346);
   U455 : OAI222_X1 port map( A1 => n2201, A2 => n3007, B1 => n2197, B2 => 
                           n2367, C1 => n2193, C2 => n2559, ZN => n1331);
   U456 : OAI222_X1 port map( A1 => n2201, A2 => n3006, B1 => n2197, B2 => 
                           n2366, C1 => n2193, C2 => n2558, ZN => n1316);
   U457 : OAI222_X1 port map( A1 => n2201, A2 => n3005, B1 => n2197, B2 => 
                           n2365, C1 => n2193, C2 => n2557, ZN => n1301);
   U458 : OAI222_X1 port map( A1 => n2201, A2 => n3004, B1 => n2197, B2 => 
                           n2364, C1 => n2193, C2 => n2556, ZN => n1286);
   U459 : OAI222_X1 port map( A1 => n2201, A2 => n3003, B1 => n2197, B2 => 
                           n2363, C1 => n2193, C2 => n2555, ZN => n1271);
   U460 : OAI222_X1 port map( A1 => n2201, A2 => n3002, B1 => n2197, B2 => 
                           n2362, C1 => n2193, C2 => n2554, ZN => n1256);
   U461 : OAI222_X1 port map( A1 => n2201, A2 => n3001, B1 => n2197, B2 => 
                           n2361, C1 => n2193, C2 => n2553, ZN => n1241);
   U462 : OAI222_X1 port map( A1 => n2202, A2 => n3000, B1 => n2198, B2 => 
                           n2360, C1 => n2194, C2 => n2552, ZN => n1226);
   U463 : OAI222_X1 port map( A1 => n2202, A2 => n2999, B1 => n2198, B2 => 
                           n2359, C1 => n2194, C2 => n2551, ZN => n1211);
   U464 : OAI222_X1 port map( A1 => n2202, A2 => n2998, B1 => n2198, B2 => 
                           n2358, C1 => n2194, C2 => n2550, ZN => n1196);
   U465 : OAI222_X1 port map( A1 => n2202, A2 => n2997, B1 => n2198, B2 => 
                           n2357, C1 => n2194, C2 => n2549, ZN => n1181);
   U466 : OAI222_X1 port map( A1 => n2202, A2 => n2996, B1 => n2198, B2 => 
                           n2356, C1 => n2194, C2 => n2548, ZN => n1166);
   U467 : OAI222_X1 port map( A1 => n2202, A2 => n2995, B1 => n2198, B2 => 
                           n2355, C1 => n2194, C2 => n2547, ZN => n1151);
   U468 : OAI222_X1 port map( A1 => n2202, A2 => n2994, B1 => n2198, B2 => 
                           n2354, C1 => n2194, C2 => n2546, ZN => n1136);
   U469 : OAI222_X1 port map( A1 => n2202, A2 => n2993, B1 => n2198, B2 => 
                           n2353, C1 => n2194, C2 => n2545, ZN => n1121);
   U470 : OAI222_X1 port map( A1 => n2202, A2 => n2992, B1 => n2198, B2 => 
                           n2352, C1 => n2194, C2 => n2544, ZN => n1106);
   U471 : OAI222_X1 port map( A1 => n2202, A2 => n2991, B1 => n2198, B2 => 
                           n2351, C1 => n2194, C2 => n2543, ZN => n1091);
   U472 : OAI222_X1 port map( A1 => n2202, A2 => n2990, B1 => n2198, B2 => 
                           n2350, C1 => n2194, C2 => n2542, ZN => n1076);
   U473 : OAI222_X1 port map( A1 => n2202, A2 => n2989, B1 => n2198, B2 => 
                           n2349, C1 => n2194, C2 => n2541, ZN => n1061);
   U474 : OAI222_X1 port map( A1 => n2203, A2 => n2988, B1 => n2199, B2 => 
                           n2348, C1 => n2195, C2 => n2540, ZN => n1046);
   U475 : OAI222_X1 port map( A1 => n2203, A2 => n2987, B1 => n2199, B2 => 
                           n2347, C1 => n2195, C2 => n2539, ZN => n1031);
   U476 : OAI222_X1 port map( A1 => n2203, A2 => n2986, B1 => n2199, B2 => 
                           n2346, C1 => n2195, C2 => n2538, ZN => n1016);
   U477 : OAI222_X1 port map( A1 => n2203, A2 => n2985, B1 => n2199, B2 => 
                           n2345, C1 => n2195, C2 => n2537, ZN => n1001);
   U478 : OAI222_X1 port map( A1 => n2203, A2 => n2984, B1 => n2199, B2 => 
                           n2344, C1 => n2195, C2 => n2536, ZN => n986);
   U479 : OAI222_X1 port map( A1 => n2203, A2 => n2983, B1 => n2199, B2 => 
                           n2343, C1 => n2195, C2 => n2535, ZN => n971);
   U480 : OAI222_X1 port map( A1 => n2203, A2 => n2982, B1 => n2199, B2 => 
                           n2342, C1 => n2195, C2 => n2534, ZN => n956);
   U481 : OAI222_X1 port map( A1 => n2203, A2 => n2981, B1 => n2199, B2 => 
                           n2341, C1 => n2195, C2 => n2533, ZN => n909);
   U482 : OAI222_X1 port map( A1 => n3012, A2 => n2073, B1 => n2372, B2 => 
                           n2069, C1 => n2564, C2 => n2065, ZN => n1921);
   U483 : OAI222_X1 port map( A1 => n3011, A2 => n2073, B1 => n2371, B2 => 
                           n2069, C1 => n2563, C2 => n2065, ZN => n1906);
   U484 : OAI222_X1 port map( A1 => n3010, A2 => n2073, B1 => n2370, B2 => 
                           n2069, C1 => n2562, C2 => n2065, ZN => n1891);
   U485 : OAI222_X1 port map( A1 => n3009, A2 => n2073, B1 => n2369, B2 => 
                           n2069, C1 => n2561, C2 => n2065, ZN => n1876);
   U486 : OAI222_X1 port map( A1 => n3008, A2 => n2073, B1 => n2368, B2 => 
                           n2069, C1 => n2560, C2 => n2065, ZN => n1861);
   U487 : OAI222_X1 port map( A1 => n3007, A2 => n2073, B1 => n2367, B2 => 
                           n2069, C1 => n2559, C2 => n2065, ZN => n1846);
   U488 : OAI222_X1 port map( A1 => n3006, A2 => n2073, B1 => n2366, B2 => 
                           n2069, C1 => n2558, C2 => n2065, ZN => n1831);
   U489 : OAI222_X1 port map( A1 => n3005, A2 => n2073, B1 => n2365, B2 => 
                           n2069, C1 => n2557, C2 => n2065, ZN => n1816);
   U490 : OAI222_X1 port map( A1 => n3004, A2 => n2073, B1 => n2364, B2 => 
                           n2069, C1 => n2556, C2 => n2065, ZN => n1801);
   U491 : OAI222_X1 port map( A1 => n3003, A2 => n2073, B1 => n2363, B2 => 
                           n2069, C1 => n2555, C2 => n2065, ZN => n1786);
   U492 : OAI222_X1 port map( A1 => n3002, A2 => n2073, B1 => n2362, B2 => 
                           n2069, C1 => n2554, C2 => n2065, ZN => n1771);
   U493 : OAI222_X1 port map( A1 => n3001, A2 => n2073, B1 => n2361, B2 => 
                           n2069, C1 => n2553, C2 => n2065, ZN => n1756);
   U494 : OAI222_X1 port map( A1 => n3000, A2 => n2074, B1 => n2360, B2 => 
                           n2070, C1 => n2552, C2 => n2066, ZN => n1741);
   U495 : OAI222_X1 port map( A1 => n2999, A2 => n2074, B1 => n2359, B2 => 
                           n2070, C1 => n2551, C2 => n2066, ZN => n1726);
   U496 : OAI222_X1 port map( A1 => n2998, A2 => n2074, B1 => n2358, B2 => 
                           n2070, C1 => n2550, C2 => n2066, ZN => n1711);
   U497 : OAI222_X1 port map( A1 => n2997, A2 => n2074, B1 => n2357, B2 => 
                           n2070, C1 => n2549, C2 => n2066, ZN => n1696);
   U498 : OAI222_X1 port map( A1 => n2996, A2 => n2074, B1 => n2356, B2 => 
                           n2070, C1 => n2548, C2 => n2066, ZN => n1681);
   U499 : OAI222_X1 port map( A1 => n2995, A2 => n2074, B1 => n2355, B2 => 
                           n2070, C1 => n2547, C2 => n2066, ZN => n1666);
   U500 : OAI222_X1 port map( A1 => n2994, A2 => n2074, B1 => n2354, B2 => 
                           n2070, C1 => n2546, C2 => n2066, ZN => n1651);
   U501 : OAI222_X1 port map( A1 => n2993, A2 => n2074, B1 => n2353, B2 => 
                           n2070, C1 => n2545, C2 => n2066, ZN => n1636);
   U502 : OAI222_X1 port map( A1 => n2992, A2 => n2074, B1 => n2352, B2 => 
                           n2070, C1 => n2544, C2 => n2066, ZN => n1621);
   U503 : OAI222_X1 port map( A1 => n2991, A2 => n2074, B1 => n2351, B2 => 
                           n2070, C1 => n2543, C2 => n2066, ZN => n1606);
   U504 : OAI222_X1 port map( A1 => n2990, A2 => n2074, B1 => n2350, B2 => 
                           n2070, C1 => n2542, C2 => n2066, ZN => n1591);
   U505 : OAI222_X1 port map( A1 => n2989, A2 => n2074, B1 => n2349, B2 => 
                           n2070, C1 => n2541, C2 => n2066, ZN => n1576);
   U506 : OAI222_X1 port map( A1 => n2988, A2 => n2075, B1 => n2348, B2 => 
                           n2071, C1 => n2540, C2 => n2067, ZN => n1561);
   U507 : OAI222_X1 port map( A1 => n2987, A2 => n2075, B1 => n2347, B2 => 
                           n2071, C1 => n2539, C2 => n2067, ZN => n1546);
   U508 : OAI222_X1 port map( A1 => n2986, A2 => n2075, B1 => n2346, B2 => 
                           n2071, C1 => n2538, C2 => n2067, ZN => n1531);
   U509 : OAI222_X1 port map( A1 => n2985, A2 => n2075, B1 => n2345, B2 => 
                           n2071, C1 => n2537, C2 => n2067, ZN => n1516);
   U510 : OAI222_X1 port map( A1 => n2984, A2 => n2075, B1 => n2344, B2 => 
                           n2071, C1 => n2536, C2 => n2067, ZN => n1501);
   U511 : OAI222_X1 port map( A1 => n2983, A2 => n2075, B1 => n2343, B2 => 
                           n2071, C1 => n2535, C2 => n2067, ZN => n1486);
   U512 : OAI222_X1 port map( A1 => n2982, A2 => n2075, B1 => n2342, B2 => 
                           n2071, C1 => n2534, C2 => n2067, ZN => n1471);
   U513 : OAI222_X1 port map( A1 => n2981, A2 => n2075, B1 => n2341, B2 => 
                           n2071, C1 => n2533, C2 => n2067, ZN => n1424);
   U514 : OAI222_X1 port map( A1 => n2189, A2 => n2436, B1 => n2185, B2 => 
                           n3108, C1 => n2181, C2 => n3076, ZN => n1405);
   U515 : OAI222_X1 port map( A1 => n2109, A2 => n2820, B1 => n2105, B2 => 
                           n2852, C1 => n2101, C2 => n2756, ZN => n1411);
   U516 : OAI222_X1 port map( A1 => n2189, A2 => n2435, B1 => n2185, B2 => 
                           n3107, C1 => n2181, C2 => n3075, ZN => n1390);
   U517 : OAI222_X1 port map( A1 => n2109, A2 => n2819, B1 => n2105, B2 => 
                           n2851, C1 => n2101, C2 => n2755, ZN => n1394);
   U518 : OAI222_X1 port map( A1 => n2189, A2 => n2434, B1 => n2185, B2 => 
                           n3106, C1 => n2181, C2 => n3074, ZN => n1375);
   U519 : OAI222_X1 port map( A1 => n2109, A2 => n2818, B1 => n2105, B2 => 
                           n2850, C1 => n2101, C2 => n2754, ZN => n1379);
   U520 : OAI222_X1 port map( A1 => n2189, A2 => n2433, B1 => n2185, B2 => 
                           n3105, C1 => n2181, C2 => n3073, ZN => n1360);
   U521 : OAI222_X1 port map( A1 => n2109, A2 => n2817, B1 => n2105, B2 => 
                           n2849, C1 => n2101, C2 => n2753, ZN => n1364);
   U522 : OAI222_X1 port map( A1 => n2189, A2 => n2432, B1 => n2185, B2 => 
                           n3104, C1 => n2181, C2 => n3072, ZN => n1345);
   U523 : OAI222_X1 port map( A1 => n2109, A2 => n2816, B1 => n2105, B2 => 
                           n2848, C1 => n2101, C2 => n2752, ZN => n1349);
   U524 : OAI222_X1 port map( A1 => n2189, A2 => n2431, B1 => n2185, B2 => 
                           n3103, C1 => n2181, C2 => n3071, ZN => n1330);
   U525 : OAI222_X1 port map( A1 => n2109, A2 => n2815, B1 => n2105, B2 => 
                           n2847, C1 => n2101, C2 => n2751, ZN => n1334);
   U526 : OAI222_X1 port map( A1 => n2189, A2 => n2430, B1 => n2185, B2 => 
                           n3102, C1 => n2181, C2 => n3070, ZN => n1315);
   U527 : OAI222_X1 port map( A1 => n2109, A2 => n2814, B1 => n2105, B2 => 
                           n2846, C1 => n2101, C2 => n2750, ZN => n1319);
   U528 : OAI222_X1 port map( A1 => n2189, A2 => n2429, B1 => n2185, B2 => 
                           n3101, C1 => n2181, C2 => n3069, ZN => n1300);
   U529 : OAI222_X1 port map( A1 => n2109, A2 => n2813, B1 => n2105, B2 => 
                           n2845, C1 => n2101, C2 => n2749, ZN => n1304);
   U530 : OAI222_X1 port map( A1 => n2189, A2 => n2428, B1 => n2185, B2 => 
                           n3100, C1 => n2181, C2 => n3068, ZN => n1285);
   U531 : OAI222_X1 port map( A1 => n2109, A2 => n2812, B1 => n2105, B2 => 
                           n2844, C1 => n2101, C2 => n2748, ZN => n1289);
   U532 : OAI222_X1 port map( A1 => n2189, A2 => n2427, B1 => n2185, B2 => 
                           n3099, C1 => n2181, C2 => n3067, ZN => n1270);
   U533 : OAI222_X1 port map( A1 => n2109, A2 => n2811, B1 => n2105, B2 => 
                           n2843, C1 => n2101, C2 => n2747, ZN => n1274);
   U534 : OAI222_X1 port map( A1 => n2189, A2 => n2426, B1 => n2185, B2 => 
                           n3098, C1 => n2181, C2 => n3066, ZN => n1255);
   U535 : OAI222_X1 port map( A1 => n2109, A2 => n2810, B1 => n2105, B2 => 
                           n2842, C1 => n2101, C2 => n2746, ZN => n1259);
   U536 : OAI222_X1 port map( A1 => n2189, A2 => n2425, B1 => n2185, B2 => 
                           n3097, C1 => n2181, C2 => n3065, ZN => n1240);
   U537 : OAI222_X1 port map( A1 => n2109, A2 => n2809, B1 => n2105, B2 => 
                           n2841, C1 => n2101, C2 => n2745, ZN => n1244);
   U538 : OAI222_X1 port map( A1 => n2190, A2 => n2424, B1 => n2186, B2 => 
                           n3096, C1 => n2182, C2 => n3064, ZN => n1225);
   U539 : OAI222_X1 port map( A1 => n2110, A2 => n2808, B1 => n2106, B2 => 
                           n2840, C1 => n2102, C2 => n2744, ZN => n1229);
   U540 : OAI222_X1 port map( A1 => n2190, A2 => n2423, B1 => n2186, B2 => 
                           n3095, C1 => n2182, C2 => n3063, ZN => n1210);
   U541 : OAI222_X1 port map( A1 => n2110, A2 => n2807, B1 => n2106, B2 => 
                           n2839, C1 => n2102, C2 => n2743, ZN => n1214);
   U542 : OAI222_X1 port map( A1 => n2190, A2 => n2422, B1 => n2186, B2 => 
                           n3094, C1 => n2182, C2 => n3062, ZN => n1195);
   U543 : OAI222_X1 port map( A1 => n2110, A2 => n2806, B1 => n2106, B2 => 
                           n2838, C1 => n2102, C2 => n2742, ZN => n1199);
   U544 : OAI222_X1 port map( A1 => n2190, A2 => n2421, B1 => n2186, B2 => 
                           n3093, C1 => n2182, C2 => n3061, ZN => n1180);
   U545 : OAI222_X1 port map( A1 => n2110, A2 => n2805, B1 => n2106, B2 => 
                           n2837, C1 => n2102, C2 => n2741, ZN => n1184);
   U546 : OAI222_X1 port map( A1 => n2190, A2 => n2420, B1 => n2186, B2 => 
                           n3092, C1 => n2182, C2 => n3060, ZN => n1165);
   U547 : OAI222_X1 port map( A1 => n2110, A2 => n2804, B1 => n2106, B2 => 
                           n2836, C1 => n2102, C2 => n2740, ZN => n1169);
   U548 : OAI222_X1 port map( A1 => n2190, A2 => n2419, B1 => n2186, B2 => 
                           n3091, C1 => n2182, C2 => n3059, ZN => n1150);
   U549 : OAI222_X1 port map( A1 => n2110, A2 => n2803, B1 => n2106, B2 => 
                           n2835, C1 => n2102, C2 => n2739, ZN => n1154);
   U550 : OAI222_X1 port map( A1 => n2190, A2 => n2418, B1 => n2186, B2 => 
                           n3090, C1 => n2182, C2 => n3058, ZN => n1135);
   U551 : OAI222_X1 port map( A1 => n2110, A2 => n2802, B1 => n2106, B2 => 
                           n2834, C1 => n2102, C2 => n2738, ZN => n1139);
   U552 : OAI222_X1 port map( A1 => n2190, A2 => n2417, B1 => n2186, B2 => 
                           n3089, C1 => n2182, C2 => n3057, ZN => n1120);
   U553 : OAI222_X1 port map( A1 => n2110, A2 => n2801, B1 => n2106, B2 => 
                           n2833, C1 => n2102, C2 => n2737, ZN => n1124);
   U554 : OAI222_X1 port map( A1 => n2190, A2 => n2416, B1 => n2186, B2 => 
                           n3088, C1 => n2182, C2 => n3056, ZN => n1105);
   U555 : OAI222_X1 port map( A1 => n2110, A2 => n2800, B1 => n2106, B2 => 
                           n2832, C1 => n2102, C2 => n2736, ZN => n1109);
   U556 : OAI222_X1 port map( A1 => n2190, A2 => n2415, B1 => n2186, B2 => 
                           n3087, C1 => n2182, C2 => n3055, ZN => n1090);
   U557 : OAI222_X1 port map( A1 => n2110, A2 => n2799, B1 => n2106, B2 => 
                           n2831, C1 => n2102, C2 => n2735, ZN => n1094);
   U558 : OAI222_X1 port map( A1 => n2190, A2 => n2414, B1 => n2186, B2 => 
                           n3086, C1 => n2182, C2 => n3054, ZN => n1075);
   U559 : OAI222_X1 port map( A1 => n2110, A2 => n2798, B1 => n2106, B2 => 
                           n2830, C1 => n2102, C2 => n2734, ZN => n1079);
   U560 : OAI222_X1 port map( A1 => n2190, A2 => n2413, B1 => n2186, B2 => 
                           n3085, C1 => n2182, C2 => n3053, ZN => n1060);
   U561 : OAI222_X1 port map( A1 => n2110, A2 => n2797, B1 => n2106, B2 => 
                           n2829, C1 => n2102, C2 => n2733, ZN => n1064);
   U562 : OAI222_X1 port map( A1 => n2191, A2 => n2412, B1 => n2187, B2 => 
                           n3084, C1 => n2183, C2 => n3052, ZN => n1045);
   U563 : OAI222_X1 port map( A1 => n2111, A2 => n2796, B1 => n2107, B2 => 
                           n2828, C1 => n2103, C2 => n2732, ZN => n1049);
   U564 : OAI222_X1 port map( A1 => n2191, A2 => n2411, B1 => n2187, B2 => 
                           n3083, C1 => n2183, C2 => n3051, ZN => n1030);
   U565 : OAI222_X1 port map( A1 => n2111, A2 => n2795, B1 => n2107, B2 => 
                           n2827, C1 => n2103, C2 => n2731, ZN => n1034);
   U566 : OAI222_X1 port map( A1 => n2191, A2 => n2410, B1 => n2187, B2 => 
                           n3082, C1 => n2183, C2 => n3050, ZN => n1015);
   U567 : OAI222_X1 port map( A1 => n2111, A2 => n2794, B1 => n2107, B2 => 
                           n2826, C1 => n2103, C2 => n2730, ZN => n1019);
   U568 : OAI222_X1 port map( A1 => n2191, A2 => n2409, B1 => n2187, B2 => 
                           n3081, C1 => n2183, C2 => n3049, ZN => n1000);
   U569 : OAI222_X1 port map( A1 => n2111, A2 => n2793, B1 => n2107, B2 => 
                           n2825, C1 => n2103, C2 => n2729, ZN => n1004);
   U570 : OAI222_X1 port map( A1 => n2191, A2 => n2408, B1 => n2187, B2 => 
                           n3080, C1 => n2183, C2 => n3048, ZN => n985);
   U571 : OAI222_X1 port map( A1 => n2111, A2 => n2792, B1 => n2107, B2 => 
                           n2824, C1 => n2103, C2 => n2728, ZN => n989);
   U572 : OAI222_X1 port map( A1 => n2191, A2 => n2407, B1 => n2187, B2 => 
                           n3079, C1 => n2183, C2 => n3047, ZN => n970);
   U573 : OAI222_X1 port map( A1 => n2111, A2 => n2791, B1 => n2107, B2 => 
                           n2823, C1 => n2103, C2 => n2727, ZN => n974);
   U574 : OAI222_X1 port map( A1 => n2191, A2 => n2406, B1 => n2187, B2 => 
                           n3078, C1 => n2183, C2 => n3046, ZN => n955);
   U575 : OAI222_X1 port map( A1 => n2111, A2 => n2790, B1 => n2107, B2 => 
                           n2822, C1 => n2103, C2 => n2726, ZN => n959);
   U576 : OAI222_X1 port map( A1 => n2191, A2 => n2405, B1 => n2187, B2 => 
                           n3077, C1 => n2183, C2 => n3045, ZN => n908);
   U577 : OAI222_X1 port map( A1 => n2111, A2 => n2789, B1 => n2107, B2 => 
                           n2821, C1 => n2103, C2 => n2725, ZN => n924);
   U578 : OAI222_X1 port map( A1 => n2436, A2 => n2061, B1 => n3108, B2 => 
                           n2057, C1 => n3076, C2 => n2053, ZN => n1920);
   U579 : OAI222_X1 port map( A1 => n2820, A2 => n1981, B1 => n2852, B2 => 
                           n1977, C1 => n2756, C2 => n1973, ZN => n1926);
   U580 : OAI222_X1 port map( A1 => n2435, A2 => n2061, B1 => n3107, B2 => 
                           n2057, C1 => n3075, C2 => n2053, ZN => n1905);
   U581 : OAI222_X1 port map( A1 => n2819, A2 => n1981, B1 => n2851, B2 => 
                           n1977, C1 => n2755, C2 => n1973, ZN => n1909);
   U582 : OAI222_X1 port map( A1 => n2434, A2 => n2061, B1 => n3106, B2 => 
                           n2057, C1 => n3074, C2 => n2053, ZN => n1890);
   U583 : OAI222_X1 port map( A1 => n2818, A2 => n1981, B1 => n2850, B2 => 
                           n1977, C1 => n2754, C2 => n1973, ZN => n1894);
   U584 : OAI222_X1 port map( A1 => n2433, A2 => n2061, B1 => n3105, B2 => 
                           n2057, C1 => n3073, C2 => n2053, ZN => n1875);
   U585 : OAI222_X1 port map( A1 => n2817, A2 => n1981, B1 => n2849, B2 => 
                           n1977, C1 => n2753, C2 => n1973, ZN => n1879);
   U586 : OAI222_X1 port map( A1 => n2432, A2 => n2061, B1 => n3104, B2 => 
                           n2057, C1 => n3072, C2 => n2053, ZN => n1860);
   U587 : OAI222_X1 port map( A1 => n2816, A2 => n1981, B1 => n2848, B2 => 
                           n1977, C1 => n2752, C2 => n1973, ZN => n1864);
   U588 : OAI222_X1 port map( A1 => n2431, A2 => n2061, B1 => n3103, B2 => 
                           n2057, C1 => n3071, C2 => n2053, ZN => n1845);
   U589 : OAI222_X1 port map( A1 => n2815, A2 => n1981, B1 => n2847, B2 => 
                           n1977, C1 => n2751, C2 => n1973, ZN => n1849);
   U590 : OAI222_X1 port map( A1 => n2430, A2 => n2061, B1 => n3102, B2 => 
                           n2057, C1 => n3070, C2 => n2053, ZN => n1830);
   U591 : OAI222_X1 port map( A1 => n2814, A2 => n1981, B1 => n2846, B2 => 
                           n1977, C1 => n2750, C2 => n1973, ZN => n1834);
   U592 : OAI222_X1 port map( A1 => n2429, A2 => n2061, B1 => n3101, B2 => 
                           n2057, C1 => n3069, C2 => n2053, ZN => n1815);
   U593 : OAI222_X1 port map( A1 => n2813, A2 => n1981, B1 => n2845, B2 => 
                           n1977, C1 => n2749, C2 => n1973, ZN => n1819);
   U594 : OAI222_X1 port map( A1 => n2428, A2 => n2061, B1 => n3100, B2 => 
                           n2057, C1 => n3068, C2 => n2053, ZN => n1800);
   U595 : OAI222_X1 port map( A1 => n2812, A2 => n1981, B1 => n2844, B2 => 
                           n1977, C1 => n2748, C2 => n1973, ZN => n1804);
   U596 : OAI222_X1 port map( A1 => n2427, A2 => n2061, B1 => n3099, B2 => 
                           n2057, C1 => n3067, C2 => n2053, ZN => n1785);
   U597 : OAI222_X1 port map( A1 => n2811, A2 => n1981, B1 => n2843, B2 => 
                           n1977, C1 => n2747, C2 => n1973, ZN => n1789);
   U598 : OAI222_X1 port map( A1 => n2426, A2 => n2061, B1 => n3098, B2 => 
                           n2057, C1 => n3066, C2 => n2053, ZN => n1770);
   U599 : OAI222_X1 port map( A1 => n2810, A2 => n1981, B1 => n2842, B2 => 
                           n1977, C1 => n2746, C2 => n1973, ZN => n1774);
   U600 : OAI222_X1 port map( A1 => n2425, A2 => n2061, B1 => n3097, B2 => 
                           n2057, C1 => n3065, C2 => n2053, ZN => n1755);
   U601 : OAI222_X1 port map( A1 => n2809, A2 => n1981, B1 => n2841, B2 => 
                           n1977, C1 => n2745, C2 => n1973, ZN => n1759);
   U602 : OAI222_X1 port map( A1 => n2424, A2 => n2062, B1 => n3096, B2 => 
                           n2058, C1 => n3064, C2 => n2054, ZN => n1740);
   U603 : OAI222_X1 port map( A1 => n2808, A2 => n1982, B1 => n2840, B2 => 
                           n1978, C1 => n2744, C2 => n1974, ZN => n1744);
   U604 : OAI222_X1 port map( A1 => n2423, A2 => n2062, B1 => n3095, B2 => 
                           n2058, C1 => n3063, C2 => n2054, ZN => n1725);
   U605 : OAI222_X1 port map( A1 => n2807, A2 => n1982, B1 => n2839, B2 => 
                           n1978, C1 => n2743, C2 => n1974, ZN => n1729);
   U606 : OAI222_X1 port map( A1 => n2422, A2 => n2062, B1 => n3094, B2 => 
                           n2058, C1 => n3062, C2 => n2054, ZN => n1710);
   U607 : OAI222_X1 port map( A1 => n2806, A2 => n1982, B1 => n2838, B2 => 
                           n1978, C1 => n2742, C2 => n1974, ZN => n1714);
   U608 : OAI222_X1 port map( A1 => n2421, A2 => n2062, B1 => n3093, B2 => 
                           n2058, C1 => n3061, C2 => n2054, ZN => n1695);
   U609 : OAI222_X1 port map( A1 => n2805, A2 => n1982, B1 => n2837, B2 => 
                           n1978, C1 => n2741, C2 => n1974, ZN => n1699);
   U610 : OAI222_X1 port map( A1 => n2420, A2 => n2062, B1 => n3092, B2 => 
                           n2058, C1 => n3060, C2 => n2054, ZN => n1680);
   U611 : OAI222_X1 port map( A1 => n2804, A2 => n1982, B1 => n2836, B2 => 
                           n1978, C1 => n2740, C2 => n1974, ZN => n1684);
   U612 : OAI222_X1 port map( A1 => n2419, A2 => n2062, B1 => n3091, B2 => 
                           n2058, C1 => n3059, C2 => n2054, ZN => n1665);
   U613 : OAI222_X1 port map( A1 => n2803, A2 => n1982, B1 => n2835, B2 => 
                           n1978, C1 => n2739, C2 => n1974, ZN => n1669);
   U614 : OAI222_X1 port map( A1 => n2418, A2 => n2062, B1 => n3090, B2 => 
                           n2058, C1 => n3058, C2 => n2054, ZN => n1650);
   U615 : OAI222_X1 port map( A1 => n2802, A2 => n1982, B1 => n2834, B2 => 
                           n1978, C1 => n2738, C2 => n1974, ZN => n1654);
   U616 : OAI222_X1 port map( A1 => n2417, A2 => n2062, B1 => n3089, B2 => 
                           n2058, C1 => n3057, C2 => n2054, ZN => n1635);
   U617 : OAI222_X1 port map( A1 => n2801, A2 => n1982, B1 => n2833, B2 => 
                           n1978, C1 => n2737, C2 => n1974, ZN => n1639);
   U618 : OAI222_X1 port map( A1 => n2416, A2 => n2062, B1 => n3088, B2 => 
                           n2058, C1 => n3056, C2 => n2054, ZN => n1620);
   U619 : OAI222_X1 port map( A1 => n2800, A2 => n1982, B1 => n2832, B2 => 
                           n1978, C1 => n2736, C2 => n1974, ZN => n1624);
   U620 : OAI222_X1 port map( A1 => n2415, A2 => n2062, B1 => n3087, B2 => 
                           n2058, C1 => n3055, C2 => n2054, ZN => n1605);
   U621 : OAI222_X1 port map( A1 => n2799, A2 => n1982, B1 => n2831, B2 => 
                           n1978, C1 => n2735, C2 => n1974, ZN => n1609);
   U622 : OAI222_X1 port map( A1 => n2414, A2 => n2062, B1 => n3086, B2 => 
                           n2058, C1 => n3054, C2 => n2054, ZN => n1590);
   U623 : OAI222_X1 port map( A1 => n2798, A2 => n1982, B1 => n2830, B2 => 
                           n1978, C1 => n2734, C2 => n1974, ZN => n1594);
   U624 : OAI222_X1 port map( A1 => n2413, A2 => n2062, B1 => n3085, B2 => 
                           n2058, C1 => n3053, C2 => n2054, ZN => n1575);
   U625 : OAI222_X1 port map( A1 => n2797, A2 => n1982, B1 => n2829, B2 => 
                           n1978, C1 => n2733, C2 => n1974, ZN => n1579);
   U626 : OAI222_X1 port map( A1 => n2412, A2 => n2063, B1 => n3084, B2 => 
                           n2059, C1 => n3052, C2 => n2055, ZN => n1560);
   U627 : OAI222_X1 port map( A1 => n2796, A2 => n1983, B1 => n2828, B2 => 
                           n1979, C1 => n2732, C2 => n1975, ZN => n1564);
   U628 : OAI222_X1 port map( A1 => n2411, A2 => n2063, B1 => n3083, B2 => 
                           n2059, C1 => n3051, C2 => n2055, ZN => n1545);
   U629 : OAI222_X1 port map( A1 => n2795, A2 => n1983, B1 => n2827, B2 => 
                           n1979, C1 => n2731, C2 => n1975, ZN => n1549);
   U630 : OAI222_X1 port map( A1 => n2410, A2 => n2063, B1 => n3082, B2 => 
                           n2059, C1 => n3050, C2 => n2055, ZN => n1530);
   U631 : OAI222_X1 port map( A1 => n2794, A2 => n1983, B1 => n2826, B2 => 
                           n1979, C1 => n2730, C2 => n1975, ZN => n1534);
   U632 : OAI222_X1 port map( A1 => n2409, A2 => n2063, B1 => n3081, B2 => 
                           n2059, C1 => n3049, C2 => n2055, ZN => n1515);
   U633 : OAI222_X1 port map( A1 => n2793, A2 => n1983, B1 => n2825, B2 => 
                           n1979, C1 => n2729, C2 => n1975, ZN => n1519);
   U634 : OAI222_X1 port map( A1 => n2408, A2 => n2063, B1 => n3080, B2 => 
                           n2059, C1 => n3048, C2 => n2055, ZN => n1500);
   U635 : OAI222_X1 port map( A1 => n2792, A2 => n1983, B1 => n2824, B2 => 
                           n1979, C1 => n2728, C2 => n1975, ZN => n1504);
   U636 : OAI222_X1 port map( A1 => n2407, A2 => n2063, B1 => n3079, B2 => 
                           n2059, C1 => n3047, C2 => n2055, ZN => n1485);
   U637 : OAI222_X1 port map( A1 => n2791, A2 => n1983, B1 => n2823, B2 => 
                           n1979, C1 => n2727, C2 => n1975, ZN => n1489);
   U638 : OAI222_X1 port map( A1 => n2406, A2 => n2063, B1 => n3078, B2 => 
                           n2059, C1 => n3046, C2 => n2055, ZN => n1470);
   U639 : OAI222_X1 port map( A1 => n2790, A2 => n1983, B1 => n2822, B2 => 
                           n1979, C1 => n2726, C2 => n1975, ZN => n1474);
   U640 : OAI222_X1 port map( A1 => n2405, A2 => n2063, B1 => n3077, B2 => 
                           n2059, C1 => n3045, C2 => n2055, ZN => n1423);
   U641 : OAI222_X1 port map( A1 => n2789, A2 => n1983, B1 => n2821, B2 => 
                           n1979, C1 => n2725, C2 => n1975, ZN => n1439);
   U642 : OAI222_X1 port map( A1 => n2177, A2 => n3172, B1 => n2173, B2 => 
                           n2532, C1 => n2169, C2 => n2468, ZN => n1404);
   U643 : OAI222_X1 port map( A1 => n2097, A2 => n2724, B1 => n2093, B2 => 
                           n2788, C1 => n2089, C2 => n2916, ZN => n1410);
   U644 : OAI222_X1 port map( A1 => n2177, A2 => n3171, B1 => n2173, B2 => 
                           n2531, C1 => n2169, C2 => n2467, ZN => n1389);
   U645 : OAI222_X1 port map( A1 => n2097, A2 => n2723, B1 => n2093, B2 => 
                           n2787, C1 => n2089, C2 => n2915, ZN => n1393);
   U646 : OAI222_X1 port map( A1 => n2177, A2 => n3170, B1 => n2173, B2 => 
                           n2530, C1 => n2169, C2 => n2466, ZN => n1374);
   U647 : OAI222_X1 port map( A1 => n2097, A2 => n2722, B1 => n2093, B2 => 
                           n2786, C1 => n2089, C2 => n2914, ZN => n1378);
   U648 : OAI222_X1 port map( A1 => n2177, A2 => n3169, B1 => n2173, B2 => 
                           n2529, C1 => n2169, C2 => n2465, ZN => n1359);
   U649 : OAI222_X1 port map( A1 => n2097, A2 => n2721, B1 => n2093, B2 => 
                           n2785, C1 => n2089, C2 => n2913, ZN => n1363);
   U650 : OAI222_X1 port map( A1 => n2177, A2 => n3168, B1 => n2173, B2 => 
                           n2528, C1 => n2169, C2 => n2464, ZN => n1344);
   U651 : OAI222_X1 port map( A1 => n2097, A2 => n2720, B1 => n2093, B2 => 
                           n2784, C1 => n2089, C2 => n2912, ZN => n1348);
   U652 : OAI222_X1 port map( A1 => n2177, A2 => n3167, B1 => n2173, B2 => 
                           n2527, C1 => n2169, C2 => n2463, ZN => n1329);
   U653 : OAI222_X1 port map( A1 => n2097, A2 => n2719, B1 => n2093, B2 => 
                           n2783, C1 => n2089, C2 => n2911, ZN => n1333);
   U654 : OAI222_X1 port map( A1 => n2177, A2 => n3166, B1 => n2173, B2 => 
                           n2526, C1 => n2169, C2 => n2462, ZN => n1314);
   U655 : OAI222_X1 port map( A1 => n2097, A2 => n2718, B1 => n2093, B2 => 
                           n2782, C1 => n2089, C2 => n2910, ZN => n1318);
   U656 : OAI222_X1 port map( A1 => n2177, A2 => n3165, B1 => n2173, B2 => 
                           n2525, C1 => n2169, C2 => n2461, ZN => n1299);
   U657 : OAI222_X1 port map( A1 => n2097, A2 => n2717, B1 => n2093, B2 => 
                           n2781, C1 => n2089, C2 => n2909, ZN => n1303);
   U658 : OAI222_X1 port map( A1 => n2177, A2 => n3164, B1 => n2173, B2 => 
                           n2524, C1 => n2169, C2 => n2460, ZN => n1284);
   U659 : OAI222_X1 port map( A1 => n2097, A2 => n2716, B1 => n2093, B2 => 
                           n2780, C1 => n2089, C2 => n2908, ZN => n1288);
   U660 : OAI222_X1 port map( A1 => n2177, A2 => n3163, B1 => n2173, B2 => 
                           n2523, C1 => n2169, C2 => n2459, ZN => n1269);
   U661 : OAI222_X1 port map( A1 => n2097, A2 => n2715, B1 => n2093, B2 => 
                           n2779, C1 => n2089, C2 => n2907, ZN => n1273);
   U662 : OAI222_X1 port map( A1 => n2177, A2 => n3162, B1 => n2173, B2 => 
                           n2522, C1 => n2169, C2 => n2458, ZN => n1254);
   U663 : OAI222_X1 port map( A1 => n2097, A2 => n2714, B1 => n2093, B2 => 
                           n2778, C1 => n2089, C2 => n2906, ZN => n1258);
   U664 : OAI222_X1 port map( A1 => n2177, A2 => n3161, B1 => n2173, B2 => 
                           n2521, C1 => n2169, C2 => n2457, ZN => n1239);
   U665 : OAI222_X1 port map( A1 => n2097, A2 => n2713, B1 => n2093, B2 => 
                           n2777, C1 => n2089, C2 => n2905, ZN => n1243);
   U666 : OAI222_X1 port map( A1 => n2178, A2 => n3160, B1 => n2174, B2 => 
                           n2520, C1 => n2170, C2 => n2456, ZN => n1224);
   U667 : OAI222_X1 port map( A1 => n2098, A2 => n2712, B1 => n2094, B2 => 
                           n2776, C1 => n2090, C2 => n2904, ZN => n1228);
   U668 : OAI222_X1 port map( A1 => n2178, A2 => n3159, B1 => n2174, B2 => 
                           n2519, C1 => n2170, C2 => n2455, ZN => n1209);
   U669 : OAI222_X1 port map( A1 => n2098, A2 => n2711, B1 => n2094, B2 => 
                           n2775, C1 => n2090, C2 => n2903, ZN => n1213);
   U670 : OAI222_X1 port map( A1 => n2178, A2 => n3158, B1 => n2174, B2 => 
                           n2518, C1 => n2170, C2 => n2454, ZN => n1194);
   U671 : OAI222_X1 port map( A1 => n2098, A2 => n2710, B1 => n2094, B2 => 
                           n2774, C1 => n2090, C2 => n2902, ZN => n1198);
   U672 : OAI222_X1 port map( A1 => n2178, A2 => n3157, B1 => n2174, B2 => 
                           n2517, C1 => n2170, C2 => n2453, ZN => n1179);
   U673 : OAI222_X1 port map( A1 => n2098, A2 => n2709, B1 => n2094, B2 => 
                           n2773, C1 => n2090, C2 => n2901, ZN => n1183);
   U674 : OAI222_X1 port map( A1 => n2178, A2 => n3156, B1 => n2174, B2 => 
                           n2516, C1 => n2170, C2 => n2452, ZN => n1164);
   U675 : OAI222_X1 port map( A1 => n2098, A2 => n2708, B1 => n2094, B2 => 
                           n2772, C1 => n2090, C2 => n2900, ZN => n1168);
   U676 : OAI222_X1 port map( A1 => n2178, A2 => n3155, B1 => n2174, B2 => 
                           n2515, C1 => n2170, C2 => n2451, ZN => n1149);
   U677 : OAI222_X1 port map( A1 => n2098, A2 => n2707, B1 => n2094, B2 => 
                           n2771, C1 => n2090, C2 => n2899, ZN => n1153);
   U678 : OAI222_X1 port map( A1 => n2178, A2 => n3154, B1 => n2174, B2 => 
                           n2514, C1 => n2170, C2 => n2450, ZN => n1134);
   U679 : OAI222_X1 port map( A1 => n2098, A2 => n2706, B1 => n2094, B2 => 
                           n2770, C1 => n2090, C2 => n2898, ZN => n1138);
   U680 : OAI222_X1 port map( A1 => n2178, A2 => n3153, B1 => n2174, B2 => 
                           n2513, C1 => n2170, C2 => n2449, ZN => n1119);
   U681 : OAI222_X1 port map( A1 => n2098, A2 => n2705, B1 => n2094, B2 => 
                           n2769, C1 => n2090, C2 => n2897, ZN => n1123);
   U682 : OAI222_X1 port map( A1 => n2178, A2 => n3152, B1 => n2174, B2 => 
                           n2512, C1 => n2170, C2 => n2448, ZN => n1104);
   U683 : OAI222_X1 port map( A1 => n2098, A2 => n2704, B1 => n2094, B2 => 
                           n2768, C1 => n2090, C2 => n2896, ZN => n1108);
   U684 : OAI222_X1 port map( A1 => n2178, A2 => n3151, B1 => n2174, B2 => 
                           n2511, C1 => n2170, C2 => n2447, ZN => n1089);
   U685 : OAI222_X1 port map( A1 => n2098, A2 => n2703, B1 => n2094, B2 => 
                           n2767, C1 => n2090, C2 => n2895, ZN => n1093);
   U686 : OAI222_X1 port map( A1 => n2178, A2 => n3150, B1 => n2174, B2 => 
                           n2510, C1 => n2170, C2 => n2446, ZN => n1074);
   U687 : OAI222_X1 port map( A1 => n2098, A2 => n2702, B1 => n2094, B2 => 
                           n2766, C1 => n2090, C2 => n2894, ZN => n1078);
   U688 : OAI222_X1 port map( A1 => n2178, A2 => n3149, B1 => n2174, B2 => 
                           n2509, C1 => n2170, C2 => n2445, ZN => n1059);
   U689 : OAI222_X1 port map( A1 => n2098, A2 => n2701, B1 => n2094, B2 => 
                           n2765, C1 => n2090, C2 => n2893, ZN => n1063);
   U690 : OAI222_X1 port map( A1 => n2179, A2 => n3148, B1 => n2175, B2 => 
                           n2508, C1 => n2171, C2 => n2444, ZN => n1044);
   U691 : OAI222_X1 port map( A1 => n2099, A2 => n2700, B1 => n2095, B2 => 
                           n2764, C1 => n2091, C2 => n2892, ZN => n1048);
   U692 : OAI222_X1 port map( A1 => n2179, A2 => n3147, B1 => n2175, B2 => 
                           n2507, C1 => n2171, C2 => n2443, ZN => n1029);
   U693 : OAI222_X1 port map( A1 => n2099, A2 => n2699, B1 => n2095, B2 => 
                           n2763, C1 => n2091, C2 => n2891, ZN => n1033);
   U694 : OAI222_X1 port map( A1 => n2179, A2 => n3146, B1 => n2175, B2 => 
                           n2506, C1 => n2171, C2 => n2442, ZN => n1014);
   U695 : OAI222_X1 port map( A1 => n2099, A2 => n2698, B1 => n2095, B2 => 
                           n2762, C1 => n2091, C2 => n2890, ZN => n1018);
   U696 : OAI222_X1 port map( A1 => n2179, A2 => n3145, B1 => n2175, B2 => 
                           n2505, C1 => n2171, C2 => n2441, ZN => n999);
   U697 : OAI222_X1 port map( A1 => n2099, A2 => n2697, B1 => n2095, B2 => 
                           n2761, C1 => n2091, C2 => n2889, ZN => n1003);
   U698 : OAI222_X1 port map( A1 => n2179, A2 => n3144, B1 => n2175, B2 => 
                           n2504, C1 => n2171, C2 => n2440, ZN => n984);
   U699 : OAI222_X1 port map( A1 => n2099, A2 => n2696, B1 => n2095, B2 => 
                           n2760, C1 => n2091, C2 => n2888, ZN => n988);
   U700 : OAI222_X1 port map( A1 => n2179, A2 => n3143, B1 => n2175, B2 => 
                           n2503, C1 => n2171, C2 => n2439, ZN => n969);
   U701 : OAI222_X1 port map( A1 => n2099, A2 => n2695, B1 => n2095, B2 => 
                           n2759, C1 => n2091, C2 => n2887, ZN => n973);
   U702 : OAI222_X1 port map( A1 => n2179, A2 => n3142, B1 => n2175, B2 => 
                           n2502, C1 => n2171, C2 => n2438, ZN => n954);
   U703 : OAI222_X1 port map( A1 => n2099, A2 => n2694, B1 => n2095, B2 => 
                           n2758, C1 => n2091, C2 => n2886, ZN => n958);
   U704 : OAI222_X1 port map( A1 => n2179, A2 => n3141, B1 => n2175, B2 => 
                           n2501, C1 => n2171, C2 => n2437, ZN => n907);
   U705 : OAI222_X1 port map( A1 => n2099, A2 => n2693, B1 => n2095, B2 => 
                           n2757, C1 => n2091, C2 => n2885, ZN => n923);
   U706 : OAI222_X1 port map( A1 => n3172, A2 => n2049, B1 => n2532, B2 => 
                           n2045, C1 => n2468, C2 => n2041, ZN => n1919);
   U707 : OAI222_X1 port map( A1 => n2724, A2 => n1969, B1 => n2788, B2 => 
                           n1965, C1 => n2916, C2 => n1961, ZN => n1925);
   U708 : OAI222_X1 port map( A1 => n3171, A2 => n2049, B1 => n2531, B2 => 
                           n2045, C1 => n2467, C2 => n2041, ZN => n1904);
   U709 : OAI222_X1 port map( A1 => n2723, A2 => n1969, B1 => n2787, B2 => 
                           n1965, C1 => n2915, C2 => n1961, ZN => n1908);
   U710 : OAI222_X1 port map( A1 => n3170, A2 => n2049, B1 => n2530, B2 => 
                           n2045, C1 => n2466, C2 => n2041, ZN => n1889);
   U711 : OAI222_X1 port map( A1 => n2722, A2 => n1969, B1 => n2786, B2 => 
                           n1965, C1 => n2914, C2 => n1961, ZN => n1893);
   U712 : OAI222_X1 port map( A1 => n3169, A2 => n2049, B1 => n2529, B2 => 
                           n2045, C1 => n2465, C2 => n2041, ZN => n1874);
   U713 : OAI222_X1 port map( A1 => n2721, A2 => n1969, B1 => n2785, B2 => 
                           n1965, C1 => n2913, C2 => n1961, ZN => n1878);
   U714 : OAI222_X1 port map( A1 => n3168, A2 => n2049, B1 => n2528, B2 => 
                           n2045, C1 => n2464, C2 => n2041, ZN => n1859);
   U715 : OAI222_X1 port map( A1 => n2720, A2 => n1969, B1 => n2784, B2 => 
                           n1965, C1 => n2912, C2 => n1961, ZN => n1863);
   U716 : OAI222_X1 port map( A1 => n3167, A2 => n2049, B1 => n2527, B2 => 
                           n2045, C1 => n2463, C2 => n2041, ZN => n1844);
   U717 : OAI222_X1 port map( A1 => n2719, A2 => n1969, B1 => n2783, B2 => 
                           n1965, C1 => n2911, C2 => n1961, ZN => n1848);
   U718 : OAI222_X1 port map( A1 => n3166, A2 => n2049, B1 => n2526, B2 => 
                           n2045, C1 => n2462, C2 => n2041, ZN => n1829);
   U719 : OAI222_X1 port map( A1 => n2718, A2 => n1969, B1 => n2782, B2 => 
                           n1965, C1 => n2910, C2 => n1961, ZN => n1833);
   U720 : OAI222_X1 port map( A1 => n3165, A2 => n2049, B1 => n2525, B2 => 
                           n2045, C1 => n2461, C2 => n2041, ZN => n1814);
   U721 : OAI222_X1 port map( A1 => n2717, A2 => n1969, B1 => n2781, B2 => 
                           n1965, C1 => n2909, C2 => n1961, ZN => n1818);
   U722 : OAI222_X1 port map( A1 => n3164, A2 => n2049, B1 => n2524, B2 => 
                           n2045, C1 => n2460, C2 => n2041, ZN => n1799);
   U723 : OAI222_X1 port map( A1 => n2716, A2 => n1969, B1 => n2780, B2 => 
                           n1965, C1 => n2908, C2 => n1961, ZN => n1803);
   U724 : OAI222_X1 port map( A1 => n3163, A2 => n2049, B1 => n2523, B2 => 
                           n2045, C1 => n2459, C2 => n2041, ZN => n1784);
   U725 : OAI222_X1 port map( A1 => n2715, A2 => n1969, B1 => n2779, B2 => 
                           n1965, C1 => n2907, C2 => n1961, ZN => n1788);
   U726 : OAI222_X1 port map( A1 => n3162, A2 => n2049, B1 => n2522, B2 => 
                           n2045, C1 => n2458, C2 => n2041, ZN => n1769);
   U727 : OAI222_X1 port map( A1 => n2714, A2 => n1969, B1 => n2778, B2 => 
                           n1965, C1 => n2906, C2 => n1961, ZN => n1773);
   U728 : OAI222_X1 port map( A1 => n3161, A2 => n2049, B1 => n2521, B2 => 
                           n2045, C1 => n2457, C2 => n2041, ZN => n1754);
   U729 : OAI222_X1 port map( A1 => n2713, A2 => n1969, B1 => n2777, B2 => 
                           n1965, C1 => n2905, C2 => n1961, ZN => n1758);
   U730 : OAI222_X1 port map( A1 => n3160, A2 => n2050, B1 => n2520, B2 => 
                           n2046, C1 => n2456, C2 => n2042, ZN => n1739);
   U731 : OAI222_X1 port map( A1 => n2712, A2 => n1970, B1 => n2776, B2 => 
                           n1966, C1 => n2904, C2 => n1962, ZN => n1743);
   U732 : OAI222_X1 port map( A1 => n3159, A2 => n2050, B1 => n2519, B2 => 
                           n2046, C1 => n2455, C2 => n2042, ZN => n1724);
   U733 : OAI222_X1 port map( A1 => n2711, A2 => n1970, B1 => n2775, B2 => 
                           n1966, C1 => n2903, C2 => n1962, ZN => n1728);
   U734 : OAI222_X1 port map( A1 => n3158, A2 => n2050, B1 => n2518, B2 => 
                           n2046, C1 => n2454, C2 => n2042, ZN => n1709);
   U735 : OAI222_X1 port map( A1 => n2710, A2 => n1970, B1 => n2774, B2 => 
                           n1966, C1 => n2902, C2 => n1962, ZN => n1713);
   U736 : OAI222_X1 port map( A1 => n3157, A2 => n2050, B1 => n2517, B2 => 
                           n2046, C1 => n2453, C2 => n2042, ZN => n1694);
   U737 : OAI222_X1 port map( A1 => n2709, A2 => n1970, B1 => n2773, B2 => 
                           n1966, C1 => n2901, C2 => n1962, ZN => n1698);
   U738 : OAI222_X1 port map( A1 => n3156, A2 => n2050, B1 => n2516, B2 => 
                           n2046, C1 => n2452, C2 => n2042, ZN => n1679);
   U739 : OAI222_X1 port map( A1 => n2708, A2 => n1970, B1 => n2772, B2 => 
                           n1966, C1 => n2900, C2 => n1962, ZN => n1683);
   U740 : OAI222_X1 port map( A1 => n3155, A2 => n2050, B1 => n2515, B2 => 
                           n2046, C1 => n2451, C2 => n2042, ZN => n1664);
   U741 : OAI222_X1 port map( A1 => n2707, A2 => n1970, B1 => n2771, B2 => 
                           n1966, C1 => n2899, C2 => n1962, ZN => n1668);
   U742 : OAI222_X1 port map( A1 => n3154, A2 => n2050, B1 => n2514, B2 => 
                           n2046, C1 => n2450, C2 => n2042, ZN => n1649);
   U743 : OAI222_X1 port map( A1 => n2706, A2 => n1970, B1 => n2770, B2 => 
                           n1966, C1 => n2898, C2 => n1962, ZN => n1653);
   U744 : OAI222_X1 port map( A1 => n3153, A2 => n2050, B1 => n2513, B2 => 
                           n2046, C1 => n2449, C2 => n2042, ZN => n1634);
   U745 : OAI222_X1 port map( A1 => n2705, A2 => n1970, B1 => n2769, B2 => 
                           n1966, C1 => n2897, C2 => n1962, ZN => n1638);
   U746 : OAI222_X1 port map( A1 => n3152, A2 => n2050, B1 => n2512, B2 => 
                           n2046, C1 => n2448, C2 => n2042, ZN => n1619);
   U747 : OAI222_X1 port map( A1 => n2704, A2 => n1970, B1 => n2768, B2 => 
                           n1966, C1 => n2896, C2 => n1962, ZN => n1623);
   U748 : OAI222_X1 port map( A1 => n3151, A2 => n2050, B1 => n2511, B2 => 
                           n2046, C1 => n2447, C2 => n2042, ZN => n1604);
   U749 : OAI222_X1 port map( A1 => n2703, A2 => n1970, B1 => n2767, B2 => 
                           n1966, C1 => n2895, C2 => n1962, ZN => n1608);
   U750 : OAI222_X1 port map( A1 => n3150, A2 => n2050, B1 => n2510, B2 => 
                           n2046, C1 => n2446, C2 => n2042, ZN => n1589);
   U751 : OAI222_X1 port map( A1 => n2702, A2 => n1970, B1 => n2766, B2 => 
                           n1966, C1 => n2894, C2 => n1962, ZN => n1593);
   U752 : OAI222_X1 port map( A1 => n3149, A2 => n2050, B1 => n2509, B2 => 
                           n2046, C1 => n2445, C2 => n2042, ZN => n1574);
   U753 : OAI222_X1 port map( A1 => n2701, A2 => n1970, B1 => n2765, B2 => 
                           n1966, C1 => n2893, C2 => n1962, ZN => n1578);
   U754 : OAI222_X1 port map( A1 => n3148, A2 => n2051, B1 => n2508, B2 => 
                           n2047, C1 => n2444, C2 => n2043, ZN => n1559);
   U755 : OAI222_X1 port map( A1 => n2700, A2 => n1971, B1 => n2764, B2 => 
                           n1967, C1 => n2892, C2 => n1963, ZN => n1563);
   U756 : OAI222_X1 port map( A1 => n3147, A2 => n2051, B1 => n2507, B2 => 
                           n2047, C1 => n2443, C2 => n2043, ZN => n1544);
   U757 : OAI222_X1 port map( A1 => n2699, A2 => n1971, B1 => n2763, B2 => 
                           n1967, C1 => n2891, C2 => n1963, ZN => n1548);
   U758 : OAI222_X1 port map( A1 => n3146, A2 => n2051, B1 => n2506, B2 => 
                           n2047, C1 => n2442, C2 => n2043, ZN => n1529);
   U759 : OAI222_X1 port map( A1 => n2698, A2 => n1971, B1 => n2762, B2 => 
                           n1967, C1 => n2890, C2 => n1963, ZN => n1533);
   U760 : OAI222_X1 port map( A1 => n3145, A2 => n2051, B1 => n2505, B2 => 
                           n2047, C1 => n2441, C2 => n2043, ZN => n1514);
   U761 : OAI222_X1 port map( A1 => n2697, A2 => n1971, B1 => n2761, B2 => 
                           n1967, C1 => n2889, C2 => n1963, ZN => n1518);
   U762 : OAI222_X1 port map( A1 => n3144, A2 => n2051, B1 => n2504, B2 => 
                           n2047, C1 => n2440, C2 => n2043, ZN => n1499);
   U763 : OAI222_X1 port map( A1 => n2696, A2 => n1971, B1 => n2760, B2 => 
                           n1967, C1 => n2888, C2 => n1963, ZN => n1503);
   U764 : OAI222_X1 port map( A1 => n3143, A2 => n2051, B1 => n2503, B2 => 
                           n2047, C1 => n2439, C2 => n2043, ZN => n1484);
   U765 : OAI222_X1 port map( A1 => n2695, A2 => n1971, B1 => n2759, B2 => 
                           n1967, C1 => n2887, C2 => n1963, ZN => n1488);
   U766 : OAI222_X1 port map( A1 => n3142, A2 => n2051, B1 => n2502, B2 => 
                           n2047, C1 => n2438, C2 => n2043, ZN => n1469);
   U767 : OAI222_X1 port map( A1 => n2694, A2 => n1971, B1 => n2758, B2 => 
                           n1967, C1 => n2886, C2 => n1963, ZN => n1473);
   U768 : OAI222_X1 port map( A1 => n3141, A2 => n2051, B1 => n2501, B2 => 
                           n2047, C1 => n2437, C2 => n2043, ZN => n1422);
   U769 : OAI222_X1 port map( A1 => n2693, A2 => n1971, B1 => n2757, B2 => 
                           n1967, C1 => n2885, C2 => n1963, ZN => n1438);
   U770 : OAI222_X1 port map( A1 => n2165, A2 => n3044, B1 => n2161, B2 => 
                           n2404, C1 => n2157, C2 => n2980, ZN => n1403);
   U771 : OAI222_X1 port map( A1 => n2085, A2 => n2500, B1 => n2081, B2 => 
                           n3204, C1 => n2077, C2 => n3140, ZN => n1409);
   U772 : OAI222_X1 port map( A1 => n2165, A2 => n3043, B1 => n2161, B2 => 
                           n2403, C1 => n2157, C2 => n2979, ZN => n1388);
   U773 : OAI222_X1 port map( A1 => n2085, A2 => n2499, B1 => n2081, B2 => 
                           n3203, C1 => n2077, C2 => n3139, ZN => n1392);
   U774 : OAI222_X1 port map( A1 => n2165, A2 => n3042, B1 => n2161, B2 => 
                           n2402, C1 => n2157, C2 => n2978, ZN => n1373);
   U775 : OAI222_X1 port map( A1 => n2085, A2 => n2498, B1 => n2081, B2 => 
                           n3202, C1 => n2077, C2 => n3138, ZN => n1377);
   U776 : OAI222_X1 port map( A1 => n2165, A2 => n3041, B1 => n2161, B2 => 
                           n2401, C1 => n2157, C2 => n2977, ZN => n1358);
   U777 : OAI222_X1 port map( A1 => n2085, A2 => n2497, B1 => n2081, B2 => 
                           n3201, C1 => n2077, C2 => n3137, ZN => n1362);
   U778 : OAI222_X1 port map( A1 => n2165, A2 => n3040, B1 => n2161, B2 => 
                           n2400, C1 => n2157, C2 => n2976, ZN => n1343);
   U779 : OAI222_X1 port map( A1 => n2085, A2 => n2496, B1 => n2081, B2 => 
                           n3200, C1 => n2077, C2 => n3136, ZN => n1347);
   U780 : OAI222_X1 port map( A1 => n2165, A2 => n3039, B1 => n2161, B2 => 
                           n2399, C1 => n2157, C2 => n2975, ZN => n1328);
   U781 : OAI222_X1 port map( A1 => n2085, A2 => n2495, B1 => n2081, B2 => 
                           n3199, C1 => n2077, C2 => n3135, ZN => n1332);
   U782 : OAI222_X1 port map( A1 => n2165, A2 => n3038, B1 => n2161, B2 => 
                           n2398, C1 => n2157, C2 => n2974, ZN => n1313);
   U783 : OAI222_X1 port map( A1 => n2085, A2 => n2494, B1 => n2081, B2 => 
                           n3198, C1 => n2077, C2 => n3134, ZN => n1317);
   U784 : OAI222_X1 port map( A1 => n2165, A2 => n3037, B1 => n2161, B2 => 
                           n2397, C1 => n2157, C2 => n2973, ZN => n1298);
   U785 : OAI222_X1 port map( A1 => n2085, A2 => n2493, B1 => n2081, B2 => 
                           n3197, C1 => n2077, C2 => n3133, ZN => n1302);
   U786 : OAI222_X1 port map( A1 => n2165, A2 => n3036, B1 => n2161, B2 => 
                           n2396, C1 => n2157, C2 => n2972, ZN => n1283);
   U787 : OAI222_X1 port map( A1 => n2085, A2 => n2492, B1 => n2081, B2 => 
                           n3196, C1 => n2077, C2 => n3132, ZN => n1287);
   U788 : OAI222_X1 port map( A1 => n2165, A2 => n3035, B1 => n2161, B2 => 
                           n2395, C1 => n2157, C2 => n2971, ZN => n1268);
   U789 : OAI222_X1 port map( A1 => n2085, A2 => n2491, B1 => n2081, B2 => 
                           n3195, C1 => n2077, C2 => n3131, ZN => n1272);
   U790 : OAI222_X1 port map( A1 => n2165, A2 => n3034, B1 => n2161, B2 => 
                           n2394, C1 => n2157, C2 => n2970, ZN => n1253);
   U791 : OAI222_X1 port map( A1 => n2085, A2 => n2490, B1 => n2081, B2 => 
                           n3194, C1 => n2077, C2 => n3130, ZN => n1257);
   U792 : OAI222_X1 port map( A1 => n2165, A2 => n3033, B1 => n2161, B2 => 
                           n2393, C1 => n2157, C2 => n2969, ZN => n1238);
   U793 : OAI222_X1 port map( A1 => n2085, A2 => n2489, B1 => n2081, B2 => 
                           n3193, C1 => n2077, C2 => n3129, ZN => n1242);
   U794 : OAI222_X1 port map( A1 => n2166, A2 => n3032, B1 => n2162, B2 => 
                           n2392, C1 => n2158, C2 => n2968, ZN => n1223);
   U795 : OAI222_X1 port map( A1 => n2086, A2 => n2488, B1 => n2082, B2 => 
                           n3192, C1 => n2078, C2 => n3128, ZN => n1227);
   U796 : OAI222_X1 port map( A1 => n2166, A2 => n3031, B1 => n2162, B2 => 
                           n2391, C1 => n2158, C2 => n2967, ZN => n1208);
   U797 : OAI222_X1 port map( A1 => n2086, A2 => n2487, B1 => n2082, B2 => 
                           n3191, C1 => n2078, C2 => n3127, ZN => n1212);
   U798 : OAI222_X1 port map( A1 => n2166, A2 => n3030, B1 => n2162, B2 => 
                           n2390, C1 => n2158, C2 => n2966, ZN => n1193);
   U799 : OAI222_X1 port map( A1 => n2086, A2 => n2486, B1 => n2082, B2 => 
                           n3190, C1 => n2078, C2 => n3126, ZN => n1197);
   U800 : OAI222_X1 port map( A1 => n2166, A2 => n3029, B1 => n2162, B2 => 
                           n2389, C1 => n2158, C2 => n2965, ZN => n1178);
   U801 : OAI222_X1 port map( A1 => n2086, A2 => n2485, B1 => n2082, B2 => 
                           n3189, C1 => n2078, C2 => n3125, ZN => n1182);
   U802 : OAI222_X1 port map( A1 => n2166, A2 => n3028, B1 => n2162, B2 => 
                           n2388, C1 => n2158, C2 => n2964, ZN => n1163);
   U803 : OAI222_X1 port map( A1 => n2086, A2 => n2484, B1 => n2082, B2 => 
                           n3188, C1 => n2078, C2 => n3124, ZN => n1167);
   U804 : OAI222_X1 port map( A1 => n2166, A2 => n3027, B1 => n2162, B2 => 
                           n2387, C1 => n2158, C2 => n2963, ZN => n1148);
   U805 : OAI222_X1 port map( A1 => n2086, A2 => n2483, B1 => n2082, B2 => 
                           n3187, C1 => n2078, C2 => n3123, ZN => n1152);
   U806 : OAI222_X1 port map( A1 => n2166, A2 => n3026, B1 => n2162, B2 => 
                           n2386, C1 => n2158, C2 => n2962, ZN => n1133);
   U807 : OAI222_X1 port map( A1 => n2086, A2 => n2482, B1 => n2082, B2 => 
                           n3186, C1 => n2078, C2 => n3122, ZN => n1137);
   U808 : OAI222_X1 port map( A1 => n2166, A2 => n3025, B1 => n2162, B2 => 
                           n2385, C1 => n2158, C2 => n2961, ZN => n1118);
   U809 : OAI222_X1 port map( A1 => n2086, A2 => n2481, B1 => n2082, B2 => 
                           n3185, C1 => n2078, C2 => n3121, ZN => n1122);
   U810 : OAI222_X1 port map( A1 => n2166, A2 => n3024, B1 => n2162, B2 => 
                           n2384, C1 => n2158, C2 => n2960, ZN => n1103);
   U811 : OAI222_X1 port map( A1 => n2086, A2 => n2480, B1 => n2082, B2 => 
                           n3184, C1 => n2078, C2 => n3120, ZN => n1107);
   U812 : OAI222_X1 port map( A1 => n2166, A2 => n3023, B1 => n2162, B2 => 
                           n2383, C1 => n2158, C2 => n2959, ZN => n1088);
   U813 : OAI222_X1 port map( A1 => n2086, A2 => n2479, B1 => n2082, B2 => 
                           n3183, C1 => n2078, C2 => n3119, ZN => n1092);
   U814 : OAI222_X1 port map( A1 => n2166, A2 => n3022, B1 => n2162, B2 => 
                           n2382, C1 => n2158, C2 => n2958, ZN => n1073);
   U815 : OAI222_X1 port map( A1 => n2086, A2 => n2478, B1 => n2082, B2 => 
                           n3182, C1 => n2078, C2 => n3118, ZN => n1077);
   U816 : OAI222_X1 port map( A1 => n2166, A2 => n3021, B1 => n2162, B2 => 
                           n2381, C1 => n2158, C2 => n2957, ZN => n1058);
   U817 : OAI222_X1 port map( A1 => n2086, A2 => n2477, B1 => n2082, B2 => 
                           n3181, C1 => n2078, C2 => n3117, ZN => n1062);
   U818 : OAI222_X1 port map( A1 => n2167, A2 => n3020, B1 => n2163, B2 => 
                           n2380, C1 => n2159, C2 => n2956, ZN => n1043);
   U819 : OAI222_X1 port map( A1 => n2087, A2 => n2476, B1 => n2083, B2 => 
                           n3180, C1 => n2079, C2 => n3116, ZN => n1047);
   U820 : OAI222_X1 port map( A1 => n2167, A2 => n3019, B1 => n2163, B2 => 
                           n2379, C1 => n2159, C2 => n2955, ZN => n1028);
   U821 : OAI222_X1 port map( A1 => n2087, A2 => n2475, B1 => n2083, B2 => 
                           n3179, C1 => n2079, C2 => n3115, ZN => n1032);
   U822 : OAI222_X1 port map( A1 => n2167, A2 => n3018, B1 => n2163, B2 => 
                           n2378, C1 => n2159, C2 => n2954, ZN => n1013);
   U823 : OAI222_X1 port map( A1 => n2087, A2 => n2474, B1 => n2083, B2 => 
                           n3178, C1 => n2079, C2 => n3114, ZN => n1017);
   U824 : OAI222_X1 port map( A1 => n2167, A2 => n3017, B1 => n2163, B2 => 
                           n2377, C1 => n2159, C2 => n2953, ZN => n998);
   U825 : OAI222_X1 port map( A1 => n2087, A2 => n2473, B1 => n2083, B2 => 
                           n3177, C1 => n2079, C2 => n3113, ZN => n1002);
   U826 : OAI222_X1 port map( A1 => n2167, A2 => n3016, B1 => n2163, B2 => 
                           n2376, C1 => n2159, C2 => n2952, ZN => n983);
   U827 : OAI222_X1 port map( A1 => n2087, A2 => n2472, B1 => n2083, B2 => 
                           n3176, C1 => n2079, C2 => n3112, ZN => n987);
   U828 : OAI222_X1 port map( A1 => n2167, A2 => n3015, B1 => n2163, B2 => 
                           n2375, C1 => n2159, C2 => n2951, ZN => n968);
   U829 : OAI222_X1 port map( A1 => n2087, A2 => n2471, B1 => n2083, B2 => 
                           n3175, C1 => n2079, C2 => n3111, ZN => n972);
   U830 : OAI222_X1 port map( A1 => n2167, A2 => n3014, B1 => n2163, B2 => 
                           n2374, C1 => n2159, C2 => n2950, ZN => n953);
   U831 : OAI222_X1 port map( A1 => n2087, A2 => n2470, B1 => n2083, B2 => 
                           n3174, C1 => n2079, C2 => n3110, ZN => n957);
   U832 : OAI222_X1 port map( A1 => n2167, A2 => n3013, B1 => n2163, B2 => 
                           n2373, C1 => n2159, C2 => n2949, ZN => n906);
   U833 : OAI222_X1 port map( A1 => n2087, A2 => n2469, B1 => n2083, B2 => 
                           n3173, C1 => n2079, C2 => n3109, ZN => n922);
   U834 : OAI222_X1 port map( A1 => n3044, A2 => n2037, B1 => n2404, B2 => 
                           n2033, C1 => n2980, C2 => n2029, ZN => n1918);
   U835 : OAI222_X1 port map( A1 => n2500, A2 => n1957, B1 => n3204, B2 => 
                           n1953, C1 => n3140, C2 => n1949, ZN => n1924);
   U836 : OAI222_X1 port map( A1 => n3043, A2 => n2037, B1 => n2403, B2 => 
                           n2033, C1 => n2979, C2 => n2029, ZN => n1903);
   U837 : OAI222_X1 port map( A1 => n2499, A2 => n1957, B1 => n3203, B2 => 
                           n1953, C1 => n3139, C2 => n1949, ZN => n1907);
   U838 : OAI222_X1 port map( A1 => n3042, A2 => n2037, B1 => n2402, B2 => 
                           n2033, C1 => n2978, C2 => n2029, ZN => n1888);
   U839 : OAI222_X1 port map( A1 => n2498, A2 => n1957, B1 => n3202, B2 => 
                           n1953, C1 => n3138, C2 => n1949, ZN => n1892);
   U840 : OAI222_X1 port map( A1 => n3041, A2 => n2037, B1 => n2401, B2 => 
                           n2033, C1 => n2977, C2 => n2029, ZN => n1873);
   U841 : OAI222_X1 port map( A1 => n2497, A2 => n1957, B1 => n3201, B2 => 
                           n1953, C1 => n3137, C2 => n1949, ZN => n1877);
   U842 : OAI222_X1 port map( A1 => n3040, A2 => n2037, B1 => n2400, B2 => 
                           n2033, C1 => n2976, C2 => n2029, ZN => n1858);
   U843 : OAI222_X1 port map( A1 => n2496, A2 => n1957, B1 => n3200, B2 => 
                           n1953, C1 => n3136, C2 => n1949, ZN => n1862);
   U844 : OAI222_X1 port map( A1 => n3039, A2 => n2037, B1 => n2399, B2 => 
                           n2033, C1 => n2975, C2 => n2029, ZN => n1843);
   U845 : OAI222_X1 port map( A1 => n2495, A2 => n1957, B1 => n3199, B2 => 
                           n1953, C1 => n3135, C2 => n1949, ZN => n1847);
   U846 : OAI222_X1 port map( A1 => n3038, A2 => n2037, B1 => n2398, B2 => 
                           n2033, C1 => n2974, C2 => n2029, ZN => n1828);
   U847 : OAI222_X1 port map( A1 => n2494, A2 => n1957, B1 => n3198, B2 => 
                           n1953, C1 => n3134, C2 => n1949, ZN => n1832);
   U848 : OAI222_X1 port map( A1 => n3037, A2 => n2037, B1 => n2397, B2 => 
                           n2033, C1 => n2973, C2 => n2029, ZN => n1813);
   U849 : OAI222_X1 port map( A1 => n2493, A2 => n1957, B1 => n3197, B2 => 
                           n1953, C1 => n3133, C2 => n1949, ZN => n1817);
   U850 : OAI222_X1 port map( A1 => n3036, A2 => n2037, B1 => n2396, B2 => 
                           n2033, C1 => n2972, C2 => n2029, ZN => n1798);
   U851 : OAI222_X1 port map( A1 => n2492, A2 => n1957, B1 => n3196, B2 => 
                           n1953, C1 => n3132, C2 => n1949, ZN => n1802);
   U852 : OAI222_X1 port map( A1 => n3035, A2 => n2037, B1 => n2395, B2 => 
                           n2033, C1 => n2971, C2 => n2029, ZN => n1783);
   U853 : OAI222_X1 port map( A1 => n2491, A2 => n1957, B1 => n3195, B2 => 
                           n1953, C1 => n3131, C2 => n1949, ZN => n1787);
   U854 : OAI222_X1 port map( A1 => n3034, A2 => n2037, B1 => n2394, B2 => 
                           n2033, C1 => n2970, C2 => n2029, ZN => n1768);
   U855 : OAI222_X1 port map( A1 => n2490, A2 => n1957, B1 => n3194, B2 => 
                           n1953, C1 => n3130, C2 => n1949, ZN => n1772);
   U856 : OAI222_X1 port map( A1 => n3033, A2 => n2037, B1 => n2393, B2 => 
                           n2033, C1 => n2969, C2 => n2029, ZN => n1753);
   U857 : OAI222_X1 port map( A1 => n2489, A2 => n1957, B1 => n3193, B2 => 
                           n1953, C1 => n3129, C2 => n1949, ZN => n1757);
   U858 : OAI222_X1 port map( A1 => n3032, A2 => n2038, B1 => n2392, B2 => 
                           n2034, C1 => n2968, C2 => n2030, ZN => n1738);
   U859 : OAI222_X1 port map( A1 => n2488, A2 => n1958, B1 => n3192, B2 => 
                           n1954, C1 => n3128, C2 => n1950, ZN => n1742);
   U860 : OAI222_X1 port map( A1 => n3031, A2 => n2038, B1 => n2391, B2 => 
                           n2034, C1 => n2967, C2 => n2030, ZN => n1723);
   U861 : OAI222_X1 port map( A1 => n2487, A2 => n1958, B1 => n3191, B2 => 
                           n1954, C1 => n3127, C2 => n1950, ZN => n1727);
   U862 : OAI222_X1 port map( A1 => n3030, A2 => n2038, B1 => n2390, B2 => 
                           n2034, C1 => n2966, C2 => n2030, ZN => n1708);
   U863 : OAI222_X1 port map( A1 => n2486, A2 => n1958, B1 => n3190, B2 => 
                           n1954, C1 => n3126, C2 => n1950, ZN => n1712);
   U864 : OAI222_X1 port map( A1 => n3029, A2 => n2038, B1 => n2389, B2 => 
                           n2034, C1 => n2965, C2 => n2030, ZN => n1693);
   U865 : OAI222_X1 port map( A1 => n2485, A2 => n1958, B1 => n3189, B2 => 
                           n1954, C1 => n3125, C2 => n1950, ZN => n1697);
   U866 : OAI222_X1 port map( A1 => n3028, A2 => n2038, B1 => n2388, B2 => 
                           n2034, C1 => n2964, C2 => n2030, ZN => n1678);
   U867 : OAI222_X1 port map( A1 => n2484, A2 => n1958, B1 => n3188, B2 => 
                           n1954, C1 => n3124, C2 => n1950, ZN => n1682);
   U868 : OAI222_X1 port map( A1 => n3027, A2 => n2038, B1 => n2387, B2 => 
                           n2034, C1 => n2963, C2 => n2030, ZN => n1663);
   U869 : OAI222_X1 port map( A1 => n2483, A2 => n1958, B1 => n3187, B2 => 
                           n1954, C1 => n3123, C2 => n1950, ZN => n1667);
   U870 : OAI222_X1 port map( A1 => n3026, A2 => n2038, B1 => n2386, B2 => 
                           n2034, C1 => n2962, C2 => n2030, ZN => n1648);
   U871 : OAI222_X1 port map( A1 => n2482, A2 => n1958, B1 => n3186, B2 => 
                           n1954, C1 => n3122, C2 => n1950, ZN => n1652);
   U872 : OAI222_X1 port map( A1 => n3025, A2 => n2038, B1 => n2385, B2 => 
                           n2034, C1 => n2961, C2 => n2030, ZN => n1633);
   U873 : OAI222_X1 port map( A1 => n2481, A2 => n1958, B1 => n3185, B2 => 
                           n1954, C1 => n3121, C2 => n1950, ZN => n1637);
   U874 : OAI222_X1 port map( A1 => n3024, A2 => n2038, B1 => n2384, B2 => 
                           n2034, C1 => n2960, C2 => n2030, ZN => n1618);
   U875 : OAI222_X1 port map( A1 => n2480, A2 => n1958, B1 => n3184, B2 => 
                           n1954, C1 => n3120, C2 => n1950, ZN => n1622);
   U876 : OAI222_X1 port map( A1 => n3023, A2 => n2038, B1 => n2383, B2 => 
                           n2034, C1 => n2959, C2 => n2030, ZN => n1603);
   U877 : OAI222_X1 port map( A1 => n2479, A2 => n1958, B1 => n3183, B2 => 
                           n1954, C1 => n3119, C2 => n1950, ZN => n1607);
   U878 : OAI222_X1 port map( A1 => n3022, A2 => n2038, B1 => n2382, B2 => 
                           n2034, C1 => n2958, C2 => n2030, ZN => n1588);
   U879 : OAI222_X1 port map( A1 => n2478, A2 => n1958, B1 => n3182, B2 => 
                           n1954, C1 => n3118, C2 => n1950, ZN => n1592);
   U880 : OAI222_X1 port map( A1 => n3021, A2 => n2038, B1 => n2381, B2 => 
                           n2034, C1 => n2957, C2 => n2030, ZN => n1573);
   U881 : OAI222_X1 port map( A1 => n2477, A2 => n1958, B1 => n3181, B2 => 
                           n1954, C1 => n3117, C2 => n1950, ZN => n1577);
   U882 : OAI222_X1 port map( A1 => n3020, A2 => n2039, B1 => n2380, B2 => 
                           n2035, C1 => n2956, C2 => n2031, ZN => n1558);
   U883 : OAI222_X1 port map( A1 => n2476, A2 => n1959, B1 => n3180, B2 => 
                           n1955, C1 => n3116, C2 => n1951, ZN => n1562);
   U884 : OAI222_X1 port map( A1 => n3019, A2 => n2039, B1 => n2379, B2 => 
                           n2035, C1 => n2955, C2 => n2031, ZN => n1543);
   U885 : OAI222_X1 port map( A1 => n2475, A2 => n1959, B1 => n3179, B2 => 
                           n1955, C1 => n3115, C2 => n1951, ZN => n1547);
   U886 : OAI222_X1 port map( A1 => n3018, A2 => n2039, B1 => n2378, B2 => 
                           n2035, C1 => n2954, C2 => n2031, ZN => n1528);
   U887 : OAI222_X1 port map( A1 => n2474, A2 => n1959, B1 => n3178, B2 => 
                           n1955, C1 => n3114, C2 => n1951, ZN => n1532);
   U888 : OAI222_X1 port map( A1 => n3017, A2 => n2039, B1 => n2377, B2 => 
                           n2035, C1 => n2953, C2 => n2031, ZN => n1513);
   U889 : OAI222_X1 port map( A1 => n2473, A2 => n1959, B1 => n3177, B2 => 
                           n1955, C1 => n3113, C2 => n1951, ZN => n1517);
   U890 : OAI222_X1 port map( A1 => n3016, A2 => n2039, B1 => n2376, B2 => 
                           n2035, C1 => n2952, C2 => n2031, ZN => n1498);
   U891 : OAI222_X1 port map( A1 => n2472, A2 => n1959, B1 => n3176, B2 => 
                           n1955, C1 => n3112, C2 => n1951, ZN => n1502);
   U892 : OAI222_X1 port map( A1 => n3015, A2 => n2039, B1 => n2375, B2 => 
                           n2035, C1 => n2951, C2 => n2031, ZN => n1483);
   U893 : OAI222_X1 port map( A1 => n2471, A2 => n1959, B1 => n3175, B2 => 
                           n1955, C1 => n3111, C2 => n1951, ZN => n1487);
   U894 : OAI222_X1 port map( A1 => n3014, A2 => n2039, B1 => n2374, B2 => 
                           n2035, C1 => n2950, C2 => n2031, ZN => n1468);
   U895 : OAI222_X1 port map( A1 => n2470, A2 => n1959, B1 => n3174, B2 => 
                           n1955, C1 => n3110, C2 => n1951, ZN => n1472);
   U896 : OAI222_X1 port map( A1 => n3013, A2 => n2039, B1 => n2373, B2 => 
                           n2035, C1 => n2949, C2 => n2031, ZN => n1421);
   U897 : OAI222_X1 port map( A1 => n2469, A2 => n1959, B1 => n3173, B2 => 
                           n1955, C1 => n3109, C2 => n1951, ZN => n1437);
   U898 : AND3_X1 port map( A1 => n3219, A2 => n3218, A3 => ADD_RD2(2), ZN => 
                           n1934);
   U899 : AOI21_X1 port map( B1 => n1401, B2 => n1402, A => n1942, ZN => N291);
   U900 : NOR4_X1 port map( A1 => n1409, A2 => n1410, A3 => n1411, A4 => n1412,
                           ZN => n1401);
   U901 : NOR4_X1 port map( A1 => n1403, A2 => n1404, A3 => n1405, A4 => n1406,
                           ZN => n1402);
   U902 : OAI221_X1 port map( B1 => n2153, B2 => n2948, C1 => n2149, C2 => 
                           n2884, A => n1413, ZN => n1412);
   U903 : AOI21_X1 port map( B1 => n1386, B2 => n1387, A => n1942, ZN => N292);
   U904 : NOR4_X1 port map( A1 => n1392, A2 => n1393, A3 => n1394, A4 => n1395,
                           ZN => n1386);
   U905 : NOR4_X1 port map( A1 => n1388, A2 => n1389, A3 => n1390, A4 => n1391,
                           ZN => n1387);
   U906 : OAI221_X1 port map( B1 => n2153, B2 => n2947, C1 => n2149, C2 => 
                           n2883, A => n1396, ZN => n1395);
   U907 : AOI21_X1 port map( B1 => n1371, B2 => n1372, A => n1942, ZN => N293);
   U908 : NOR4_X1 port map( A1 => n1377, A2 => n1378, A3 => n1379, A4 => n1380,
                           ZN => n1371);
   U909 : NOR4_X1 port map( A1 => n1373, A2 => n1374, A3 => n1375, A4 => n1376,
                           ZN => n1372);
   U910 : OAI221_X1 port map( B1 => n2153, B2 => n2946, C1 => n2149, C2 => 
                           n2882, A => n1381, ZN => n1380);
   U911 : AOI21_X1 port map( B1 => n1356, B2 => n1357, A => n1942, ZN => N294);
   U912 : NOR4_X1 port map( A1 => n1362, A2 => n1363, A3 => n1364, A4 => n1365,
                           ZN => n1356);
   U913 : NOR4_X1 port map( A1 => n1358, A2 => n1359, A3 => n1360, A4 => n1361,
                           ZN => n1357);
   U914 : OAI221_X1 port map( B1 => n2153, B2 => n2945, C1 => n2149, C2 => 
                           n2881, A => n1366, ZN => n1365);
   U915 : AOI21_X1 port map( B1 => n1341, B2 => n1342, A => n1942, ZN => N295);
   U916 : NOR4_X1 port map( A1 => n1347, A2 => n1348, A3 => n1349, A4 => n1350,
                           ZN => n1341);
   U917 : NOR4_X1 port map( A1 => n1343, A2 => n1344, A3 => n1345, A4 => n1346,
                           ZN => n1342);
   U918 : OAI221_X1 port map( B1 => n2153, B2 => n2944, C1 => n2149, C2 => 
                           n2880, A => n1351, ZN => n1350);
   U919 : AOI21_X1 port map( B1 => n1326, B2 => n1327, A => n1942, ZN => N296);
   U920 : NOR4_X1 port map( A1 => n1332, A2 => n1333, A3 => n1334, A4 => n1335,
                           ZN => n1326);
   U921 : NOR4_X1 port map( A1 => n1328, A2 => n1329, A3 => n1330, A4 => n1331,
                           ZN => n1327);
   U922 : OAI221_X1 port map( B1 => n2153, B2 => n2943, C1 => n2149, C2 => 
                           n2879, A => n1336, ZN => n1335);
   U923 : AOI21_X1 port map( B1 => n1311, B2 => n1312, A => n1942, ZN => N297);
   U924 : NOR4_X1 port map( A1 => n1317, A2 => n1318, A3 => n1319, A4 => n1320,
                           ZN => n1311);
   U925 : NOR4_X1 port map( A1 => n1313, A2 => n1314, A3 => n1315, A4 => n1316,
                           ZN => n1312);
   U926 : OAI221_X1 port map( B1 => n2153, B2 => n2942, C1 => n2149, C2 => 
                           n2878, A => n1321, ZN => n1320);
   U927 : AOI21_X1 port map( B1 => n1296, B2 => n1297, A => n1942, ZN => N298);
   U928 : NOR4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1304, A4 => n1305,
                           ZN => n1296);
   U929 : NOR4_X1 port map( A1 => n1298, A2 => n1299, A3 => n1300, A4 => n1301,
                           ZN => n1297);
   U930 : OAI221_X1 port map( B1 => n2153, B2 => n2941, C1 => n2149, C2 => 
                           n2877, A => n1306, ZN => n1305);
   U931 : AOI21_X1 port map( B1 => n1281, B2 => n1282, A => n1942, ZN => N299);
   U932 : NOR4_X1 port map( A1 => n1287, A2 => n1288, A3 => n1289, A4 => n1290,
                           ZN => n1281);
   U933 : NOR4_X1 port map( A1 => n1283, A2 => n1284, A3 => n1285, A4 => n1286,
                           ZN => n1282);
   U934 : OAI221_X1 port map( B1 => n2153, B2 => n2940, C1 => n2149, C2 => 
                           n2876, A => n1291, ZN => n1290);
   U935 : AOI21_X1 port map( B1 => n1266, B2 => n1267, A => n1942, ZN => N300);
   U936 : NOR4_X1 port map( A1 => n1272, A2 => n1273, A3 => n1274, A4 => n1275,
                           ZN => n1266);
   U937 : NOR4_X1 port map( A1 => n1268, A2 => n1269, A3 => n1270, A4 => n1271,
                           ZN => n1267);
   U938 : OAI221_X1 port map( B1 => n2153, B2 => n2939, C1 => n2149, C2 => 
                           n2875, A => n1276, ZN => n1275);
   U939 : AOI21_X1 port map( B1 => n1251, B2 => n1252, A => n1942, ZN => N301);
   U940 : NOR4_X1 port map( A1 => n1257, A2 => n1258, A3 => n1259, A4 => n1260,
                           ZN => n1251);
   U941 : NOR4_X1 port map( A1 => n1253, A2 => n1254, A3 => n1255, A4 => n1256,
                           ZN => n1252);
   U942 : OAI221_X1 port map( B1 => n2153, B2 => n2938, C1 => n2149, C2 => 
                           n2874, A => n1261, ZN => n1260);
   U943 : AOI21_X1 port map( B1 => n1236, B2 => n1237, A => n1942, ZN => N302);
   U944 : NOR4_X1 port map( A1 => n1242, A2 => n1243, A3 => n1244, A4 => n1245,
                           ZN => n1236);
   U945 : NOR4_X1 port map( A1 => n1238, A2 => n1239, A3 => n1240, A4 => n1241,
                           ZN => n1237);
   U946 : OAI221_X1 port map( B1 => n2153, B2 => n2937, C1 => n2149, C2 => 
                           n2873, A => n1246, ZN => n1245);
   U947 : AOI21_X1 port map( B1 => n1221, B2 => n1222, A => n1943, ZN => N303);
   U948 : NOR4_X1 port map( A1 => n1227, A2 => n1228, A3 => n1229, A4 => n1230,
                           ZN => n1221);
   U949 : NOR4_X1 port map( A1 => n1223, A2 => n1224, A3 => n1225, A4 => n1226,
                           ZN => n1222);
   U950 : OAI221_X1 port map( B1 => n2154, B2 => n2936, C1 => n2150, C2 => 
                           n2872, A => n1231, ZN => n1230);
   U951 : AOI21_X1 port map( B1 => n1206, B2 => n1207, A => n1943, ZN => N304);
   U952 : NOR4_X1 port map( A1 => n1212, A2 => n1213, A3 => n1214, A4 => n1215,
                           ZN => n1206);
   U953 : NOR4_X1 port map( A1 => n1208, A2 => n1209, A3 => n1210, A4 => n1211,
                           ZN => n1207);
   U954 : OAI221_X1 port map( B1 => n2154, B2 => n2935, C1 => n2150, C2 => 
                           n2871, A => n1216, ZN => n1215);
   U955 : AOI21_X1 port map( B1 => n1191, B2 => n1192, A => n1943, ZN => N305);
   U956 : NOR4_X1 port map( A1 => n1197, A2 => n1198, A3 => n1199, A4 => n1200,
                           ZN => n1191);
   U957 : NOR4_X1 port map( A1 => n1193, A2 => n1194, A3 => n1195, A4 => n1196,
                           ZN => n1192);
   U958 : OAI221_X1 port map( B1 => n2154, B2 => n2934, C1 => n2150, C2 => 
                           n2870, A => n1201, ZN => n1200);
   U959 : AOI21_X1 port map( B1 => n1176, B2 => n1177, A => n1943, ZN => N306);
   U960 : NOR4_X1 port map( A1 => n1182, A2 => n1183, A3 => n1184, A4 => n1185,
                           ZN => n1176);
   U961 : NOR4_X1 port map( A1 => n1178, A2 => n1179, A3 => n1180, A4 => n1181,
                           ZN => n1177);
   U962 : OAI221_X1 port map( B1 => n2154, B2 => n2933, C1 => n2150, C2 => 
                           n2869, A => n1186, ZN => n1185);
   U963 : AOI21_X1 port map( B1 => n1161, B2 => n1162, A => n1943, ZN => N307);
   U964 : NOR4_X1 port map( A1 => n1167, A2 => n1168, A3 => n1169, A4 => n1170,
                           ZN => n1161);
   U965 : NOR4_X1 port map( A1 => n1163, A2 => n1164, A3 => n1165, A4 => n1166,
                           ZN => n1162);
   U966 : OAI221_X1 port map( B1 => n2154, B2 => n2932, C1 => n2150, C2 => 
                           n2868, A => n1171, ZN => n1170);
   U967 : AOI21_X1 port map( B1 => n1146, B2 => n1147, A => n1943, ZN => N308);
   U968 : NOR4_X1 port map( A1 => n1152, A2 => n1153, A3 => n1154, A4 => n1155,
                           ZN => n1146);
   U969 : NOR4_X1 port map( A1 => n1148, A2 => n1149, A3 => n1150, A4 => n1151,
                           ZN => n1147);
   U970 : OAI221_X1 port map( B1 => n2154, B2 => n2931, C1 => n2150, C2 => 
                           n2867, A => n1156, ZN => n1155);
   U971 : AOI21_X1 port map( B1 => n1131, B2 => n1132, A => n1943, ZN => N309);
   U972 : NOR4_X1 port map( A1 => n1137, A2 => n1138, A3 => n1139, A4 => n1140,
                           ZN => n1131);
   U973 : NOR4_X1 port map( A1 => n1133, A2 => n1134, A3 => n1135, A4 => n1136,
                           ZN => n1132);
   U974 : OAI221_X1 port map( B1 => n2154, B2 => n2930, C1 => n2150, C2 => 
                           n2866, A => n1141, ZN => n1140);
   U975 : AOI21_X1 port map( B1 => n1116, B2 => n1117, A => n1943, ZN => N310);
   U976 : NOR4_X1 port map( A1 => n1122, A2 => n1123, A3 => n1124, A4 => n1125,
                           ZN => n1116);
   U977 : NOR4_X1 port map( A1 => n1118, A2 => n1119, A3 => n1120, A4 => n1121,
                           ZN => n1117);
   U978 : OAI221_X1 port map( B1 => n2154, B2 => n2929, C1 => n2150, C2 => 
                           n2865, A => n1126, ZN => n1125);
   U979 : AOI21_X1 port map( B1 => n1101, B2 => n1102, A => n1943, ZN => N311);
   U980 : NOR4_X1 port map( A1 => n1107, A2 => n1108, A3 => n1109, A4 => n1110,
                           ZN => n1101);
   U981 : NOR4_X1 port map( A1 => n1103, A2 => n1104, A3 => n1105, A4 => n1106,
                           ZN => n1102);
   U982 : OAI221_X1 port map( B1 => n2154, B2 => n2928, C1 => n2150, C2 => 
                           n2864, A => n1111, ZN => n1110);
   U983 : AOI21_X1 port map( B1 => n1086, B2 => n1087, A => n1943, ZN => N312);
   U984 : NOR4_X1 port map( A1 => n1092, A2 => n1093, A3 => n1094, A4 => n1095,
                           ZN => n1086);
   U985 : NOR4_X1 port map( A1 => n1088, A2 => n1089, A3 => n1090, A4 => n1091,
                           ZN => n1087);
   U986 : OAI221_X1 port map( B1 => n2154, B2 => n2927, C1 => n2150, C2 => 
                           n2863, A => n1096, ZN => n1095);
   U987 : AOI21_X1 port map( B1 => n1071, B2 => n1072, A => n1943, ZN => N313);
   U988 : NOR4_X1 port map( A1 => n1077, A2 => n1078, A3 => n1079, A4 => n1080,
                           ZN => n1071);
   U989 : NOR4_X1 port map( A1 => n1073, A2 => n1074, A3 => n1075, A4 => n1076,
                           ZN => n1072);
   U990 : OAI221_X1 port map( B1 => n2154, B2 => n2926, C1 => n2150, C2 => 
                           n2862, A => n1081, ZN => n1080);
   U991 : AOI21_X1 port map( B1 => n1056, B2 => n1057, A => n1943, ZN => N314);
   U992 : NOR4_X1 port map( A1 => n1062, A2 => n1063, A3 => n1064, A4 => n1065,
                           ZN => n1056);
   U993 : NOR4_X1 port map( A1 => n1058, A2 => n1059, A3 => n1060, A4 => n1061,
                           ZN => n1057);
   U994 : OAI221_X1 port map( B1 => n2154, B2 => n2925, C1 => n2150, C2 => 
                           n2861, A => n1066, ZN => n1065);
   U995 : AOI21_X1 port map( B1 => n1041, B2 => n1042, A => n1944, ZN => N315);
   U996 : NOR4_X1 port map( A1 => n1047, A2 => n1048, A3 => n1049, A4 => n1050,
                           ZN => n1041);
   U997 : NOR4_X1 port map( A1 => n1043, A2 => n1044, A3 => n1045, A4 => n1046,
                           ZN => n1042);
   U998 : OAI221_X1 port map( B1 => n2155, B2 => n2924, C1 => n2151, C2 => 
                           n2860, A => n1051, ZN => n1050);
   U999 : AOI21_X1 port map( B1 => n1026, B2 => n1027, A => n1944, ZN => N316);
   U1000 : NOR4_X1 port map( A1 => n1032, A2 => n1033, A3 => n1034, A4 => n1035
                           , ZN => n1026);
   U1001 : NOR4_X1 port map( A1 => n1028, A2 => n1029, A3 => n1030, A4 => n1031
                           , ZN => n1027);
   U1002 : OAI221_X1 port map( B1 => n2155, B2 => n2923, C1 => n2151, C2 => 
                           n2859, A => n1036, ZN => n1035);
   U1003 : AOI21_X1 port map( B1 => n1011, B2 => n1012, A => n1944, ZN => N317)
                           ;
   U1004 : NOR4_X1 port map( A1 => n1017, A2 => n1018, A3 => n1019, A4 => n1020
                           , ZN => n1011);
   U1005 : NOR4_X1 port map( A1 => n1013, A2 => n1014, A3 => n1015, A4 => n1016
                           , ZN => n1012);
   U1006 : OAI221_X1 port map( B1 => n2155, B2 => n2922, C1 => n2151, C2 => 
                           n2858, A => n1021, ZN => n1020);
   U1007 : AOI21_X1 port map( B1 => n996, B2 => n997, A => n1944, ZN => N318);
   U1008 : NOR4_X1 port map( A1 => n1002, A2 => n1003, A3 => n1004, A4 => n1005
                           , ZN => n996);
   U1009 : NOR4_X1 port map( A1 => n998, A2 => n999, A3 => n1000, A4 => n1001, 
                           ZN => n997);
   U1010 : OAI221_X1 port map( B1 => n2155, B2 => n2921, C1 => n2151, C2 => 
                           n2857, A => n1006, ZN => n1005);
   U1011 : AOI21_X1 port map( B1 => n981, B2 => n982, A => n1944, ZN => N319);
   U1012 : NOR4_X1 port map( A1 => n987, A2 => n988, A3 => n989, A4 => n990, ZN
                           => n981);
   U1013 : NOR4_X1 port map( A1 => n983, A2 => n984, A3 => n985, A4 => n986, ZN
                           => n982);
   U1014 : OAI221_X1 port map( B1 => n2155, B2 => n2920, C1 => n2151, C2 => 
                           n2856, A => n991, ZN => n990);
   U1015 : AOI21_X1 port map( B1 => n966, B2 => n967, A => n1944, ZN => N320);
   U1016 : NOR4_X1 port map( A1 => n972, A2 => n973, A3 => n974, A4 => n975, ZN
                           => n966);
   U1017 : NOR4_X1 port map( A1 => n968, A2 => n969, A3 => n970, A4 => n971, ZN
                           => n967);
   U1018 : OAI221_X1 port map( B1 => n2155, B2 => n2919, C1 => n2151, C2 => 
                           n2855, A => n976, ZN => n975);
   U1019 : AOI21_X1 port map( B1 => n951, B2 => n952, A => n1944, ZN => N321);
   U1020 : NOR4_X1 port map( A1 => n957, A2 => n958, A3 => n959, A4 => n960, ZN
                           => n951);
   U1021 : NOR4_X1 port map( A1 => n953, A2 => n954, A3 => n955, A4 => n956, ZN
                           => n952);
   U1022 : OAI221_X1 port map( B1 => n2155, B2 => n2918, C1 => n2151, C2 => 
                           n2854, A => n961, ZN => n960);
   U1023 : AOI21_X1 port map( B1 => n904, B2 => n905, A => n1944, ZN => N322);
   U1024 : NOR4_X1 port map( A1 => n922, A2 => n923, A3 => n924, A4 => n925, ZN
                           => n904);
   U1025 : NOR4_X1 port map( A1 => n906, A2 => n907, A3 => n908, A4 => n909, ZN
                           => n905);
   U1026 : OAI221_X1 port map( B1 => n2155, B2 => n2917, C1 => n2151, C2 => 
                           n2853, A => n928, ZN => n925);
   U1027 : AOI21_X1 port map( B1 => n1916, B2 => n1917, A => n1945, ZN => N225)
                           ;
   U1028 : NOR4_X1 port map( A1 => n1924, A2 => n1925, A3 => n1926, A4 => n1927
                           , ZN => n1916);
   U1029 : NOR4_X1 port map( A1 => n1918, A2 => n1919, A3 => n1920, A4 => n1921
                           , ZN => n1917);
   U1030 : OAI221_X1 port map( B1 => n2948, B2 => n2025, C1 => n2884, C2 => 
                           n2021, A => n1928, ZN => n1927);
   U1031 : AOI21_X1 port map( B1 => n1901, B2 => n1902, A => n1945, ZN => N226)
                           ;
   U1032 : NOR4_X1 port map( A1 => n1907, A2 => n1908, A3 => n1909, A4 => n1910
                           , ZN => n1901);
   U1033 : NOR4_X1 port map( A1 => n1903, A2 => n1904, A3 => n1905, A4 => n1906
                           , ZN => n1902);
   U1034 : OAI221_X1 port map( B1 => n2947, B2 => n2025, C1 => n2883, C2 => 
                           n2021, A => n1911, ZN => n1910);
   U1035 : AOI21_X1 port map( B1 => n1886, B2 => n1887, A => n1945, ZN => N227)
                           ;
   U1036 : NOR4_X1 port map( A1 => n1892, A2 => n1893, A3 => n1894, A4 => n1895
                           , ZN => n1886);
   U1037 : NOR4_X1 port map( A1 => n1888, A2 => n1889, A3 => n1890, A4 => n1891
                           , ZN => n1887);
   U1038 : OAI221_X1 port map( B1 => n2946, B2 => n2025, C1 => n2882, C2 => 
                           n2021, A => n1896, ZN => n1895);
   U1039 : AOI21_X1 port map( B1 => n1871, B2 => n1872, A => n1945, ZN => N228)
                           ;
   U1040 : NOR4_X1 port map( A1 => n1877, A2 => n1878, A3 => n1879, A4 => n1880
                           , ZN => n1871);
   U1041 : NOR4_X1 port map( A1 => n1873, A2 => n1874, A3 => n1875, A4 => n1876
                           , ZN => n1872);
   U1042 : OAI221_X1 port map( B1 => n2945, B2 => n2025, C1 => n2881, C2 => 
                           n2021, A => n1881, ZN => n1880);
   U1043 : AOI21_X1 port map( B1 => n1856, B2 => n1857, A => n1945, ZN => N229)
                           ;
   U1044 : NOR4_X1 port map( A1 => n1862, A2 => n1863, A3 => n1864, A4 => n1865
                           , ZN => n1856);
   U1045 : NOR4_X1 port map( A1 => n1858, A2 => n1859, A3 => n1860, A4 => n1861
                           , ZN => n1857);
   U1046 : OAI221_X1 port map( B1 => n2944, B2 => n2025, C1 => n2880, C2 => 
                           n2021, A => n1866, ZN => n1865);
   U1047 : AOI21_X1 port map( B1 => n1841, B2 => n1842, A => n1945, ZN => N230)
                           ;
   U1048 : NOR4_X1 port map( A1 => n1847, A2 => n1848, A3 => n1849, A4 => n1850
                           , ZN => n1841);
   U1049 : NOR4_X1 port map( A1 => n1843, A2 => n1844, A3 => n1845, A4 => n1846
                           , ZN => n1842);
   U1050 : OAI221_X1 port map( B1 => n2943, B2 => n2025, C1 => n2879, C2 => 
                           n2021, A => n1851, ZN => n1850);
   U1051 : AOI21_X1 port map( B1 => n1826, B2 => n1827, A => n1945, ZN => N231)
                           ;
   U1052 : NOR4_X1 port map( A1 => n1832, A2 => n1833, A3 => n1834, A4 => n1835
                           , ZN => n1826);
   U1053 : NOR4_X1 port map( A1 => n1828, A2 => n1829, A3 => n1830, A4 => n1831
                           , ZN => n1827);
   U1054 : OAI221_X1 port map( B1 => n2942, B2 => n2025, C1 => n2878, C2 => 
                           n2021, A => n1836, ZN => n1835);
   U1055 : AOI21_X1 port map( B1 => n1811, B2 => n1812, A => n1945, ZN => N232)
                           ;
   U1056 : NOR4_X1 port map( A1 => n1817, A2 => n1818, A3 => n1819, A4 => n1820
                           , ZN => n1811);
   U1057 : NOR4_X1 port map( A1 => n1813, A2 => n1814, A3 => n1815, A4 => n1816
                           , ZN => n1812);
   U1058 : OAI221_X1 port map( B1 => n2941, B2 => n2025, C1 => n2877, C2 => 
                           n2021, A => n1821, ZN => n1820);
   U1059 : AOI21_X1 port map( B1 => n1796, B2 => n1797, A => n1945, ZN => N233)
                           ;
   U1060 : NOR4_X1 port map( A1 => n1802, A2 => n1803, A3 => n1804, A4 => n1805
                           , ZN => n1796);
   U1061 : NOR4_X1 port map( A1 => n1798, A2 => n1799, A3 => n1800, A4 => n1801
                           , ZN => n1797);
   U1062 : OAI221_X1 port map( B1 => n2940, B2 => n2025, C1 => n2876, C2 => 
                           n2021, A => n1806, ZN => n1805);
   U1063 : AOI21_X1 port map( B1 => n1781, B2 => n1782, A => n1945, ZN => N234)
                           ;
   U1064 : NOR4_X1 port map( A1 => n1787, A2 => n1788, A3 => n1789, A4 => n1790
                           , ZN => n1781);
   U1065 : NOR4_X1 port map( A1 => n1783, A2 => n1784, A3 => n1785, A4 => n1786
                           , ZN => n1782);
   U1066 : OAI221_X1 port map( B1 => n2939, B2 => n2025, C1 => n2875, C2 => 
                           n2021, A => n1791, ZN => n1790);
   U1067 : AOI21_X1 port map( B1 => n1766, B2 => n1767, A => n1945, ZN => N235)
                           ;
   U1068 : NOR4_X1 port map( A1 => n1772, A2 => n1773, A3 => n1774, A4 => n1775
                           , ZN => n1766);
   U1069 : NOR4_X1 port map( A1 => n1768, A2 => n1769, A3 => n1770, A4 => n1771
                           , ZN => n1767);
   U1070 : OAI221_X1 port map( B1 => n2938, B2 => n2025, C1 => n2874, C2 => 
                           n2021, A => n1776, ZN => n1775);
   U1071 : AOI21_X1 port map( B1 => n1751, B2 => n1752, A => n1945, ZN => N236)
                           ;
   U1072 : NOR4_X1 port map( A1 => n1757, A2 => n1758, A3 => n1759, A4 => n1760
                           , ZN => n1751);
   U1073 : NOR4_X1 port map( A1 => n1753, A2 => n1754, A3 => n1755, A4 => n1756
                           , ZN => n1752);
   U1074 : OAI221_X1 port map( B1 => n2937, B2 => n2025, C1 => n2873, C2 => 
                           n2021, A => n1761, ZN => n1760);
   U1075 : AOI21_X1 port map( B1 => n1736, B2 => n1737, A => n1946, ZN => N237)
                           ;
   U1076 : NOR4_X1 port map( A1 => n1742, A2 => n1743, A3 => n1744, A4 => n1745
                           , ZN => n1736);
   U1077 : NOR4_X1 port map( A1 => n1738, A2 => n1739, A3 => n1740, A4 => n1741
                           , ZN => n1737);
   U1078 : OAI221_X1 port map( B1 => n2936, B2 => n2026, C1 => n2872, C2 => 
                           n2022, A => n1746, ZN => n1745);
   U1079 : AOI21_X1 port map( B1 => n1721, B2 => n1722, A => n1946, ZN => N238)
                           ;
   U1080 : NOR4_X1 port map( A1 => n1727, A2 => n1728, A3 => n1729, A4 => n1730
                           , ZN => n1721);
   U1081 : NOR4_X1 port map( A1 => n1723, A2 => n1724, A3 => n1725, A4 => n1726
                           , ZN => n1722);
   U1082 : OAI221_X1 port map( B1 => n2935, B2 => n2026, C1 => n2871, C2 => 
                           n2022, A => n1731, ZN => n1730);
   U1083 : AOI21_X1 port map( B1 => n1706, B2 => n1707, A => n1946, ZN => N239)
                           ;
   U1084 : NOR4_X1 port map( A1 => n1712, A2 => n1713, A3 => n1714, A4 => n1715
                           , ZN => n1706);
   U1085 : NOR4_X1 port map( A1 => n1708, A2 => n1709, A3 => n1710, A4 => n1711
                           , ZN => n1707);
   U1086 : OAI221_X1 port map( B1 => n2934, B2 => n2026, C1 => n2870, C2 => 
                           n2022, A => n1716, ZN => n1715);
   U1087 : AOI21_X1 port map( B1 => n1691, B2 => n1692, A => n1946, ZN => N240)
                           ;
   U1088 : NOR4_X1 port map( A1 => n1697, A2 => n1698, A3 => n1699, A4 => n1700
                           , ZN => n1691);
   U1089 : NOR4_X1 port map( A1 => n1693, A2 => n1694, A3 => n1695, A4 => n1696
                           , ZN => n1692);
   U1090 : OAI221_X1 port map( B1 => n2933, B2 => n2026, C1 => n2869, C2 => 
                           n2022, A => n1701, ZN => n1700);
   U1091 : AOI21_X1 port map( B1 => n1676, B2 => n1677, A => n1946, ZN => N241)
                           ;
   U1092 : NOR4_X1 port map( A1 => n1682, A2 => n1683, A3 => n1684, A4 => n1685
                           , ZN => n1676);
   U1093 : NOR4_X1 port map( A1 => n1678, A2 => n1679, A3 => n1680, A4 => n1681
                           , ZN => n1677);
   U1094 : OAI221_X1 port map( B1 => n2932, B2 => n2026, C1 => n2868, C2 => 
                           n2022, A => n1686, ZN => n1685);
   U1095 : AOI21_X1 port map( B1 => n1661, B2 => n1662, A => n1946, ZN => N242)
                           ;
   U1096 : NOR4_X1 port map( A1 => n1667, A2 => n1668, A3 => n1669, A4 => n1670
                           , ZN => n1661);
   U1097 : NOR4_X1 port map( A1 => n1663, A2 => n1664, A3 => n1665, A4 => n1666
                           , ZN => n1662);
   U1098 : OAI221_X1 port map( B1 => n2931, B2 => n2026, C1 => n2867, C2 => 
                           n2022, A => n1671, ZN => n1670);
   U1099 : AOI21_X1 port map( B1 => n1646, B2 => n1647, A => n1946, ZN => N243)
                           ;
   U1100 : NOR4_X1 port map( A1 => n1652, A2 => n1653, A3 => n1654, A4 => n1655
                           , ZN => n1646);
   U1101 : NOR4_X1 port map( A1 => n1648, A2 => n1649, A3 => n1650, A4 => n1651
                           , ZN => n1647);
   U1102 : OAI221_X1 port map( B1 => n2930, B2 => n2026, C1 => n2866, C2 => 
                           n2022, A => n1656, ZN => n1655);
   U1103 : AOI21_X1 port map( B1 => n1631, B2 => n1632, A => n1946, ZN => N244)
                           ;
   U1104 : NOR4_X1 port map( A1 => n1637, A2 => n1638, A3 => n1639, A4 => n1640
                           , ZN => n1631);
   U1105 : NOR4_X1 port map( A1 => n1633, A2 => n1634, A3 => n1635, A4 => n1636
                           , ZN => n1632);
   U1106 : OAI221_X1 port map( B1 => n2929, B2 => n2026, C1 => n2865, C2 => 
                           n2022, A => n1641, ZN => n1640);
   U1107 : AOI21_X1 port map( B1 => n1616, B2 => n1617, A => n1946, ZN => N245)
                           ;
   U1108 : NOR4_X1 port map( A1 => n1622, A2 => n1623, A3 => n1624, A4 => n1625
                           , ZN => n1616);
   U1109 : NOR4_X1 port map( A1 => n1618, A2 => n1619, A3 => n1620, A4 => n1621
                           , ZN => n1617);
   U1110 : OAI221_X1 port map( B1 => n2928, B2 => n2026, C1 => n2864, C2 => 
                           n2022, A => n1626, ZN => n1625);
   U1111 : AOI21_X1 port map( B1 => n1601, B2 => n1602, A => n1946, ZN => N246)
                           ;
   U1112 : NOR4_X1 port map( A1 => n1607, A2 => n1608, A3 => n1609, A4 => n1610
                           , ZN => n1601);
   U1113 : NOR4_X1 port map( A1 => n1603, A2 => n1604, A3 => n1605, A4 => n1606
                           , ZN => n1602);
   U1114 : OAI221_X1 port map( B1 => n2927, B2 => n2026, C1 => n2863, C2 => 
                           n2022, A => n1611, ZN => n1610);
   U1115 : AOI21_X1 port map( B1 => n1586, B2 => n1587, A => n1946, ZN => N247)
                           ;
   U1116 : NOR4_X1 port map( A1 => n1592, A2 => n1593, A3 => n1594, A4 => n1595
                           , ZN => n1586);
   U1117 : NOR4_X1 port map( A1 => n1588, A2 => n1589, A3 => n1590, A4 => n1591
                           , ZN => n1587);
   U1118 : OAI221_X1 port map( B1 => n2926, B2 => n2026, C1 => n2862, C2 => 
                           n2022, A => n1596, ZN => n1595);
   U1119 : AOI21_X1 port map( B1 => n1571, B2 => n1572, A => n1946, ZN => N248)
                           ;
   U1120 : NOR4_X1 port map( A1 => n1577, A2 => n1578, A3 => n1579, A4 => n1580
                           , ZN => n1571);
   U1121 : NOR4_X1 port map( A1 => n1573, A2 => n1574, A3 => n1575, A4 => n1576
                           , ZN => n1572);
   U1122 : OAI221_X1 port map( B1 => n2925, B2 => n2026, C1 => n2861, C2 => 
                           n2022, A => n1581, ZN => n1580);
   U1123 : AOI21_X1 port map( B1 => n1556, B2 => n1557, A => n1947, ZN => N249)
                           ;
   U1124 : NOR4_X1 port map( A1 => n1562, A2 => n1563, A3 => n1564, A4 => n1565
                           , ZN => n1556);
   U1125 : NOR4_X1 port map( A1 => n1558, A2 => n1559, A3 => n1560, A4 => n1561
                           , ZN => n1557);
   U1126 : OAI221_X1 port map( B1 => n2924, B2 => n2027, C1 => n2860, C2 => 
                           n2023, A => n1566, ZN => n1565);
   U1127 : AOI21_X1 port map( B1 => n1541, B2 => n1542, A => n1947, ZN => N250)
                           ;
   U1128 : NOR4_X1 port map( A1 => n1547, A2 => n1548, A3 => n1549, A4 => n1550
                           , ZN => n1541);
   U1129 : NOR4_X1 port map( A1 => n1543, A2 => n1544, A3 => n1545, A4 => n1546
                           , ZN => n1542);
   U1130 : OAI221_X1 port map( B1 => n2923, B2 => n2027, C1 => n2859, C2 => 
                           n2023, A => n1551, ZN => n1550);
   U1131 : AOI21_X1 port map( B1 => n1526, B2 => n1527, A => n1947, ZN => N251)
                           ;
   U1132 : NOR4_X1 port map( A1 => n1532, A2 => n1533, A3 => n1534, A4 => n1535
                           , ZN => n1526);
   U1133 : NOR4_X1 port map( A1 => n1528, A2 => n1529, A3 => n1530, A4 => n1531
                           , ZN => n1527);
   U1134 : OAI221_X1 port map( B1 => n2922, B2 => n2027, C1 => n2858, C2 => 
                           n2023, A => n1536, ZN => n1535);
   U1135 : AOI21_X1 port map( B1 => n1511, B2 => n1512, A => n1947, ZN => N252)
                           ;
   U1136 : NOR4_X1 port map( A1 => n1517, A2 => n1518, A3 => n1519, A4 => n1520
                           , ZN => n1511);
   U1137 : NOR4_X1 port map( A1 => n1513, A2 => n1514, A3 => n1515, A4 => n1516
                           , ZN => n1512);
   U1138 : OAI221_X1 port map( B1 => n2921, B2 => n2027, C1 => n2857, C2 => 
                           n2023, A => n1521, ZN => n1520);
   U1139 : AOI21_X1 port map( B1 => n1496, B2 => n1497, A => n1947, ZN => N253)
                           ;
   U1140 : NOR4_X1 port map( A1 => n1502, A2 => n1503, A3 => n1504, A4 => n1505
                           , ZN => n1496);
   U1141 : NOR4_X1 port map( A1 => n1498, A2 => n1499, A3 => n1500, A4 => n1501
                           , ZN => n1497);
   U1142 : OAI221_X1 port map( B1 => n2920, B2 => n2027, C1 => n2856, C2 => 
                           n2023, A => n1506, ZN => n1505);
   U1143 : AOI21_X1 port map( B1 => n1481, B2 => n1482, A => n1947, ZN => N254)
                           ;
   U1144 : NOR4_X1 port map( A1 => n1487, A2 => n1488, A3 => n1489, A4 => n1490
                           , ZN => n1481);
   U1145 : NOR4_X1 port map( A1 => n1483, A2 => n1484, A3 => n1485, A4 => n1486
                           , ZN => n1482);
   U1146 : OAI221_X1 port map( B1 => n2919, B2 => n2027, C1 => n2855, C2 => 
                           n2023, A => n1491, ZN => n1490);
   U1147 : AOI21_X1 port map( B1 => n1466, B2 => n1467, A => n1947, ZN => N255)
                           ;
   U1148 : NOR4_X1 port map( A1 => n1472, A2 => n1473, A3 => n1474, A4 => n1475
                           , ZN => n1466);
   U1149 : NOR4_X1 port map( A1 => n1468, A2 => n1469, A3 => n1470, A4 => n1471
                           , ZN => n1467);
   U1150 : OAI221_X1 port map( B1 => n2918, B2 => n2027, C1 => n2854, C2 => 
                           n2023, A => n1476, ZN => n1475);
   U1151 : AOI21_X1 port map( B1 => n1419, B2 => n1420, A => n1947, ZN => N256)
                           ;
   U1152 : NOR4_X1 port map( A1 => n1437, A2 => n1438, A3 => n1439, A4 => n1440
                           , ZN => n1419);
   U1153 : NOR4_X1 port map( A1 => n1421, A2 => n1422, A3 => n1423, A4 => n1424
                           , ZN => n1420);
   U1154 : OAI221_X1 port map( B1 => n2917, B2 => n2027, C1 => n2853, C2 => 
                           n2023, A => n1443, ZN => n1440);
   U1155 : NAND2_X1 port map( A1 => n2143, A2 => n1407, ZN => n912);
   U1156 : NAND2_X1 port map( A1 => n2130, A2 => n1407, ZN => n911);
   U1157 : NAND2_X1 port map( A1 => n2134, A2 => n1407, ZN => n913);
   U1158 : NAND2_X1 port map( A1 => n2123, A2 => n1407, ZN => n918);
   U1159 : NAND2_X1 port map( A1 => n2127, A2 => n1407, ZN => n917);
   U1160 : NAND2_X1 port map( A1 => n2118, A2 => n1407, ZN => n920);
   U1161 : NAND2_X1 port map( A1 => n2139, A2 => n1407, ZN => n948);
   U1162 : NAND2_X1 port map( A1 => n2015, A2 => n1922, ZN => n1427);
   U1163 : NAND2_X1 port map( A1 => n2000, A2 => n1922, ZN => n1426);
   U1164 : NAND2_X1 port map( A1 => n2006, A2 => n1922, ZN => n1428);
   U1165 : NAND2_X1 port map( A1 => n1995, A2 => n1922, ZN => n1433);
   U1166 : NAND2_X1 port map( A1 => n1999, A2 => n1922, ZN => n1432);
   U1167 : NAND2_X1 port map( A1 => n1990, A2 => n1922, ZN => n1435);
   U1168 : NAND2_X1 port map( A1 => n2011, A2 => n1922, ZN => n1463);
   U1169 : NAND2_X1 port map( A1 => n1418, A2 => n2128, ZN => n944);
   U1170 : NAND2_X1 port map( A1 => n1418, A2 => n2123, ZN => n943);
   U1171 : NAND2_X1 port map( A1 => n1418, A2 => n2134, ZN => n942);
   U1172 : NAND2_X1 port map( A1 => n1418, A2 => n2127, ZN => n947);
   U1173 : NAND2_X1 port map( A1 => n1418, A2 => n2118, ZN => n946);
   U1174 : NAND2_X1 port map( A1 => n1418, A2 => n2112, ZN => n945);
   U1175 : NAND2_X1 port map( A1 => n1418, A2 => n2143, ZN => n926);
   U1176 : NAND2_X1 port map( A1 => n1418, A2 => n2139, ZN => n927);
   U1177 : NAND2_X1 port map( A1 => n1933, A2 => n2000, ZN => n1459);
   U1178 : NAND2_X1 port map( A1 => n1933, A2 => n1995, ZN => n1458);
   U1179 : NAND2_X1 port map( A1 => n1933, A2 => n2004, ZN => n1457);
   U1180 : NAND2_X1 port map( A1 => n1933, A2 => n1999, ZN => n1462);
   U1181 : NAND2_X1 port map( A1 => n1933, A2 => n1988, ZN => n1461);
   U1182 : NAND2_X1 port map( A1 => n1933, A2 => n1984, ZN => n1460);
   U1183 : NAND2_X1 port map( A1 => n1933, A2 => n2011, ZN => n1442);
   U1184 : NAND2_X1 port map( A1 => n1933, A2 => n2015, ZN => n1441);
   U1185 : NAND2_X1 port map( A1 => n2336, A2 => n3220, ZN => n892);
   U1186 : INV_X1 port map( A => RD2, ZN => n3205);
   U1187 : INV_X1 port map( A => RD1, ZN => n3206);
   U1188 : BUF_X1 port map( A => n1991, Z => n1988);
   U1189 : BUF_X1 port map( A => n1991, Z => n1989);
   U1190 : BUF_X1 port map( A => n2119, Z => n2116);
   U1191 : BUF_X1 port map( A => n2119, Z => n2117);
   U1192 : BUF_X1 port map( A => n2007, Z => n2004);
   U1193 : BUF_X1 port map( A => n2131, Z => n2128);
   U1194 : BUF_X1 port map( A => n2115, Z => n2112);
   U1195 : BUF_X1 port map( A => n2131, Z => n2129);
   U1196 : BUF_X1 port map( A => n2115, Z => n2113);
   U1197 : BUF_X1 port map( A => n2007, Z => n2005);
   U1198 : BUF_X1 port map( A => n2003, Z => n2000);
   U1199 : BUF_X1 port map( A => n1987, Z => n1984);
   U1200 : BUF_X1 port map( A => n2003, Z => n2001);
   U1201 : BUF_X1 port map( A => n1987, Z => n1985);
   U1202 : BUF_X1 port map( A => n2147, Z => n2144);
   U1203 : BUF_X1 port map( A => n2147, Z => n2145);
   U1204 : BUF_X1 port map( A => n2019, Z => n2016);
   U1205 : BUF_X1 port map( A => n2019, Z => n2017);
   U1206 : BUF_X1 port map( A => n2119, Z => n2118);
   U1207 : BUF_X1 port map( A => n2131, Z => n2130);
   U1208 : BUF_X1 port map( A => n2115, Z => n2114);
   U1209 : BUF_X1 port map( A => n1991, Z => n1990);
   U1210 : BUF_X1 port map( A => n2007, Z => n2006);
   U1211 : BUF_X1 port map( A => n2003, Z => n2002);
   U1212 : BUF_X1 port map( A => n2147, Z => n2146);
   U1213 : BUF_X1 port map( A => n2019, Z => n2018);
   U1214 : BUF_X1 port map( A => n1987, Z => n1986);
   U1215 : BUF_X1 port map( A => n1939, Z => n2127);
   U1216 : BUF_X1 port map( A => n1940, Z => n2143);
   U1217 : BUF_X1 port map( A => n1941, Z => n2139);
   U1218 : BUF_X1 port map( A => n1937, Z => n1995);
   U1219 : BUF_X1 port map( A => n1938, Z => n1999);
   U1220 : BUF_X1 port map( A => n1935, Z => n2011);
   U1221 : BUF_X1 port map( A => n1936, Z => n2015);
   U1222 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n2134, B1 => 
                           REGISTERS_9_0_port, B2 => n2128, ZN => n1416);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n2134, B1 => 
                           REGISTERS_9_1_port, B2 => n2130, ZN => n1399);
   U1224 : AOI22_X1 port map( A1 => REGISTERS_11_2_port, A2 => n2134, B1 => 
                           REGISTERS_9_2_port, B2 => n2130, ZN => n1384);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n2134, B1 => 
                           REGISTERS_9_3_port, B2 => n2130, ZN => n1369);
   U1226 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n2134, B1 => 
                           REGISTERS_9_4_port, B2 => n2130, ZN => n1354);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n2134, B1 => 
                           REGISTERS_9_5_port, B2 => n2130, ZN => n1339);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n2134, B1 => 
                           REGISTERS_9_6_port, B2 => n2130, ZN => n1324);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n2134, B1 => 
                           REGISTERS_9_7_port, B2 => n2130, ZN => n1309);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n2133, B1 => 
                           REGISTERS_9_8_port, B2 => n2130, ZN => n1294);
   U1231 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n2133, B1 => 
                           REGISTERS_9_9_port, B2 => n2130, ZN => n1279);
   U1232 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n2133, B1 => 
                           REGISTERS_9_10_port, B2 => n2129, ZN => n1264);
   U1233 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n2133, B1 => 
                           REGISTERS_9_11_port, B2 => n2129, ZN => n1249);
   U1234 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n2133, B1 => 
                           REGISTERS_9_12_port, B2 => n2129, ZN => n1234);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_11_13_port, A2 => n2133, B1 => 
                           REGISTERS_9_13_port, B2 => n2129, ZN => n1219);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n2133, B1 => 
                           REGISTERS_9_14_port, B2 => n2129, ZN => n1204);
   U1237 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n2133, B1 => 
                           REGISTERS_9_15_port, B2 => n2129, ZN => n1189);
   U1238 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n2133, B1 => 
                           REGISTERS_9_16_port, B2 => n2129, ZN => n1174);
   U1239 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n2133, B1 => 
                           REGISTERS_9_17_port, B2 => n2129, ZN => n1159);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_11_18_port, A2 => n2133, B1 => 
                           REGISTERS_9_18_port, B2 => n2129, ZN => n1144);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n2132, B1 => 
                           REGISTERS_9_19_port, B2 => n2129, ZN => n1129);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n2132, B1 => 
                           REGISTERS_9_20_port, B2 => n2129, ZN => n1114);
   U1243 : AOI22_X1 port map( A1 => REGISTERS_11_21_port, A2 => n2132, B1 => 
                           REGISTERS_9_21_port, B2 => n2128, ZN => n1099);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n2132, B1 => 
                           REGISTERS_9_22_port, B2 => n2128, ZN => n1084);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n2132, B1 => 
                           REGISTERS_9_23_port, B2 => n2128, ZN => n1069);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n2132, B1 => 
                           REGISTERS_9_24_port, B2 => n2128, ZN => n1054);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n2132, B1 => 
                           REGISTERS_9_25_port, B2 => n2128, ZN => n1039);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n2132, B1 => 
                           REGISTERS_9_26_port, B2 => n2128, ZN => n1024);
   U1249 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n2132, B1 => 
                           REGISTERS_9_27_port, B2 => n2128, ZN => n1009);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n2132, B1 => 
                           REGISTERS_9_28_port, B2 => n2128, ZN => n994);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n2132, B1 => 
                           REGISTERS_9_29_port, B2 => n2128, ZN => n979);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_11_30_port, A2 => n2132, B1 => 
                           REGISTERS_9_30_port, B2 => n2128, ZN => n964);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n2133, B1 => 
                           REGISTERS_9_31_port, B2 => n2129, ZN => n934);
   U1254 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_0_port, B1 => 
                           n2000, B2 => REGISTERS_9_0_port, ZN => n1931);
   U1255 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_1_port, B1 => 
                           n2002, B2 => REGISTERS_9_1_port, ZN => n1914);
   U1256 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_2_port, B1 => 
                           n2002, B2 => REGISTERS_9_2_port, ZN => n1899);
   U1257 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_3_port, B1 => 
                           n2002, B2 => REGISTERS_9_3_port, ZN => n1884);
   U1258 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_4_port, B1 => 
                           n2002, B2 => REGISTERS_9_4_port, ZN => n1869);
   U1259 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_5_port, B1 => 
                           n2002, B2 => REGISTERS_9_5_port, ZN => n1854);
   U1260 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_6_port, B1 => 
                           n2002, B2 => REGISTERS_9_6_port, ZN => n1839);
   U1261 : AOI22_X1 port map( A1 => n2006, A2 => REGISTERS_11_7_port, B1 => 
                           n2002, B2 => REGISTERS_9_7_port, ZN => n1824);
   U1262 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_8_port, B1 => 
                           n2002, B2 => REGISTERS_9_8_port, ZN => n1809);
   U1263 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_9_port, B1 => 
                           n2002, B2 => REGISTERS_9_9_port, ZN => n1794);
   U1264 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_10_port, B1 => 
                           n2001, B2 => REGISTERS_9_10_port, ZN => n1779);
   U1265 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_11_port, B1 => 
                           n2001, B2 => REGISTERS_9_11_port, ZN => n1764);
   U1266 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_12_port, B1 => 
                           n2001, B2 => REGISTERS_9_12_port, ZN => n1749);
   U1267 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_13_port, B1 => 
                           n2001, B2 => REGISTERS_9_13_port, ZN => n1734);
   U1268 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_14_port, B1 => 
                           n2001, B2 => REGISTERS_9_14_port, ZN => n1719);
   U1269 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_15_port, B1 => 
                           n2001, B2 => REGISTERS_9_15_port, ZN => n1704);
   U1270 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_16_port, B1 => 
                           n2001, B2 => REGISTERS_9_16_port, ZN => n1689);
   U1271 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_17_port, B1 => 
                           n2001, B2 => REGISTERS_9_17_port, ZN => n1674);
   U1272 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_18_port, B1 => 
                           n2001, B2 => REGISTERS_9_18_port, ZN => n1659);
   U1273 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_19_port, B1 => 
                           n2001, B2 => REGISTERS_9_19_port, ZN => n1644);
   U1274 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_20_port, B1 => 
                           n2001, B2 => REGISTERS_9_20_port, ZN => n1629);
   U1275 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_21_port, B1 => 
                           n2001, B2 => REGISTERS_9_21_port, ZN => n1614);
   U1276 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_22_port, B1 => 
                           n2000, B2 => REGISTERS_9_22_port, ZN => n1599);
   U1277 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_23_port, B1 => 
                           n2000, B2 => REGISTERS_9_23_port, ZN => n1584);
   U1278 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_24_port, B1 => 
                           n2000, B2 => REGISTERS_9_24_port, ZN => n1569);
   U1279 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_25_port, B1 => 
                           n2000, B2 => REGISTERS_9_25_port, ZN => n1554);
   U1280 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_26_port, B1 => 
                           n2000, B2 => REGISTERS_9_26_port, ZN => n1539);
   U1281 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_27_port, B1 => 
                           n2000, B2 => REGISTERS_9_27_port, ZN => n1524);
   U1282 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_28_port, B1 => 
                           n2000, B2 => REGISTERS_9_28_port, ZN => n1509);
   U1283 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_29_port, B1 => 
                           n2000, B2 => REGISTERS_9_29_port, ZN => n1494);
   U1284 : AOI22_X1 port map( A1 => n2004, A2 => REGISTERS_11_30_port, B1 => 
                           n2000, B2 => REGISTERS_9_30_port, ZN => n1479);
   U1285 : AOI22_X1 port map( A1 => n2005, A2 => REGISTERS_11_31_port, B1 => 
                           n2001, B2 => REGISTERS_9_31_port, ZN => n1449);
   U1286 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => n3214, A3 => ADD_RD1(0), 
                           ZN => n1935);
   U1287 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), A3 => 
                           ADD_RD1(0), ZN => n1936);
   U1288 : AND3_X1 port map( A1 => n3215, A2 => n3214, A3 => ADD_RD1(2), ZN => 
                           n1937);
   U1289 : AND3_X1 port map( A1 => ADD_RD1(1), A2 => n3215, A3 => ADD_RD1(2), 
                           ZN => n1938);
   U1290 : AND3_X1 port map( A1 => ADD_RD2(1), A2 => n3219, A3 => ADD_RD2(2), 
                           ZN => n1939);
   U1291 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => 
                           ADD_RD2(0), ZN => n1940);
   U1292 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => n3218, A3 => ADD_RD2(0), 
                           ZN => n1941);
   U1293 : OAI21_X1 port map( B1 => n1414, B2 => n1415, A => n2144, ZN => n1413
                           );
   U1294 : OAI221_X1 port map( B1 => n2124, B2 => n2660, C1 => n2120, C2 => 
                           n2596, A => n1417, ZN => n1414);
   U1295 : OAI221_X1 port map( B1 => n2140, B2 => n2692, C1 => n2136, C2 => 
                           n2628, A => n1416, ZN => n1415);
   U1296 : AOI22_X1 port map( A1 => REGISTERS_10_0_port, A2 => n2118, B1 => 
                           REGISTERS_8_0_port, B2 => n2112, ZN => n1417);
   U1297 : OAI21_X1 port map( B1 => n1397, B2 => n1398, A => n2144, ZN => n1396
                           );
   U1298 : OAI221_X1 port map( B1 => n2124, B2 => n2659, C1 => n2120, C2 => 
                           n2595, A => n1400, ZN => n1397);
   U1299 : OAI221_X1 port map( B1 => n2140, B2 => n2691, C1 => n2136, C2 => 
                           n2627, A => n1399, ZN => n1398);
   U1300 : AOI22_X1 port map( A1 => REGISTERS_10_1_port, A2 => n2118, B1 => 
                           REGISTERS_8_1_port, B2 => n2114, ZN => n1400);
   U1301 : OAI21_X1 port map( B1 => n1382, B2 => n1383, A => n2144, ZN => n1381
                           );
   U1302 : OAI221_X1 port map( B1 => n2124, B2 => n2658, C1 => n2120, C2 => 
                           n2594, A => n1385, ZN => n1382);
   U1303 : OAI221_X1 port map( B1 => n2140, B2 => n2690, C1 => n2136, C2 => 
                           n2626, A => n1384, ZN => n1383);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n2118, B1 => 
                           REGISTERS_8_2_port, B2 => n2114, ZN => n1385);
   U1305 : OAI21_X1 port map( B1 => n1367, B2 => n1368, A => n2144, ZN => n1366
                           );
   U1306 : OAI221_X1 port map( B1 => n2124, B2 => n2657, C1 => n2120, C2 => 
                           n2593, A => n1370, ZN => n1367);
   U1307 : OAI221_X1 port map( B1 => n2140, B2 => n2689, C1 => n2136, C2 => 
                           n2625, A => n1369, ZN => n1368);
   U1308 : AOI22_X1 port map( A1 => REGISTERS_10_3_port, A2 => n2118, B1 => 
                           REGISTERS_8_3_port, B2 => n2114, ZN => n1370);
   U1309 : OAI21_X1 port map( B1 => n1352, B2 => n1353, A => n2144, ZN => n1351
                           );
   U1310 : OAI221_X1 port map( B1 => n2124, B2 => n2656, C1 => n2120, C2 => 
                           n2592, A => n1355, ZN => n1352);
   U1311 : OAI221_X1 port map( B1 => n2140, B2 => n2688, C1 => n2136, C2 => 
                           n2624, A => n1354, ZN => n1353);
   U1312 : AOI22_X1 port map( A1 => REGISTERS_10_4_port, A2 => n2118, B1 => 
                           REGISTERS_8_4_port, B2 => n2114, ZN => n1355);
   U1313 : OAI21_X1 port map( B1 => n1337, B2 => n1338, A => n2144, ZN => n1336
                           );
   U1314 : OAI221_X1 port map( B1 => n2124, B2 => n2655, C1 => n2120, C2 => 
                           n2591, A => n1340, ZN => n1337);
   U1315 : OAI221_X1 port map( B1 => n2140, B2 => n2687, C1 => n2136, C2 => 
                           n2623, A => n1339, ZN => n1338);
   U1316 : AOI22_X1 port map( A1 => REGISTERS_10_5_port, A2 => n2118, B1 => 
                           REGISTERS_8_5_port, B2 => n2114, ZN => n1340);
   U1317 : OAI21_X1 port map( B1 => n1322, B2 => n1323, A => n2144, ZN => n1321
                           );
   U1318 : OAI221_X1 port map( B1 => n2124, B2 => n2654, C1 => n2120, C2 => 
                           n2590, A => n1325, ZN => n1322);
   U1319 : OAI221_X1 port map( B1 => n2140, B2 => n2686, C1 => n2136, C2 => 
                           n2622, A => n1324, ZN => n1323);
   U1320 : AOI22_X1 port map( A1 => REGISTERS_10_6_port, A2 => n2118, B1 => 
                           REGISTERS_8_6_port, B2 => n2114, ZN => n1325);
   U1321 : OAI21_X1 port map( B1 => n1307, B2 => n1308, A => n2144, ZN => n1306
                           );
   U1322 : OAI221_X1 port map( B1 => n2124, B2 => n2653, C1 => n2120, C2 => 
                           n2589, A => n1310, ZN => n1307);
   U1323 : OAI221_X1 port map( B1 => n2140, B2 => n2685, C1 => n2136, C2 => 
                           n2621, A => n1309, ZN => n1308);
   U1324 : AOI22_X1 port map( A1 => REGISTERS_10_7_port, A2 => n2118, B1 => 
                           REGISTERS_8_7_port, B2 => n2114, ZN => n1310);
   U1325 : OAI21_X1 port map( B1 => n1292, B2 => n1293, A => n2144, ZN => n1291
                           );
   U1326 : OAI221_X1 port map( B1 => n2124, B2 => n2652, C1 => n2120, C2 => 
                           n2588, A => n1295, ZN => n1292);
   U1327 : OAI221_X1 port map( B1 => n2140, B2 => n2684, C1 => n2136, C2 => 
                           n2620, A => n1294, ZN => n1293);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_10_8_port, A2 => n2117, B1 => 
                           REGISTERS_8_8_port, B2 => n2114, ZN => n1295);
   U1329 : OAI21_X1 port map( B1 => n1277, B2 => n1278, A => n2144, ZN => n1276
                           );
   U1330 : OAI221_X1 port map( B1 => n2124, B2 => n2651, C1 => n2120, C2 => 
                           n2587, A => n1280, ZN => n1277);
   U1331 : OAI221_X1 port map( B1 => n2140, B2 => n2683, C1 => n2136, C2 => 
                           n2619, A => n1279, ZN => n1278);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_10_9_port, A2 => n2117, B1 => 
                           REGISTERS_8_9_port, B2 => n2114, ZN => n1280);
   U1333 : OAI21_X1 port map( B1 => n1262, B2 => n1263, A => n2144, ZN => n1261
                           );
   U1334 : OAI221_X1 port map( B1 => n2124, B2 => n2650, C1 => n2120, C2 => 
                           n2586, A => n1265, ZN => n1262);
   U1335 : OAI221_X1 port map( B1 => n2140, B2 => n2682, C1 => n2136, C2 => 
                           n2618, A => n1264, ZN => n1263);
   U1336 : AOI22_X1 port map( A1 => REGISTERS_10_10_port, A2 => n2117, B1 => 
                           REGISTERS_8_10_port, B2 => n2113, ZN => n1265);
   U1337 : OAI21_X1 port map( B1 => n1247, B2 => n1248, A => n2144, ZN => n1246
                           );
   U1338 : OAI221_X1 port map( B1 => n2124, B2 => n2649, C1 => n2120, C2 => 
                           n2585, A => n1250, ZN => n1247);
   U1339 : OAI221_X1 port map( B1 => n2140, B2 => n2681, C1 => n2136, C2 => 
                           n2617, A => n1249, ZN => n1248);
   U1340 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n2117, B1 => 
                           REGISTERS_8_11_port, B2 => n2113, ZN => n1250);
   U1341 : OAI21_X1 port map( B1 => n1232, B2 => n1233, A => n2145, ZN => n1231
                           );
   U1342 : OAI221_X1 port map( B1 => n2125, B2 => n2648, C1 => n2121, C2 => 
                           n2584, A => n1235, ZN => n1232);
   U1343 : OAI221_X1 port map( B1 => n2141, B2 => n2680, C1 => n2137, C2 => 
                           n2616, A => n1234, ZN => n1233);
   U1344 : AOI22_X1 port map( A1 => REGISTERS_10_12_port, A2 => n2117, B1 => 
                           REGISTERS_8_12_port, B2 => n2113, ZN => n1235);
   U1345 : OAI21_X1 port map( B1 => n1217, B2 => n1218, A => n2145, ZN => n1216
                           );
   U1346 : OAI221_X1 port map( B1 => n2125, B2 => n2647, C1 => n2121, C2 => 
                           n2583, A => n1220, ZN => n1217);
   U1347 : OAI221_X1 port map( B1 => n2141, B2 => n2679, C1 => n2137, C2 => 
                           n2615, A => n1219, ZN => n1218);
   U1348 : AOI22_X1 port map( A1 => REGISTERS_10_13_port, A2 => n2117, B1 => 
                           REGISTERS_8_13_port, B2 => n2113, ZN => n1220);
   U1349 : OAI21_X1 port map( B1 => n1202, B2 => n1203, A => n2145, ZN => n1201
                           );
   U1350 : OAI221_X1 port map( B1 => n2125, B2 => n2646, C1 => n2121, C2 => 
                           n2582, A => n1205, ZN => n1202);
   U1351 : OAI221_X1 port map( B1 => n2141, B2 => n2678, C1 => n2137, C2 => 
                           n2614, A => n1204, ZN => n1203);
   U1352 : AOI22_X1 port map( A1 => REGISTERS_10_14_port, A2 => n2117, B1 => 
                           REGISTERS_8_14_port, B2 => n2113, ZN => n1205);
   U1353 : OAI21_X1 port map( B1 => n1187, B2 => n1188, A => n2145, ZN => n1186
                           );
   U1354 : OAI221_X1 port map( B1 => n2125, B2 => n2645, C1 => n2121, C2 => 
                           n2581, A => n1190, ZN => n1187);
   U1355 : OAI221_X1 port map( B1 => n2141, B2 => n2677, C1 => n2137, C2 => 
                           n2613, A => n1189, ZN => n1188);
   U1356 : AOI22_X1 port map( A1 => REGISTERS_10_15_port, A2 => n2117, B1 => 
                           REGISTERS_8_15_port, B2 => n2113, ZN => n1190);
   U1357 : OAI21_X1 port map( B1 => n1172, B2 => n1173, A => n2145, ZN => n1171
                           );
   U1358 : OAI221_X1 port map( B1 => n2124, B2 => n2644, C1 => n2121, C2 => 
                           n2580, A => n1175, ZN => n1172);
   U1359 : OAI221_X1 port map( B1 => n2140, B2 => n2676, C1 => n2137, C2 => 
                           n2612, A => n1174, ZN => n1173);
   U1360 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n2117, B1 => 
                           REGISTERS_8_16_port, B2 => n2113, ZN => n1175);
   U1361 : OAI21_X1 port map( B1 => n1157, B2 => n1158, A => n2145, ZN => n1156
                           );
   U1362 : OAI221_X1 port map( B1 => n2125, B2 => n2643, C1 => n2121, C2 => 
                           n2579, A => n1160, ZN => n1157);
   U1363 : OAI221_X1 port map( B1 => n2141, B2 => n2675, C1 => n2137, C2 => 
                           n2611, A => n1159, ZN => n1158);
   U1364 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n2117, B1 => 
                           REGISTERS_8_17_port, B2 => n2113, ZN => n1160);
   U1365 : OAI21_X1 port map( B1 => n1142, B2 => n1143, A => n2145, ZN => n1141
                           );
   U1366 : OAI221_X1 port map( B1 => n2124, B2 => n2642, C1 => n2121, C2 => 
                           n2578, A => n1145, ZN => n1142);
   U1367 : OAI221_X1 port map( B1 => n2140, B2 => n2674, C1 => n2137, C2 => 
                           n2610, A => n1144, ZN => n1143);
   U1368 : AOI22_X1 port map( A1 => REGISTERS_10_18_port, A2 => n2117, B1 => 
                           REGISTERS_8_18_port, B2 => n2113, ZN => n1145);
   U1369 : OAI21_X1 port map( B1 => n1127, B2 => n1128, A => n2145, ZN => n1126
                           );
   U1370 : OAI221_X1 port map( B1 => n2125, B2 => n2641, C1 => n2121, C2 => 
                           n2577, A => n1130, ZN => n1127);
   U1371 : OAI221_X1 port map( B1 => n2141, B2 => n2673, C1 => n2137, C2 => 
                           n2609, A => n1129, ZN => n1128);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_10_19_port, A2 => n2116, B1 => 
                           REGISTERS_8_19_port, B2 => n2113, ZN => n1130);
   U1373 : OAI21_X1 port map( B1 => n1112, B2 => n1113, A => n2145, ZN => n1111
                           );
   U1374 : OAI221_X1 port map( B1 => n2124, B2 => n2640, C1 => n2121, C2 => 
                           n2576, A => n1115, ZN => n1112);
   U1375 : OAI221_X1 port map( B1 => n2140, B2 => n2672, C1 => n2137, C2 => 
                           n2608, A => n1114, ZN => n1113);
   U1376 : AOI22_X1 port map( A1 => REGISTERS_10_20_port, A2 => n2116, B1 => 
                           REGISTERS_8_20_port, B2 => n2113, ZN => n1115);
   U1377 : OAI21_X1 port map( B1 => n1097, B2 => n1098, A => n2145, ZN => n1096
                           );
   U1378 : OAI221_X1 port map( B1 => n2125, B2 => n2639, C1 => n2121, C2 => 
                           n2575, A => n1100, ZN => n1097);
   U1379 : OAI221_X1 port map( B1 => n2141, B2 => n2671, C1 => n2137, C2 => 
                           n2607, A => n1099, ZN => n1098);
   U1380 : AOI22_X1 port map( A1 => REGISTERS_10_21_port, A2 => n2116, B1 => 
                           REGISTERS_8_21_port, B2 => n2112, ZN => n1100);
   U1381 : OAI21_X1 port map( B1 => n1082, B2 => n1083, A => n2145, ZN => n1081
                           );
   U1382 : OAI221_X1 port map( B1 => n2124, B2 => n2638, C1 => n2121, C2 => 
                           n2574, A => n1085, ZN => n1082);
   U1383 : OAI221_X1 port map( B1 => n2140, B2 => n2670, C1 => n2137, C2 => 
                           n2606, A => n1084, ZN => n1083);
   U1384 : AOI22_X1 port map( A1 => REGISTERS_10_22_port, A2 => n2116, B1 => 
                           REGISTERS_8_22_port, B2 => n2112, ZN => n1085);
   U1385 : OAI21_X1 port map( B1 => n1067, B2 => n1068, A => n2145, ZN => n1066
                           );
   U1386 : OAI221_X1 port map( B1 => n2125, B2 => n2637, C1 => n2121, C2 => 
                           n2573, A => n1070, ZN => n1067);
   U1387 : OAI221_X1 port map( B1 => n2141, B2 => n2669, C1 => n2137, C2 => 
                           n2605, A => n1069, ZN => n1068);
   U1388 : AOI22_X1 port map( A1 => REGISTERS_10_23_port, A2 => n2116, B1 => 
                           REGISTERS_8_23_port, B2 => n2112, ZN => n1070);
   U1389 : OAI21_X1 port map( B1 => n1052, B2 => n1053, A => n2146, ZN => n1051
                           );
   U1390 : OAI221_X1 port map( B1 => n2125, B2 => n2636, C1 => n2120, C2 => 
                           n2572, A => n1055, ZN => n1052);
   U1391 : OAI221_X1 port map( B1 => n2141, B2 => n2668, C1 => n2136, C2 => 
                           n2604, A => n1054, ZN => n1053);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_10_24_port, A2 => n2116, B1 => 
                           REGISTERS_8_24_port, B2 => n2112, ZN => n1055);
   U1393 : OAI21_X1 port map( B1 => n1037, B2 => n1038, A => n2146, ZN => n1036
                           );
   U1394 : OAI221_X1 port map( B1 => n2125, B2 => n2635, C1 => n2121, C2 => 
                           n2571, A => n1040, ZN => n1037);
   U1395 : OAI221_X1 port map( B1 => n2141, B2 => n2667, C1 => n2137, C2 => 
                           n2603, A => n1039, ZN => n1038);
   U1396 : AOI22_X1 port map( A1 => REGISTERS_10_25_port, A2 => n2116, B1 => 
                           REGISTERS_8_25_port, B2 => n2112, ZN => n1040);
   U1397 : OAI21_X1 port map( B1 => n1022, B2 => n1023, A => n2146, ZN => n1021
                           );
   U1398 : OAI221_X1 port map( B1 => n2125, B2 => n2634, C1 => n2120, C2 => 
                           n2570, A => n1025, ZN => n1022);
   U1399 : OAI221_X1 port map( B1 => n2141, B2 => n2666, C1 => n2136, C2 => 
                           n2602, A => n1024, ZN => n1023);
   U1400 : AOI22_X1 port map( A1 => REGISTERS_10_26_port, A2 => n2116, B1 => 
                           REGISTERS_8_26_port, B2 => n2112, ZN => n1025);
   U1401 : OAI21_X1 port map( B1 => n1007, B2 => n1008, A => n2146, ZN => n1006
                           );
   U1402 : OAI221_X1 port map( B1 => n2125, B2 => n2633, C1 => n2121, C2 => 
                           n2569, A => n1010, ZN => n1007);
   U1403 : OAI221_X1 port map( B1 => n2141, B2 => n2665, C1 => n2137, C2 => 
                           n2601, A => n1009, ZN => n1008);
   U1404 : AOI22_X1 port map( A1 => REGISTERS_10_27_port, A2 => n2116, B1 => 
                           REGISTERS_8_27_port, B2 => n2112, ZN => n1010);
   U1405 : OAI21_X1 port map( B1 => n992, B2 => n993, A => n2146, ZN => n991);
   U1406 : OAI221_X1 port map( B1 => n2125, B2 => n2632, C1 => n2120, C2 => 
                           n2568, A => n995, ZN => n992);
   U1407 : OAI221_X1 port map( B1 => n2141, B2 => n2664, C1 => n2136, C2 => 
                           n2600, A => n994, ZN => n993);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_10_28_port, A2 => n2116, B1 => 
                           REGISTERS_8_28_port, B2 => n2112, ZN => n995);
   U1409 : OAI21_X1 port map( B1 => n977, B2 => n978, A => n2146, ZN => n976);
   U1410 : OAI221_X1 port map( B1 => n2125, B2 => n2631, C1 => n2121, C2 => 
                           n2567, A => n980, ZN => n977);
   U1411 : OAI221_X1 port map( B1 => n2141, B2 => n2663, C1 => n2137, C2 => 
                           n2599, A => n979, ZN => n978);
   U1412 : AOI22_X1 port map( A1 => REGISTERS_10_29_port, A2 => n2116, B1 => 
                           REGISTERS_8_29_port, B2 => n2112, ZN => n980);
   U1413 : OAI21_X1 port map( B1 => n962, B2 => n963, A => n2146, ZN => n961);
   U1414 : OAI221_X1 port map( B1 => n2125, B2 => n2630, C1 => n2120, C2 => 
                           n2566, A => n965, ZN => n962);
   U1415 : OAI221_X1 port map( B1 => n2141, B2 => n2662, C1 => n2136, C2 => 
                           n2598, A => n964, ZN => n963);
   U1416 : AOI22_X1 port map( A1 => REGISTERS_10_30_port, A2 => n2116, B1 => 
                           REGISTERS_8_30_port, B2 => n2112, ZN => n965);
   U1417 : OAI21_X1 port map( B1 => n929, B2 => n930, A => n2146, ZN => n928);
   U1418 : OAI221_X1 port map( B1 => n2125, B2 => n2629, C1 => n2121, C2 => 
                           n2565, A => n939, ZN => n929);
   U1419 : OAI221_X1 port map( B1 => n2141, B2 => n2661, C1 => n2137, C2 => 
                           n2597, A => n934, ZN => n930);
   U1420 : AOI22_X1 port map( A1 => REGISTERS_10_31_port, A2 => n2117, B1 => 
                           REGISTERS_8_31_port, B2 => n2113, ZN => n939);
   U1421 : OAI21_X1 port map( B1 => n1929, B2 => n1930, A => n2016, ZN => n1928
                           );
   U1422 : OAI221_X1 port map( B1 => n2660, B2 => n1996, C1 => n2596, C2 => 
                           n1992, A => n1932, ZN => n1929);
   U1423 : OAI221_X1 port map( B1 => n2692, B2 => n2012, C1 => n2628, C2 => 
                           n2008, A => n1931, ZN => n1930);
   U1424 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_0_port, B1 => 
                           n1984, B2 => REGISTERS_8_0_port, ZN => n1932);
   U1425 : OAI21_X1 port map( B1 => n1912, B2 => n1913, A => n2016, ZN => n1911
                           );
   U1426 : OAI221_X1 port map( B1 => n2659, B2 => n1996, C1 => n2595, C2 => 
                           n1992, A => n1915, ZN => n1912);
   U1427 : OAI221_X1 port map( B1 => n2691, B2 => n2012, C1 => n2627, C2 => 
                           n2008, A => n1914, ZN => n1913);
   U1428 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_1_port, B1 => 
                           n1986, B2 => REGISTERS_8_1_port, ZN => n1915);
   U1429 : OAI21_X1 port map( B1 => n1897, B2 => n1898, A => n2016, ZN => n1896
                           );
   U1430 : OAI221_X1 port map( B1 => n2658, B2 => n1996, C1 => n2594, C2 => 
                           n1992, A => n1900, ZN => n1897);
   U1431 : OAI221_X1 port map( B1 => n2690, B2 => n2012, C1 => n2626, C2 => 
                           n2008, A => n1899, ZN => n1898);
   U1432 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_2_port, B1 => 
                           n1986, B2 => REGISTERS_8_2_port, ZN => n1900);
   U1433 : OAI21_X1 port map( B1 => n1882, B2 => n1883, A => n2016, ZN => n1881
                           );
   U1434 : OAI221_X1 port map( B1 => n2657, B2 => n1996, C1 => n2593, C2 => 
                           n1992, A => n1885, ZN => n1882);
   U1435 : OAI221_X1 port map( B1 => n2689, B2 => n2012, C1 => n2625, C2 => 
                           n2008, A => n1884, ZN => n1883);
   U1436 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_3_port, B1 => 
                           n1986, B2 => REGISTERS_8_3_port, ZN => n1885);
   U1437 : OAI21_X1 port map( B1 => n1867, B2 => n1868, A => n2016, ZN => n1866
                           );
   U1438 : OAI221_X1 port map( B1 => n2656, B2 => n1996, C1 => n2592, C2 => 
                           n1992, A => n1870, ZN => n1867);
   U1439 : OAI221_X1 port map( B1 => n2688, B2 => n2012, C1 => n2624, C2 => 
                           n2008, A => n1869, ZN => n1868);
   U1440 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_4_port, B1 => 
                           n1986, B2 => REGISTERS_8_4_port, ZN => n1870);
   U1441 : OAI21_X1 port map( B1 => n1852, B2 => n1853, A => n2016, ZN => n1851
                           );
   U1442 : OAI221_X1 port map( B1 => n2655, B2 => n1996, C1 => n2591, C2 => 
                           n1992, A => n1855, ZN => n1852);
   U1443 : OAI221_X1 port map( B1 => n2687, B2 => n2012, C1 => n2623, C2 => 
                           n2008, A => n1854, ZN => n1853);
   U1444 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_5_port, B1 => 
                           n1986, B2 => REGISTERS_8_5_port, ZN => n1855);
   U1445 : OAI21_X1 port map( B1 => n1837, B2 => n1838, A => n2016, ZN => n1836
                           );
   U1446 : OAI221_X1 port map( B1 => n2654, B2 => n1996, C1 => n2590, C2 => 
                           n1992, A => n1840, ZN => n1837);
   U1447 : OAI221_X1 port map( B1 => n2686, B2 => n2012, C1 => n2622, C2 => 
                           n2008, A => n1839, ZN => n1838);
   U1448 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_6_port, B1 => 
                           n1986, B2 => REGISTERS_8_6_port, ZN => n1840);
   U1449 : OAI21_X1 port map( B1 => n1822, B2 => n1823, A => n2016, ZN => n1821
                           );
   U1450 : OAI221_X1 port map( B1 => n2653, B2 => n1996, C1 => n2589, C2 => 
                           n1992, A => n1825, ZN => n1822);
   U1451 : OAI221_X1 port map( B1 => n2685, B2 => n2012, C1 => n2621, C2 => 
                           n2008, A => n1824, ZN => n1823);
   U1452 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_7_port, B1 => 
                           n1986, B2 => REGISTERS_8_7_port, ZN => n1825);
   U1453 : OAI21_X1 port map( B1 => n1807, B2 => n1808, A => n2016, ZN => n1806
                           );
   U1454 : OAI221_X1 port map( B1 => n2652, B2 => n1996, C1 => n2588, C2 => 
                           n1992, A => n1810, ZN => n1807);
   U1455 : OAI221_X1 port map( B1 => n2684, B2 => n2012, C1 => n2620, C2 => 
                           n2008, A => n1809, ZN => n1808);
   U1456 : AOI22_X1 port map( A1 => n1990, A2 => REGISTERS_10_8_port, B1 => 
                           n1986, B2 => REGISTERS_8_8_port, ZN => n1810);
   U1457 : OAI21_X1 port map( B1 => n1792, B2 => n1793, A => n2016, ZN => n1791
                           );
   U1458 : OAI221_X1 port map( B1 => n2651, B2 => n1996, C1 => n2587, C2 => 
                           n1992, A => n1795, ZN => n1792);
   U1459 : OAI221_X1 port map( B1 => n2683, B2 => n2012, C1 => n2619, C2 => 
                           n2008, A => n1794, ZN => n1793);
   U1460 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_9_port, B1 => 
                           n1985, B2 => REGISTERS_8_9_port, ZN => n1795);
   U1461 : OAI21_X1 port map( B1 => n1777, B2 => n1778, A => n2016, ZN => n1776
                           );
   U1462 : OAI221_X1 port map( B1 => n2650, B2 => n1996, C1 => n2586, C2 => 
                           n1992, A => n1780, ZN => n1777);
   U1463 : OAI221_X1 port map( B1 => n2682, B2 => n2012, C1 => n2618, C2 => 
                           n2008, A => n1779, ZN => n1778);
   U1464 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_10_port, B1 => 
                           n1985, B2 => REGISTERS_8_10_port, ZN => n1780);
   U1465 : OAI21_X1 port map( B1 => n1762, B2 => n1763, A => n2016, ZN => n1761
                           );
   U1466 : OAI221_X1 port map( B1 => n2649, B2 => n1996, C1 => n2585, C2 => 
                           n1992, A => n1765, ZN => n1762);
   U1467 : OAI221_X1 port map( B1 => n2681, B2 => n2012, C1 => n2617, C2 => 
                           n2008, A => n1764, ZN => n1763);
   U1468 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_11_port, B1 => 
                           n1985, B2 => REGISTERS_8_11_port, ZN => n1765);
   U1469 : OAI21_X1 port map( B1 => n1747, B2 => n1748, A => n2017, ZN => n1746
                           );
   U1470 : OAI221_X1 port map( B1 => n2648, B2 => n1997, C1 => n2584, C2 => 
                           n1993, A => n1750, ZN => n1747);
   U1471 : OAI221_X1 port map( B1 => n2680, B2 => n2013, C1 => n2616, C2 => 
                           n2009, A => n1749, ZN => n1748);
   U1472 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_12_port, B1 => 
                           n1985, B2 => REGISTERS_8_12_port, ZN => n1750);
   U1473 : OAI21_X1 port map( B1 => n1732, B2 => n1733, A => n2017, ZN => n1731
                           );
   U1474 : OAI221_X1 port map( B1 => n2647, B2 => n1997, C1 => n2583, C2 => 
                           n1993, A => n1735, ZN => n1732);
   U1475 : OAI221_X1 port map( B1 => n2679, B2 => n2013, C1 => n2615, C2 => 
                           n2009, A => n1734, ZN => n1733);
   U1476 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_13_port, B1 => 
                           n1985, B2 => REGISTERS_8_13_port, ZN => n1735);
   U1477 : OAI21_X1 port map( B1 => n1717, B2 => n1718, A => n2017, ZN => n1716
                           );
   U1478 : OAI221_X1 port map( B1 => n2646, B2 => n1997, C1 => n2582, C2 => 
                           n1993, A => n1720, ZN => n1717);
   U1479 : OAI221_X1 port map( B1 => n2678, B2 => n2013, C1 => n2614, C2 => 
                           n2009, A => n1719, ZN => n1718);
   U1480 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_14_port, B1 => 
                           n1985, B2 => REGISTERS_8_14_port, ZN => n1720);
   U1481 : OAI21_X1 port map( B1 => n1702, B2 => n1703, A => n2017, ZN => n1701
                           );
   U1482 : OAI221_X1 port map( B1 => n2645, B2 => n1997, C1 => n2581, C2 => 
                           n1993, A => n1705, ZN => n1702);
   U1483 : OAI221_X1 port map( B1 => n2677, B2 => n2013, C1 => n2613, C2 => 
                           n2009, A => n1704, ZN => n1703);
   U1484 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_15_port, B1 => 
                           n1985, B2 => REGISTERS_8_15_port, ZN => n1705);
   U1485 : OAI21_X1 port map( B1 => n1687, B2 => n1688, A => n2017, ZN => n1686
                           );
   U1486 : OAI221_X1 port map( B1 => n2644, B2 => n1996, C1 => n2580, C2 => 
                           n1993, A => n1690, ZN => n1687);
   U1487 : OAI221_X1 port map( B1 => n2676, B2 => n2012, C1 => n2612, C2 => 
                           n2009, A => n1689, ZN => n1688);
   U1488 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_16_port, B1 => 
                           n1985, B2 => REGISTERS_8_16_port, ZN => n1690);
   U1489 : OAI21_X1 port map( B1 => n1672, B2 => n1673, A => n2017, ZN => n1671
                           );
   U1490 : OAI221_X1 port map( B1 => n2643, B2 => n1997, C1 => n2579, C2 => 
                           n1993, A => n1675, ZN => n1672);
   U1491 : OAI221_X1 port map( B1 => n2675, B2 => n2013, C1 => n2611, C2 => 
                           n2009, A => n1674, ZN => n1673);
   U1492 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_17_port, B1 => 
                           n1985, B2 => REGISTERS_8_17_port, ZN => n1675);
   U1493 : OAI21_X1 port map( B1 => n1657, B2 => n1658, A => n2017, ZN => n1656
                           );
   U1494 : OAI221_X1 port map( B1 => n2642, B2 => n1996, C1 => n2578, C2 => 
                           n1993, A => n1660, ZN => n1657);
   U1495 : OAI221_X1 port map( B1 => n2674, B2 => n2012, C1 => n2610, C2 => 
                           n2009, A => n1659, ZN => n1658);
   U1496 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_18_port, B1 => 
                           n1985, B2 => REGISTERS_8_18_port, ZN => n1660);
   U1497 : OAI21_X1 port map( B1 => n1642, B2 => n1643, A => n2017, ZN => n1641
                           );
   U1498 : OAI221_X1 port map( B1 => n2641, B2 => n1997, C1 => n2577, C2 => 
                           n1993, A => n1645, ZN => n1642);
   U1499 : OAI221_X1 port map( B1 => n2673, B2 => n2013, C1 => n2609, C2 => 
                           n2009, A => n1644, ZN => n1643);
   U1500 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_19_port, B1 => 
                           n1985, B2 => REGISTERS_8_19_port, ZN => n1645);
   U1501 : OAI21_X1 port map( B1 => n1627, B2 => n1628, A => n2017, ZN => n1626
                           );
   U1502 : OAI221_X1 port map( B1 => n2640, B2 => n1996, C1 => n2576, C2 => 
                           n1993, A => n1630, ZN => n1627);
   U1503 : OAI221_X1 port map( B1 => n2672, B2 => n2012, C1 => n2608, C2 => 
                           n2009, A => n1629, ZN => n1628);
   U1504 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_20_port, B1 => 
                           n1985, B2 => REGISTERS_8_20_port, ZN => n1630);
   U1505 : OAI21_X1 port map( B1 => n1612, B2 => n1613, A => n2017, ZN => n1611
                           );
   U1506 : OAI221_X1 port map( B1 => n2639, B2 => n1997, C1 => n2575, C2 => 
                           n1993, A => n1615, ZN => n1612);
   U1507 : OAI221_X1 port map( B1 => n2671, B2 => n2013, C1 => n2607, C2 => 
                           n2009, A => n1614, ZN => n1613);
   U1508 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_21_port, B1 => 
                           n1984, B2 => REGISTERS_8_21_port, ZN => n1615);
   U1509 : OAI21_X1 port map( B1 => n1597, B2 => n1598, A => n2017, ZN => n1596
                           );
   U1510 : OAI221_X1 port map( B1 => n2638, B2 => n1996, C1 => n2574, C2 => 
                           n1993, A => n1600, ZN => n1597);
   U1511 : OAI221_X1 port map( B1 => n2670, B2 => n2012, C1 => n2606, C2 => 
                           n2009, A => n1599, ZN => n1598);
   U1512 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_22_port, B1 => 
                           n1984, B2 => REGISTERS_8_22_port, ZN => n1600);
   U1513 : OAI21_X1 port map( B1 => n1582, B2 => n1583, A => n2017, ZN => n1581
                           );
   U1514 : OAI221_X1 port map( B1 => n2637, B2 => n1997, C1 => n2573, C2 => 
                           n1993, A => n1585, ZN => n1582);
   U1515 : OAI221_X1 port map( B1 => n2669, B2 => n2013, C1 => n2605, C2 => 
                           n2009, A => n1584, ZN => n1583);
   U1516 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_23_port, B1 => 
                           n1984, B2 => REGISTERS_8_23_port, ZN => n1585);
   U1517 : OAI21_X1 port map( B1 => n1567, B2 => n1568, A => n2018, ZN => n1566
                           );
   U1518 : OAI221_X1 port map( B1 => n2636, B2 => n1997, C1 => n2572, C2 => 
                           n1992, A => n1570, ZN => n1567);
   U1519 : OAI221_X1 port map( B1 => n2668, B2 => n2013, C1 => n2604, C2 => 
                           n2008, A => n1569, ZN => n1568);
   U1520 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_24_port, B1 => 
                           n1984, B2 => REGISTERS_8_24_port, ZN => n1570);
   U1521 : OAI21_X1 port map( B1 => n1552, B2 => n1553, A => n2018, ZN => n1551
                           );
   U1522 : OAI221_X1 port map( B1 => n2635, B2 => n1997, C1 => n2571, C2 => 
                           n1993, A => n1555, ZN => n1552);
   U1523 : OAI221_X1 port map( B1 => n2667, B2 => n2013, C1 => n2603, C2 => 
                           n2009, A => n1554, ZN => n1553);
   U1524 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_25_port, B1 => 
                           n1984, B2 => REGISTERS_8_25_port, ZN => n1555);
   U1525 : OAI21_X1 port map( B1 => n1537, B2 => n1538, A => n2018, ZN => n1536
                           );
   U1526 : OAI221_X1 port map( B1 => n2634, B2 => n1997, C1 => n2570, C2 => 
                           n1992, A => n1540, ZN => n1537);
   U1527 : OAI221_X1 port map( B1 => n2666, B2 => n2013, C1 => n2602, C2 => 
                           n2008, A => n1539, ZN => n1538);
   U1528 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_26_port, B1 => 
                           n1984, B2 => REGISTERS_8_26_port, ZN => n1540);
   U1529 : OAI21_X1 port map( B1 => n1522, B2 => n1523, A => n2018, ZN => n1521
                           );
   U1530 : OAI221_X1 port map( B1 => n2633, B2 => n1997, C1 => n2569, C2 => 
                           n1993, A => n1525, ZN => n1522);
   U1531 : OAI221_X1 port map( B1 => n2665, B2 => n2013, C1 => n2601, C2 => 
                           n2009, A => n1524, ZN => n1523);
   U1532 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_27_port, B1 => 
                           n1984, B2 => REGISTERS_8_27_port, ZN => n1525);
   U1533 : OAI21_X1 port map( B1 => n1507, B2 => n1508, A => n2018, ZN => n1506
                           );
   U1534 : OAI221_X1 port map( B1 => n2632, B2 => n1997, C1 => n2568, C2 => 
                           n1992, A => n1510, ZN => n1507);
   U1535 : OAI221_X1 port map( B1 => n2664, B2 => n2013, C1 => n2600, C2 => 
                           n2008, A => n1509, ZN => n1508);
   U1536 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_28_port, B1 => 
                           n1984, B2 => REGISTERS_8_28_port, ZN => n1510);
   U1537 : OAI21_X1 port map( B1 => n1492, B2 => n1493, A => n2018, ZN => n1491
                           );
   U1538 : OAI221_X1 port map( B1 => n2631, B2 => n1997, C1 => n2567, C2 => 
                           n1993, A => n1495, ZN => n1492);
   U1539 : OAI221_X1 port map( B1 => n2663, B2 => n2013, C1 => n2599, C2 => 
                           n2009, A => n1494, ZN => n1493);
   U1540 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_29_port, B1 => 
                           n1984, B2 => REGISTERS_8_29_port, ZN => n1495);
   U1541 : OAI21_X1 port map( B1 => n1477, B2 => n1478, A => n2018, ZN => n1476
                           );
   U1542 : OAI221_X1 port map( B1 => n2630, B2 => n1997, C1 => n2566, C2 => 
                           n1992, A => n1480, ZN => n1477);
   U1543 : OAI221_X1 port map( B1 => n2662, B2 => n2013, C1 => n2598, C2 => 
                           n2008, A => n1479, ZN => n1478);
   U1544 : AOI22_X1 port map( A1 => n1988, A2 => REGISTERS_10_30_port, B1 => 
                           n1984, B2 => REGISTERS_8_30_port, ZN => n1480);
   U1545 : OAI21_X1 port map( B1 => n1444, B2 => n1445, A => n2018, ZN => n1443
                           );
   U1546 : OAI221_X1 port map( B1 => n2629, B2 => n1997, C1 => n2565, C2 => 
                           n1993, A => n1454, ZN => n1444);
   U1547 : OAI221_X1 port map( B1 => n2661, B2 => n2013, C1 => n2597, C2 => 
                           n2009, A => n1449, ZN => n1445);
   U1548 : AOI22_X1 port map( A1 => n1989, A2 => REGISTERS_10_31_port, B1 => 
                           n1985, B2 => REGISTERS_8_31_port, ZN => n1454);
   U1549 : INV_X1 port map( A => ADD_RD2(0), ZN => n3219);
   U1550 : AND3_X1 port map( A1 => ENABLE, A2 => n3220, A3 => WR, ZN => n899);
   U1551 : INV_X1 port map( A => ADD_RD1(3), ZN => n3213);
   U1552 : INV_X1 port map( A => ADD_WR(0), ZN => n3211);
   U1553 : INV_X1 port map( A => ADD_WR(2), ZN => n3209);
   U1554 : INV_X1 port map( A => ADD_WR(1), ZN => n3210);
   U1555 : NOR3_X1 port map( A1 => n3214, A2 => ADD_RD1(2), A3 => n3215, ZN => 
                           n1450);
   U1556 : INV_X1 port map( A => REGISTERS_15_0_port, ZN => n2692);
   U1557 : INV_X1 port map( A => REGISTERS_14_0_port, ZN => n2660);
   U1558 : INV_X1 port map( A => REGISTERS_15_1_port, ZN => n2691);
   U1559 : INV_X1 port map( A => REGISTERS_14_1_port, ZN => n2659);
   U1560 : INV_X1 port map( A => REGISTERS_15_2_port, ZN => n2690);
   U1561 : INV_X1 port map( A => REGISTERS_14_2_port, ZN => n2658);
   U1562 : INV_X1 port map( A => REGISTERS_15_3_port, ZN => n2689);
   U1563 : INV_X1 port map( A => REGISTERS_14_3_port, ZN => n2657);
   U1564 : INV_X1 port map( A => REGISTERS_15_4_port, ZN => n2688);
   U1565 : INV_X1 port map( A => REGISTERS_14_4_port, ZN => n2656);
   U1566 : INV_X1 port map( A => REGISTERS_15_5_port, ZN => n2687);
   U1567 : INV_X1 port map( A => REGISTERS_14_5_port, ZN => n2655);
   U1568 : INV_X1 port map( A => REGISTERS_15_6_port, ZN => n2686);
   U1569 : INV_X1 port map( A => REGISTERS_14_6_port, ZN => n2654);
   U1570 : INV_X1 port map( A => REGISTERS_15_7_port, ZN => n2685);
   U1571 : INV_X1 port map( A => REGISTERS_14_7_port, ZN => n2653);
   U1572 : INV_X1 port map( A => REGISTERS_15_8_port, ZN => n2684);
   U1573 : INV_X1 port map( A => REGISTERS_14_8_port, ZN => n2652);
   U1574 : INV_X1 port map( A => REGISTERS_15_9_port, ZN => n2683);
   U1575 : INV_X1 port map( A => REGISTERS_14_9_port, ZN => n2651);
   U1576 : INV_X1 port map( A => REGISTERS_15_10_port, ZN => n2682);
   U1577 : INV_X1 port map( A => REGISTERS_14_10_port, ZN => n2650);
   U1578 : INV_X1 port map( A => REGISTERS_15_11_port, ZN => n2681);
   U1579 : INV_X1 port map( A => REGISTERS_14_11_port, ZN => n2649);
   U1580 : INV_X1 port map( A => REGISTERS_15_12_port, ZN => n2680);
   U1581 : INV_X1 port map( A => REGISTERS_14_12_port, ZN => n2648);
   U1582 : INV_X1 port map( A => REGISTERS_15_13_port, ZN => n2679);
   U1583 : INV_X1 port map( A => REGISTERS_14_13_port, ZN => n2647);
   U1584 : INV_X1 port map( A => REGISTERS_15_14_port, ZN => n2678);
   U1585 : INV_X1 port map( A => REGISTERS_14_14_port, ZN => n2646);
   U1586 : INV_X1 port map( A => REGISTERS_15_15_port, ZN => n2677);
   U1587 : INV_X1 port map( A => REGISTERS_14_15_port, ZN => n2645);
   U1588 : INV_X1 port map( A => REGISTERS_15_16_port, ZN => n2676);
   U1589 : INV_X1 port map( A => REGISTERS_14_16_port, ZN => n2644);
   U1590 : INV_X1 port map( A => REGISTERS_15_17_port, ZN => n2675);
   U1591 : INV_X1 port map( A => REGISTERS_14_17_port, ZN => n2643);
   U1592 : INV_X1 port map( A => REGISTERS_15_18_port, ZN => n2674);
   U1593 : INV_X1 port map( A => REGISTERS_14_18_port, ZN => n2642);
   U1594 : INV_X1 port map( A => REGISTERS_15_19_port, ZN => n2673);
   U1595 : INV_X1 port map( A => REGISTERS_14_19_port, ZN => n2641);
   U1596 : INV_X1 port map( A => REGISTERS_15_20_port, ZN => n2672);
   U1597 : INV_X1 port map( A => REGISTERS_14_20_port, ZN => n2640);
   U1598 : INV_X1 port map( A => REGISTERS_15_21_port, ZN => n2671);
   U1599 : INV_X1 port map( A => REGISTERS_14_21_port, ZN => n2639);
   U1600 : INV_X1 port map( A => REGISTERS_15_22_port, ZN => n2670);
   U1601 : INV_X1 port map( A => REGISTERS_14_22_port, ZN => n2638);
   U1602 : INV_X1 port map( A => REGISTERS_15_23_port, ZN => n2669);
   U1603 : INV_X1 port map( A => REGISTERS_14_23_port, ZN => n2637);
   U1604 : INV_X1 port map( A => REGISTERS_15_24_port, ZN => n2668);
   U1605 : INV_X1 port map( A => REGISTERS_14_24_port, ZN => n2636);
   U1606 : INV_X1 port map( A => REGISTERS_15_25_port, ZN => n2667);
   U1607 : INV_X1 port map( A => REGISTERS_14_25_port, ZN => n2635);
   U1608 : INV_X1 port map( A => REGISTERS_15_26_port, ZN => n2666);
   U1609 : INV_X1 port map( A => REGISTERS_14_26_port, ZN => n2634);
   U1610 : INV_X1 port map( A => REGISTERS_15_27_port, ZN => n2665);
   U1611 : INV_X1 port map( A => REGISTERS_14_27_port, ZN => n2633);
   U1612 : INV_X1 port map( A => REGISTERS_15_28_port, ZN => n2664);
   U1613 : INV_X1 port map( A => REGISTERS_14_28_port, ZN => n2632);
   U1614 : INV_X1 port map( A => REGISTERS_15_29_port, ZN => n2663);
   U1615 : INV_X1 port map( A => REGISTERS_14_29_port, ZN => n2631);
   U1616 : INV_X1 port map( A => REGISTERS_15_30_port, ZN => n2662);
   U1617 : INV_X1 port map( A => REGISTERS_14_30_port, ZN => n2630);
   U1618 : INV_X1 port map( A => REGISTERS_15_31_port, ZN => n2661);
   U1619 : INV_X1 port map( A => REGISTERS_14_31_port, ZN => n2629);
   U1620 : INV_X1 port map( A => REGISTERS_23_0_port, ZN => n2948);
   U1621 : INV_X1 port map( A => REGISTERS_23_1_port, ZN => n2947);
   U1622 : INV_X1 port map( A => REGISTERS_23_2_port, ZN => n2946);
   U1623 : INV_X1 port map( A => REGISTERS_23_3_port, ZN => n2945);
   U1624 : INV_X1 port map( A => REGISTERS_23_4_port, ZN => n2944);
   U1625 : INV_X1 port map( A => REGISTERS_23_5_port, ZN => n2943);
   U1626 : INV_X1 port map( A => REGISTERS_23_6_port, ZN => n2942);
   U1627 : INV_X1 port map( A => REGISTERS_23_7_port, ZN => n2941);
   U1628 : INV_X1 port map( A => REGISTERS_23_8_port, ZN => n2940);
   U1629 : INV_X1 port map( A => REGISTERS_23_9_port, ZN => n2939);
   U1630 : INV_X1 port map( A => REGISTERS_23_10_port, ZN => n2938);
   U1631 : INV_X1 port map( A => REGISTERS_23_11_port, ZN => n2937);
   U1632 : INV_X1 port map( A => REGISTERS_23_12_port, ZN => n2936);
   U1633 : INV_X1 port map( A => REGISTERS_23_13_port, ZN => n2935);
   U1634 : INV_X1 port map( A => REGISTERS_23_14_port, ZN => n2934);
   U1635 : INV_X1 port map( A => REGISTERS_23_15_port, ZN => n2933);
   U1636 : INV_X1 port map( A => REGISTERS_23_16_port, ZN => n2932);
   U1637 : INV_X1 port map( A => REGISTERS_23_17_port, ZN => n2931);
   U1638 : INV_X1 port map( A => REGISTERS_23_18_port, ZN => n2930);
   U1639 : INV_X1 port map( A => REGISTERS_23_19_port, ZN => n2929);
   U1640 : INV_X1 port map( A => REGISTERS_23_20_port, ZN => n2928);
   U1641 : INV_X1 port map( A => REGISTERS_23_21_port, ZN => n2927);
   U1642 : INV_X1 port map( A => REGISTERS_23_22_port, ZN => n2926);
   U1643 : INV_X1 port map( A => REGISTERS_23_23_port, ZN => n2925);
   U1644 : INV_X1 port map( A => REGISTERS_23_24_port, ZN => n2924);
   U1645 : INV_X1 port map( A => REGISTERS_23_25_port, ZN => n2923);
   U1646 : INV_X1 port map( A => REGISTERS_23_26_port, ZN => n2922);
   U1647 : INV_X1 port map( A => REGISTERS_23_27_port, ZN => n2921);
   U1648 : INV_X1 port map( A => REGISTERS_23_28_port, ZN => n2920);
   U1649 : INV_X1 port map( A => REGISTERS_23_29_port, ZN => n2919);
   U1650 : INV_X1 port map( A => REGISTERS_23_30_port, ZN => n2918);
   U1651 : INV_X1 port map( A => REGISTERS_23_31_port, ZN => n2917);
   U1652 : INV_X1 port map( A => REGISTERS_7_0_port, ZN => n2564);
   U1653 : INV_X1 port map( A => REGISTERS_27_0_port, ZN => n3076);
   U1654 : INV_X1 port map( A => REGISTERS_4_0_port, ZN => n2468);
   U1655 : INV_X1 port map( A => REGISTERS_24_0_port, ZN => n2980);
   U1656 : INV_X1 port map( A => REGISTERS_17_0_port, ZN => n2756);
   U1657 : INV_X1 port map( A => REGISTERS_22_0_port, ZN => n2916);
   U1658 : INV_X1 port map( A => REGISTERS_29_0_port, ZN => n3140);
   U1659 : INV_X1 port map( A => REGISTERS_7_1_port, ZN => n2563);
   U1660 : INV_X1 port map( A => REGISTERS_27_1_port, ZN => n3075);
   U1661 : INV_X1 port map( A => REGISTERS_4_1_port, ZN => n2467);
   U1662 : INV_X1 port map( A => REGISTERS_24_1_port, ZN => n2979);
   U1663 : INV_X1 port map( A => REGISTERS_17_1_port, ZN => n2755);
   U1664 : INV_X1 port map( A => REGISTERS_22_1_port, ZN => n2915);
   U1665 : INV_X1 port map( A => REGISTERS_29_1_port, ZN => n3139);
   U1666 : INV_X1 port map( A => REGISTERS_7_2_port, ZN => n2562);
   U1667 : INV_X1 port map( A => REGISTERS_27_2_port, ZN => n3074);
   U1668 : INV_X1 port map( A => REGISTERS_4_2_port, ZN => n2466);
   U1669 : INV_X1 port map( A => REGISTERS_24_2_port, ZN => n2978);
   U1670 : INV_X1 port map( A => REGISTERS_17_2_port, ZN => n2754);
   U1671 : INV_X1 port map( A => REGISTERS_22_2_port, ZN => n2914);
   U1672 : INV_X1 port map( A => REGISTERS_29_2_port, ZN => n3138);
   U1673 : INV_X1 port map( A => REGISTERS_7_3_port, ZN => n2561);
   U1674 : INV_X1 port map( A => REGISTERS_27_3_port, ZN => n3073);
   U1675 : INV_X1 port map( A => REGISTERS_4_3_port, ZN => n2465);
   U1676 : INV_X1 port map( A => REGISTERS_24_3_port, ZN => n2977);
   U1677 : INV_X1 port map( A => REGISTERS_17_3_port, ZN => n2753);
   U1678 : INV_X1 port map( A => REGISTERS_22_3_port, ZN => n2913);
   U1679 : INV_X1 port map( A => REGISTERS_29_3_port, ZN => n3137);
   U1680 : INV_X1 port map( A => REGISTERS_7_4_port, ZN => n2560);
   U1681 : INV_X1 port map( A => REGISTERS_27_4_port, ZN => n3072);
   U1682 : INV_X1 port map( A => REGISTERS_4_4_port, ZN => n2464);
   U1683 : INV_X1 port map( A => REGISTERS_24_4_port, ZN => n2976);
   U1684 : INV_X1 port map( A => REGISTERS_17_4_port, ZN => n2752);
   U1685 : INV_X1 port map( A => REGISTERS_22_4_port, ZN => n2912);
   U1686 : INV_X1 port map( A => REGISTERS_29_4_port, ZN => n3136);
   U1687 : INV_X1 port map( A => REGISTERS_7_5_port, ZN => n2559);
   U1688 : INV_X1 port map( A => REGISTERS_27_5_port, ZN => n3071);
   U1689 : INV_X1 port map( A => REGISTERS_4_5_port, ZN => n2463);
   U1690 : INV_X1 port map( A => REGISTERS_24_5_port, ZN => n2975);
   U1691 : INV_X1 port map( A => REGISTERS_17_5_port, ZN => n2751);
   U1692 : INV_X1 port map( A => REGISTERS_22_5_port, ZN => n2911);
   U1693 : INV_X1 port map( A => REGISTERS_29_5_port, ZN => n3135);
   U1694 : INV_X1 port map( A => REGISTERS_7_6_port, ZN => n2558);
   U1695 : INV_X1 port map( A => REGISTERS_27_6_port, ZN => n3070);
   U1696 : INV_X1 port map( A => REGISTERS_4_6_port, ZN => n2462);
   U1697 : INV_X1 port map( A => REGISTERS_24_6_port, ZN => n2974);
   U1698 : INV_X1 port map( A => REGISTERS_17_6_port, ZN => n2750);
   U1699 : INV_X1 port map( A => REGISTERS_22_6_port, ZN => n2910);
   U1700 : INV_X1 port map( A => REGISTERS_29_6_port, ZN => n3134);
   U1701 : INV_X1 port map( A => REGISTERS_7_7_port, ZN => n2557);
   U1702 : INV_X1 port map( A => REGISTERS_27_7_port, ZN => n3069);
   U1703 : INV_X1 port map( A => REGISTERS_4_7_port, ZN => n2461);
   U1704 : INV_X1 port map( A => REGISTERS_24_7_port, ZN => n2973);
   U1705 : INV_X1 port map( A => REGISTERS_17_7_port, ZN => n2749);
   U1706 : INV_X1 port map( A => REGISTERS_22_7_port, ZN => n2909);
   U1707 : INV_X1 port map( A => REGISTERS_29_7_port, ZN => n3133);
   U1708 : INV_X1 port map( A => REGISTERS_7_8_port, ZN => n2556);
   U1709 : INV_X1 port map( A => REGISTERS_27_8_port, ZN => n3068);
   U1710 : INV_X1 port map( A => REGISTERS_4_8_port, ZN => n2460);
   U1711 : INV_X1 port map( A => REGISTERS_24_8_port, ZN => n2972);
   U1712 : INV_X1 port map( A => REGISTERS_17_8_port, ZN => n2748);
   U1713 : INV_X1 port map( A => REGISTERS_22_8_port, ZN => n2908);
   U1714 : INV_X1 port map( A => REGISTERS_29_8_port, ZN => n3132);
   U1715 : INV_X1 port map( A => REGISTERS_7_9_port, ZN => n2555);
   U1716 : INV_X1 port map( A => REGISTERS_27_9_port, ZN => n3067);
   U1717 : INV_X1 port map( A => REGISTERS_4_9_port, ZN => n2459);
   U1718 : INV_X1 port map( A => REGISTERS_24_9_port, ZN => n2971);
   U1719 : INV_X1 port map( A => REGISTERS_17_9_port, ZN => n2747);
   U1720 : INV_X1 port map( A => REGISTERS_22_9_port, ZN => n2907);
   U1721 : INV_X1 port map( A => REGISTERS_29_9_port, ZN => n3131);
   U1722 : INV_X1 port map( A => REGISTERS_7_10_port, ZN => n2554);
   U1723 : INV_X1 port map( A => REGISTERS_27_10_port, ZN => n3066);
   U1724 : INV_X1 port map( A => REGISTERS_4_10_port, ZN => n2458);
   U1725 : INV_X1 port map( A => REGISTERS_24_10_port, ZN => n2970);
   U1726 : INV_X1 port map( A => REGISTERS_17_10_port, ZN => n2746);
   U1727 : INV_X1 port map( A => REGISTERS_22_10_port, ZN => n2906);
   U1728 : INV_X1 port map( A => REGISTERS_29_10_port, ZN => n3130);
   U1729 : INV_X1 port map( A => REGISTERS_7_11_port, ZN => n2553);
   U1730 : INV_X1 port map( A => REGISTERS_27_11_port, ZN => n3065);
   U1731 : INV_X1 port map( A => REGISTERS_4_11_port, ZN => n2457);
   U1732 : INV_X1 port map( A => REGISTERS_24_11_port, ZN => n2969);
   U1733 : INV_X1 port map( A => REGISTERS_17_11_port, ZN => n2745);
   U1734 : INV_X1 port map( A => REGISTERS_22_11_port, ZN => n2905);
   U1735 : INV_X1 port map( A => REGISTERS_29_11_port, ZN => n3129);
   U1736 : INV_X1 port map( A => REGISTERS_7_12_port, ZN => n2552);
   U1737 : INV_X1 port map( A => REGISTERS_27_12_port, ZN => n3064);
   U1738 : INV_X1 port map( A => REGISTERS_4_12_port, ZN => n2456);
   U1739 : INV_X1 port map( A => REGISTERS_24_12_port, ZN => n2968);
   U1740 : INV_X1 port map( A => REGISTERS_17_12_port, ZN => n2744);
   U1741 : INV_X1 port map( A => REGISTERS_22_12_port, ZN => n2904);
   U1742 : INV_X1 port map( A => REGISTERS_29_12_port, ZN => n3128);
   U1743 : INV_X1 port map( A => REGISTERS_7_13_port, ZN => n2551);
   U1744 : INV_X1 port map( A => REGISTERS_27_13_port, ZN => n3063);
   U1745 : INV_X1 port map( A => REGISTERS_4_13_port, ZN => n2455);
   U1746 : INV_X1 port map( A => REGISTERS_24_13_port, ZN => n2967);
   U1747 : INV_X1 port map( A => REGISTERS_17_13_port, ZN => n2743);
   U1748 : INV_X1 port map( A => REGISTERS_22_13_port, ZN => n2903);
   U1749 : INV_X1 port map( A => REGISTERS_29_13_port, ZN => n3127);
   U1750 : INV_X1 port map( A => REGISTERS_7_14_port, ZN => n2550);
   U1751 : INV_X1 port map( A => REGISTERS_27_14_port, ZN => n3062);
   U1752 : INV_X1 port map( A => REGISTERS_4_14_port, ZN => n2454);
   U1753 : INV_X1 port map( A => REGISTERS_24_14_port, ZN => n2966);
   U1754 : INV_X1 port map( A => REGISTERS_17_14_port, ZN => n2742);
   U1755 : INV_X1 port map( A => REGISTERS_22_14_port, ZN => n2902);
   U1756 : INV_X1 port map( A => REGISTERS_29_14_port, ZN => n3126);
   U1757 : INV_X1 port map( A => REGISTERS_7_15_port, ZN => n2549);
   U1758 : INV_X1 port map( A => REGISTERS_27_15_port, ZN => n3061);
   U1759 : INV_X1 port map( A => REGISTERS_4_15_port, ZN => n2453);
   U1760 : INV_X1 port map( A => REGISTERS_24_15_port, ZN => n2965);
   U1761 : INV_X1 port map( A => REGISTERS_17_15_port, ZN => n2741);
   U1762 : INV_X1 port map( A => REGISTERS_22_15_port, ZN => n2901);
   U1763 : INV_X1 port map( A => REGISTERS_29_15_port, ZN => n3125);
   U1764 : INV_X1 port map( A => REGISTERS_7_16_port, ZN => n2548);
   U1765 : INV_X1 port map( A => REGISTERS_27_16_port, ZN => n3060);
   U1766 : INV_X1 port map( A => REGISTERS_4_16_port, ZN => n2452);
   U1767 : INV_X1 port map( A => REGISTERS_24_16_port, ZN => n2964);
   U1768 : INV_X1 port map( A => REGISTERS_17_16_port, ZN => n2740);
   U1769 : INV_X1 port map( A => REGISTERS_22_16_port, ZN => n2900);
   U1770 : INV_X1 port map( A => REGISTERS_29_16_port, ZN => n3124);
   U1771 : INV_X1 port map( A => REGISTERS_7_17_port, ZN => n2547);
   U1772 : INV_X1 port map( A => REGISTERS_27_17_port, ZN => n3059);
   U1773 : INV_X1 port map( A => REGISTERS_4_17_port, ZN => n2451);
   U1774 : INV_X1 port map( A => REGISTERS_24_17_port, ZN => n2963);
   U1775 : INV_X1 port map( A => REGISTERS_17_17_port, ZN => n2739);
   U1776 : INV_X1 port map( A => REGISTERS_22_17_port, ZN => n2899);
   U1777 : INV_X1 port map( A => REGISTERS_29_17_port, ZN => n3123);
   U1778 : INV_X1 port map( A => REGISTERS_7_18_port, ZN => n2546);
   U1779 : INV_X1 port map( A => REGISTERS_27_18_port, ZN => n3058);
   U1780 : INV_X1 port map( A => REGISTERS_4_18_port, ZN => n2450);
   U1781 : INV_X1 port map( A => REGISTERS_24_18_port, ZN => n2962);
   U1782 : INV_X1 port map( A => REGISTERS_17_18_port, ZN => n2738);
   U1783 : INV_X1 port map( A => REGISTERS_22_18_port, ZN => n2898);
   U1784 : INV_X1 port map( A => REGISTERS_29_18_port, ZN => n3122);
   U1785 : INV_X1 port map( A => REGISTERS_7_19_port, ZN => n2545);
   U1786 : INV_X1 port map( A => REGISTERS_27_19_port, ZN => n3057);
   U1787 : INV_X1 port map( A => REGISTERS_4_19_port, ZN => n2449);
   U1788 : INV_X1 port map( A => REGISTERS_24_19_port, ZN => n2961);
   U1789 : INV_X1 port map( A => REGISTERS_17_19_port, ZN => n2737);
   U1790 : INV_X1 port map( A => REGISTERS_22_19_port, ZN => n2897);
   U1791 : INV_X1 port map( A => REGISTERS_29_19_port, ZN => n3121);
   U1792 : INV_X1 port map( A => REGISTERS_7_20_port, ZN => n2544);
   U1793 : INV_X1 port map( A => REGISTERS_27_20_port, ZN => n3056);
   U1794 : INV_X1 port map( A => REGISTERS_4_20_port, ZN => n2448);
   U1795 : INV_X1 port map( A => REGISTERS_24_20_port, ZN => n2960);
   U1796 : INV_X1 port map( A => REGISTERS_17_20_port, ZN => n2736);
   U1797 : INV_X1 port map( A => REGISTERS_22_20_port, ZN => n2896);
   U1798 : INV_X1 port map( A => REGISTERS_29_20_port, ZN => n3120);
   U1799 : INV_X1 port map( A => REGISTERS_7_21_port, ZN => n2543);
   U1800 : INV_X1 port map( A => REGISTERS_27_21_port, ZN => n3055);
   U1801 : INV_X1 port map( A => REGISTERS_4_21_port, ZN => n2447);
   U1802 : INV_X1 port map( A => REGISTERS_24_21_port, ZN => n2959);
   U1803 : INV_X1 port map( A => REGISTERS_17_21_port, ZN => n2735);
   U1804 : INV_X1 port map( A => REGISTERS_22_21_port, ZN => n2895);
   U1805 : INV_X1 port map( A => REGISTERS_29_21_port, ZN => n3119);
   U1806 : INV_X1 port map( A => REGISTERS_7_22_port, ZN => n2542);
   U1807 : INV_X1 port map( A => REGISTERS_27_22_port, ZN => n3054);
   U1808 : INV_X1 port map( A => REGISTERS_4_22_port, ZN => n2446);
   U1809 : INV_X1 port map( A => REGISTERS_24_22_port, ZN => n2958);
   U1810 : INV_X1 port map( A => REGISTERS_17_22_port, ZN => n2734);
   U1811 : INV_X1 port map( A => REGISTERS_22_22_port, ZN => n2894);
   U1812 : INV_X1 port map( A => REGISTERS_29_22_port, ZN => n3118);
   U1813 : INV_X1 port map( A => REGISTERS_7_23_port, ZN => n2541);
   U1814 : INV_X1 port map( A => REGISTERS_27_23_port, ZN => n3053);
   U1815 : INV_X1 port map( A => REGISTERS_4_23_port, ZN => n2445);
   U1816 : INV_X1 port map( A => REGISTERS_24_23_port, ZN => n2957);
   U1817 : INV_X1 port map( A => REGISTERS_17_23_port, ZN => n2733);
   U1818 : INV_X1 port map( A => REGISTERS_22_23_port, ZN => n2893);
   U1819 : INV_X1 port map( A => REGISTERS_29_23_port, ZN => n3117);
   U1820 : INV_X1 port map( A => REGISTERS_7_24_port, ZN => n2540);
   U1821 : INV_X1 port map( A => REGISTERS_27_24_port, ZN => n3052);
   U1822 : INV_X1 port map( A => REGISTERS_4_24_port, ZN => n2444);
   U1823 : INV_X1 port map( A => REGISTERS_24_24_port, ZN => n2956);
   U1824 : INV_X1 port map( A => REGISTERS_17_24_port, ZN => n2732);
   U1825 : INV_X1 port map( A => REGISTERS_22_24_port, ZN => n2892);
   U1826 : INV_X1 port map( A => REGISTERS_29_24_port, ZN => n3116);
   U1827 : INV_X1 port map( A => REGISTERS_7_25_port, ZN => n2539);
   U1828 : INV_X1 port map( A => REGISTERS_27_25_port, ZN => n3051);
   U1829 : INV_X1 port map( A => REGISTERS_4_25_port, ZN => n2443);
   U1830 : INV_X1 port map( A => REGISTERS_24_25_port, ZN => n2955);
   U1831 : INV_X1 port map( A => REGISTERS_17_25_port, ZN => n2731);
   U1832 : INV_X1 port map( A => REGISTERS_22_25_port, ZN => n2891);
   U1833 : INV_X1 port map( A => REGISTERS_29_25_port, ZN => n3115);
   U1834 : INV_X1 port map( A => REGISTERS_7_26_port, ZN => n2538);
   U1835 : INV_X1 port map( A => REGISTERS_27_26_port, ZN => n3050);
   U1836 : INV_X1 port map( A => REGISTERS_4_26_port, ZN => n2442);
   U1837 : INV_X1 port map( A => REGISTERS_24_26_port, ZN => n2954);
   U1838 : INV_X1 port map( A => REGISTERS_17_26_port, ZN => n2730);
   U1839 : INV_X1 port map( A => REGISTERS_22_26_port, ZN => n2890);
   U1840 : INV_X1 port map( A => REGISTERS_29_26_port, ZN => n3114);
   U1841 : INV_X1 port map( A => REGISTERS_7_27_port, ZN => n2537);
   U1842 : INV_X1 port map( A => REGISTERS_27_27_port, ZN => n3049);
   U1843 : INV_X1 port map( A => REGISTERS_4_27_port, ZN => n2441);
   U1844 : INV_X1 port map( A => REGISTERS_24_27_port, ZN => n2953);
   U1845 : INV_X1 port map( A => REGISTERS_17_27_port, ZN => n2729);
   U1846 : INV_X1 port map( A => REGISTERS_22_27_port, ZN => n2889);
   U1847 : INV_X1 port map( A => REGISTERS_29_27_port, ZN => n3113);
   U1848 : INV_X1 port map( A => REGISTERS_7_28_port, ZN => n2536);
   U1849 : INV_X1 port map( A => REGISTERS_27_28_port, ZN => n3048);
   U1850 : INV_X1 port map( A => REGISTERS_4_28_port, ZN => n2440);
   U1851 : INV_X1 port map( A => REGISTERS_24_28_port, ZN => n2952);
   U1852 : INV_X1 port map( A => REGISTERS_17_28_port, ZN => n2728);
   U1853 : INV_X1 port map( A => REGISTERS_22_28_port, ZN => n2888);
   U1854 : INV_X1 port map( A => REGISTERS_29_28_port, ZN => n3112);
   U1855 : INV_X1 port map( A => REGISTERS_7_29_port, ZN => n2535);
   U1856 : INV_X1 port map( A => REGISTERS_27_29_port, ZN => n3047);
   U1857 : INV_X1 port map( A => REGISTERS_4_29_port, ZN => n2439);
   U1858 : INV_X1 port map( A => REGISTERS_24_29_port, ZN => n2951);
   U1859 : INV_X1 port map( A => REGISTERS_17_29_port, ZN => n2727);
   U1860 : INV_X1 port map( A => REGISTERS_22_29_port, ZN => n2887);
   U1861 : INV_X1 port map( A => REGISTERS_29_29_port, ZN => n3111);
   U1862 : INV_X1 port map( A => REGISTERS_7_30_port, ZN => n2534);
   U1863 : INV_X1 port map( A => REGISTERS_27_30_port, ZN => n3046);
   U1864 : INV_X1 port map( A => REGISTERS_4_30_port, ZN => n2438);
   U1865 : INV_X1 port map( A => REGISTERS_24_30_port, ZN => n2950);
   U1866 : INV_X1 port map( A => REGISTERS_17_30_port, ZN => n2726);
   U1867 : INV_X1 port map( A => REGISTERS_22_30_port, ZN => n2886);
   U1868 : INV_X1 port map( A => REGISTERS_29_30_port, ZN => n3110);
   U1869 : INV_X1 port map( A => REGISTERS_7_31_port, ZN => n2533);
   U1870 : INV_X1 port map( A => REGISTERS_27_31_port, ZN => n3045);
   U1871 : INV_X1 port map( A => REGISTERS_4_31_port, ZN => n2437);
   U1872 : INV_X1 port map( A => REGISTERS_24_31_port, ZN => n2949);
   U1873 : INV_X1 port map( A => REGISTERS_17_31_port, ZN => n2725);
   U1874 : INV_X1 port map( A => REGISTERS_22_31_port, ZN => n2885);
   U1875 : INV_X1 port map( A => REGISTERS_29_31_port, ZN => n3109);
   U1876 : INV_X1 port map( A => REGISTERS_1_0_port, ZN => n2372);
   U1877 : INV_X1 port map( A => REGISTERS_28_0_port, ZN => n3108);
   U1878 : INV_X1 port map( A => REGISTERS_6_0_port, ZN => n2532);
   U1879 : INV_X1 port map( A => REGISTERS_2_0_port, ZN => n2404);
   U1880 : INV_X1 port map( A => REGISTERS_20_0_port, ZN => n2852);
   U1881 : INV_X1 port map( A => REGISTERS_18_0_port, ZN => n2788);
   U1882 : INV_X1 port map( A => REGISTERS_31_0_port, ZN => n3204);
   U1883 : INV_X1 port map( A => REGISTERS_1_1_port, ZN => n2371);
   U1884 : INV_X1 port map( A => REGISTERS_28_1_port, ZN => n3107);
   U1885 : INV_X1 port map( A => REGISTERS_6_1_port, ZN => n2531);
   U1886 : INV_X1 port map( A => REGISTERS_2_1_port, ZN => n2403);
   U1887 : INV_X1 port map( A => REGISTERS_20_1_port, ZN => n2851);
   U1888 : INV_X1 port map( A => REGISTERS_18_1_port, ZN => n2787);
   U1889 : INV_X1 port map( A => REGISTERS_31_1_port, ZN => n3203);
   U1890 : INV_X1 port map( A => REGISTERS_1_2_port, ZN => n2370);
   U1891 : INV_X1 port map( A => REGISTERS_28_2_port, ZN => n3106);
   U1892 : INV_X1 port map( A => REGISTERS_6_2_port, ZN => n2530);
   U1893 : INV_X1 port map( A => REGISTERS_2_2_port, ZN => n2402);
   U1894 : INV_X1 port map( A => REGISTERS_20_2_port, ZN => n2850);
   U1895 : INV_X1 port map( A => REGISTERS_18_2_port, ZN => n2786);
   U1896 : INV_X1 port map( A => REGISTERS_31_2_port, ZN => n3202);
   U1897 : INV_X1 port map( A => REGISTERS_1_3_port, ZN => n2369);
   U1898 : INV_X1 port map( A => REGISTERS_28_3_port, ZN => n3105);
   U1899 : INV_X1 port map( A => REGISTERS_6_3_port, ZN => n2529);
   U1900 : INV_X1 port map( A => REGISTERS_2_3_port, ZN => n2401);
   U1901 : INV_X1 port map( A => REGISTERS_20_3_port, ZN => n2849);
   U1902 : INV_X1 port map( A => REGISTERS_18_3_port, ZN => n2785);
   U1903 : INV_X1 port map( A => REGISTERS_31_3_port, ZN => n3201);
   U1904 : INV_X1 port map( A => REGISTERS_1_4_port, ZN => n2368);
   U1905 : INV_X1 port map( A => REGISTERS_28_4_port, ZN => n3104);
   U1906 : INV_X1 port map( A => REGISTERS_6_4_port, ZN => n2528);
   U1907 : INV_X1 port map( A => REGISTERS_2_4_port, ZN => n2400);
   U1908 : INV_X1 port map( A => REGISTERS_20_4_port, ZN => n2848);
   U1909 : INV_X1 port map( A => REGISTERS_18_4_port, ZN => n2784);
   U1910 : INV_X1 port map( A => REGISTERS_31_4_port, ZN => n3200);
   U1911 : INV_X1 port map( A => REGISTERS_1_5_port, ZN => n2367);
   U1912 : INV_X1 port map( A => REGISTERS_28_5_port, ZN => n3103);
   U1913 : INV_X1 port map( A => REGISTERS_6_5_port, ZN => n2527);
   U1914 : INV_X1 port map( A => REGISTERS_2_5_port, ZN => n2399);
   U1915 : INV_X1 port map( A => REGISTERS_20_5_port, ZN => n2847);
   U1916 : INV_X1 port map( A => REGISTERS_18_5_port, ZN => n2783);
   U1917 : INV_X1 port map( A => REGISTERS_31_5_port, ZN => n3199);
   U1918 : INV_X1 port map( A => REGISTERS_1_6_port, ZN => n2366);
   U1919 : INV_X1 port map( A => REGISTERS_28_6_port, ZN => n3102);
   U1920 : INV_X1 port map( A => REGISTERS_6_6_port, ZN => n2526);
   U1921 : INV_X1 port map( A => REGISTERS_2_6_port, ZN => n2398);
   U1922 : INV_X1 port map( A => REGISTERS_20_6_port, ZN => n2846);
   U1923 : INV_X1 port map( A => REGISTERS_18_6_port, ZN => n2782);
   U1924 : INV_X1 port map( A => REGISTERS_31_6_port, ZN => n3198);
   U1925 : INV_X1 port map( A => REGISTERS_1_7_port, ZN => n2365);
   U1926 : INV_X1 port map( A => REGISTERS_28_7_port, ZN => n3101);
   U1927 : INV_X1 port map( A => REGISTERS_6_7_port, ZN => n2525);
   U1928 : INV_X1 port map( A => REGISTERS_2_7_port, ZN => n2397);
   U1929 : INV_X1 port map( A => REGISTERS_20_7_port, ZN => n2845);
   U1930 : INV_X1 port map( A => REGISTERS_18_7_port, ZN => n2781);
   U1931 : INV_X1 port map( A => REGISTERS_31_7_port, ZN => n3197);
   U1932 : INV_X1 port map( A => REGISTERS_1_8_port, ZN => n2364);
   U1933 : INV_X1 port map( A => REGISTERS_28_8_port, ZN => n3100);
   U1934 : INV_X1 port map( A => REGISTERS_6_8_port, ZN => n2524);
   U1935 : INV_X1 port map( A => REGISTERS_2_8_port, ZN => n2396);
   U1936 : INV_X1 port map( A => REGISTERS_20_8_port, ZN => n2844);
   U1937 : INV_X1 port map( A => REGISTERS_18_8_port, ZN => n2780);
   U1938 : INV_X1 port map( A => REGISTERS_31_8_port, ZN => n3196);
   U1939 : INV_X1 port map( A => REGISTERS_1_9_port, ZN => n2363);
   U1940 : INV_X1 port map( A => REGISTERS_28_9_port, ZN => n3099);
   U1941 : INV_X1 port map( A => REGISTERS_6_9_port, ZN => n2523);
   U1942 : INV_X1 port map( A => REGISTERS_2_9_port, ZN => n2395);
   U1943 : INV_X1 port map( A => REGISTERS_20_9_port, ZN => n2843);
   U1944 : INV_X1 port map( A => REGISTERS_18_9_port, ZN => n2779);
   U1945 : INV_X1 port map( A => REGISTERS_31_9_port, ZN => n3195);
   U1946 : INV_X1 port map( A => REGISTERS_1_10_port, ZN => n2362);
   U1947 : INV_X1 port map( A => REGISTERS_28_10_port, ZN => n3098);
   U1948 : INV_X1 port map( A => REGISTERS_6_10_port, ZN => n2522);
   U1949 : INV_X1 port map( A => REGISTERS_2_10_port, ZN => n2394);
   U1950 : INV_X1 port map( A => REGISTERS_20_10_port, ZN => n2842);
   U1951 : INV_X1 port map( A => REGISTERS_18_10_port, ZN => n2778);
   U1952 : INV_X1 port map( A => REGISTERS_31_10_port, ZN => n3194);
   U1953 : INV_X1 port map( A => REGISTERS_1_11_port, ZN => n2361);
   U1954 : INV_X1 port map( A => REGISTERS_28_11_port, ZN => n3097);
   U1955 : INV_X1 port map( A => REGISTERS_6_11_port, ZN => n2521);
   U1956 : INV_X1 port map( A => REGISTERS_2_11_port, ZN => n2393);
   U1957 : INV_X1 port map( A => REGISTERS_20_11_port, ZN => n2841);
   U1958 : INV_X1 port map( A => REGISTERS_18_11_port, ZN => n2777);
   U1959 : INV_X1 port map( A => REGISTERS_31_11_port, ZN => n3193);
   U1960 : INV_X1 port map( A => REGISTERS_1_12_port, ZN => n2360);
   U1961 : INV_X1 port map( A => REGISTERS_28_12_port, ZN => n3096);
   U1962 : INV_X1 port map( A => REGISTERS_6_12_port, ZN => n2520);
   U1963 : INV_X1 port map( A => REGISTERS_2_12_port, ZN => n2392);
   U1964 : INV_X1 port map( A => REGISTERS_20_12_port, ZN => n2840);
   U1965 : INV_X1 port map( A => REGISTERS_18_12_port, ZN => n2776);
   U1966 : INV_X1 port map( A => REGISTERS_31_12_port, ZN => n3192);
   U1967 : INV_X1 port map( A => REGISTERS_1_13_port, ZN => n2359);
   U1968 : INV_X1 port map( A => REGISTERS_28_13_port, ZN => n3095);
   U1969 : INV_X1 port map( A => REGISTERS_6_13_port, ZN => n2519);
   U1970 : INV_X1 port map( A => REGISTERS_2_13_port, ZN => n2391);
   U1971 : INV_X1 port map( A => REGISTERS_20_13_port, ZN => n2839);
   U1972 : INV_X1 port map( A => REGISTERS_18_13_port, ZN => n2775);
   U1973 : INV_X1 port map( A => REGISTERS_31_13_port, ZN => n3191);
   U1974 : INV_X1 port map( A => REGISTERS_1_14_port, ZN => n2358);
   U1975 : INV_X1 port map( A => REGISTERS_28_14_port, ZN => n3094);
   U1976 : INV_X1 port map( A => REGISTERS_6_14_port, ZN => n2518);
   U1977 : INV_X1 port map( A => REGISTERS_2_14_port, ZN => n2390);
   U1978 : INV_X1 port map( A => REGISTERS_20_14_port, ZN => n2838);
   U1979 : INV_X1 port map( A => REGISTERS_18_14_port, ZN => n2774);
   U1980 : INV_X1 port map( A => REGISTERS_31_14_port, ZN => n3190);
   U1981 : INV_X1 port map( A => REGISTERS_1_15_port, ZN => n2357);
   U1982 : INV_X1 port map( A => REGISTERS_28_15_port, ZN => n3093);
   U1983 : INV_X1 port map( A => REGISTERS_6_15_port, ZN => n2517);
   U1984 : INV_X1 port map( A => REGISTERS_2_15_port, ZN => n2389);
   U1985 : INV_X1 port map( A => REGISTERS_20_15_port, ZN => n2837);
   U1986 : INV_X1 port map( A => REGISTERS_18_15_port, ZN => n2773);
   U1987 : INV_X1 port map( A => REGISTERS_31_15_port, ZN => n3189);
   U1988 : INV_X1 port map( A => REGISTERS_1_16_port, ZN => n2356);
   U1989 : INV_X1 port map( A => REGISTERS_28_16_port, ZN => n3092);
   U1990 : INV_X1 port map( A => REGISTERS_6_16_port, ZN => n2516);
   U1991 : INV_X1 port map( A => REGISTERS_2_16_port, ZN => n2388);
   U1992 : INV_X1 port map( A => REGISTERS_20_16_port, ZN => n2836);
   U1993 : INV_X1 port map( A => REGISTERS_18_16_port, ZN => n2772);
   U1994 : INV_X1 port map( A => REGISTERS_31_16_port, ZN => n3188);
   U1995 : INV_X1 port map( A => REGISTERS_1_17_port, ZN => n2355);
   U1996 : INV_X1 port map( A => REGISTERS_28_17_port, ZN => n3091);
   U1997 : INV_X1 port map( A => REGISTERS_6_17_port, ZN => n2515);
   U1998 : INV_X1 port map( A => REGISTERS_2_17_port, ZN => n2387);
   U1999 : INV_X1 port map( A => REGISTERS_20_17_port, ZN => n2835);
   U2000 : INV_X1 port map( A => REGISTERS_18_17_port, ZN => n2771);
   U2001 : INV_X1 port map( A => REGISTERS_31_17_port, ZN => n3187);
   U2002 : INV_X1 port map( A => REGISTERS_1_18_port, ZN => n2354);
   U2003 : INV_X1 port map( A => REGISTERS_28_18_port, ZN => n3090);
   U2004 : INV_X1 port map( A => REGISTERS_6_18_port, ZN => n2514);
   U2005 : INV_X1 port map( A => REGISTERS_2_18_port, ZN => n2386);
   U2006 : INV_X1 port map( A => REGISTERS_20_18_port, ZN => n2834);
   U2007 : INV_X1 port map( A => REGISTERS_18_18_port, ZN => n2770);
   U2008 : INV_X1 port map( A => REGISTERS_31_18_port, ZN => n3186);
   U2009 : INV_X1 port map( A => REGISTERS_1_19_port, ZN => n2353);
   U2010 : INV_X1 port map( A => REGISTERS_28_19_port, ZN => n3089);
   U2011 : INV_X1 port map( A => REGISTERS_6_19_port, ZN => n2513);
   U2012 : INV_X1 port map( A => REGISTERS_2_19_port, ZN => n2385);
   U2013 : INV_X1 port map( A => REGISTERS_20_19_port, ZN => n2833);
   U2014 : INV_X1 port map( A => REGISTERS_18_19_port, ZN => n2769);
   U2015 : INV_X1 port map( A => REGISTERS_31_19_port, ZN => n3185);
   U2016 : INV_X1 port map( A => REGISTERS_1_20_port, ZN => n2352);
   U2017 : INV_X1 port map( A => REGISTERS_28_20_port, ZN => n3088);
   U2018 : INV_X1 port map( A => REGISTERS_6_20_port, ZN => n2512);
   U2019 : INV_X1 port map( A => REGISTERS_2_20_port, ZN => n2384);
   U2020 : INV_X1 port map( A => REGISTERS_20_20_port, ZN => n2832);
   U2021 : INV_X1 port map( A => REGISTERS_18_20_port, ZN => n2768);
   U2022 : INV_X1 port map( A => REGISTERS_31_20_port, ZN => n3184);
   U2023 : INV_X1 port map( A => REGISTERS_1_21_port, ZN => n2351);
   U2024 : INV_X1 port map( A => REGISTERS_28_21_port, ZN => n3087);
   U2025 : INV_X1 port map( A => REGISTERS_6_21_port, ZN => n2511);
   U2026 : INV_X1 port map( A => REGISTERS_2_21_port, ZN => n2383);
   U2027 : INV_X1 port map( A => REGISTERS_20_21_port, ZN => n2831);
   U2028 : INV_X1 port map( A => REGISTERS_18_21_port, ZN => n2767);
   U2029 : INV_X1 port map( A => REGISTERS_31_21_port, ZN => n3183);
   U2030 : INV_X1 port map( A => REGISTERS_1_22_port, ZN => n2350);
   U2031 : INV_X1 port map( A => REGISTERS_28_22_port, ZN => n3086);
   U2032 : INV_X1 port map( A => REGISTERS_6_22_port, ZN => n2510);
   U2033 : INV_X1 port map( A => REGISTERS_2_22_port, ZN => n2382);
   U2034 : INV_X1 port map( A => REGISTERS_20_22_port, ZN => n2830);
   U2035 : INV_X1 port map( A => REGISTERS_18_22_port, ZN => n2766);
   U2036 : INV_X1 port map( A => REGISTERS_31_22_port, ZN => n3182);
   U2037 : INV_X1 port map( A => REGISTERS_1_23_port, ZN => n2349);
   U2038 : INV_X1 port map( A => REGISTERS_28_23_port, ZN => n3085);
   U2039 : INV_X1 port map( A => REGISTERS_6_23_port, ZN => n2509);
   U2040 : INV_X1 port map( A => REGISTERS_2_23_port, ZN => n2381);
   U2041 : INV_X1 port map( A => REGISTERS_20_23_port, ZN => n2829);
   U2042 : INV_X1 port map( A => REGISTERS_18_23_port, ZN => n2765);
   U2055 : INV_X1 port map( A => REGISTERS_31_23_port, ZN => n3181);
   U2056 : INV_X1 port map( A => REGISTERS_1_24_port, ZN => n2348);
   U2057 : INV_X1 port map( A => REGISTERS_28_24_port, ZN => n3084);
   U2058 : INV_X1 port map( A => REGISTERS_6_24_port, ZN => n2508);
   U2059 : INV_X1 port map( A => REGISTERS_2_24_port, ZN => n2380);
   U2060 : INV_X1 port map( A => REGISTERS_20_24_port, ZN => n2828);
   U2061 : INV_X1 port map( A => REGISTERS_18_24_port, ZN => n2764);
   U2062 : INV_X1 port map( A => REGISTERS_31_24_port, ZN => n3180);
   U2063 : INV_X1 port map( A => REGISTERS_1_25_port, ZN => n2347);
   U2064 : INV_X1 port map( A => REGISTERS_28_25_port, ZN => n3083);
   U2065 : INV_X1 port map( A => REGISTERS_6_25_port, ZN => n2507);
   U2066 : INV_X1 port map( A => REGISTERS_2_25_port, ZN => n2379);
   U2067 : INV_X1 port map( A => REGISTERS_20_25_port, ZN => n2827);
   U2068 : INV_X1 port map( A => REGISTERS_18_25_port, ZN => n2763);
   U2069 : INV_X1 port map( A => REGISTERS_31_25_port, ZN => n3179);
   U2070 : INV_X1 port map( A => REGISTERS_1_26_port, ZN => n2346);
   U2071 : INV_X1 port map( A => REGISTERS_28_26_port, ZN => n3082);
   U2072 : INV_X1 port map( A => REGISTERS_6_26_port, ZN => n2506);
   U2073 : INV_X1 port map( A => REGISTERS_2_26_port, ZN => n2378);
   U2074 : INV_X1 port map( A => REGISTERS_20_26_port, ZN => n2826);
   U2075 : INV_X1 port map( A => REGISTERS_18_26_port, ZN => n2762);
   U2076 : INV_X1 port map( A => REGISTERS_31_26_port, ZN => n3178);
   U2077 : INV_X1 port map( A => REGISTERS_1_27_port, ZN => n2345);
   U2078 : INV_X1 port map( A => REGISTERS_28_27_port, ZN => n3081);
   U2079 : INV_X1 port map( A => REGISTERS_6_27_port, ZN => n2505);
   U2080 : INV_X1 port map( A => REGISTERS_2_27_port, ZN => n2377);
   U2081 : INV_X1 port map( A => REGISTERS_20_27_port, ZN => n2825);
   U2082 : INV_X1 port map( A => REGISTERS_18_27_port, ZN => n2761);
   U2083 : INV_X1 port map( A => REGISTERS_31_27_port, ZN => n3177);
   U2084 : INV_X1 port map( A => REGISTERS_1_28_port, ZN => n2344);
   U2085 : INV_X1 port map( A => REGISTERS_28_28_port, ZN => n3080);
   U2086 : INV_X1 port map( A => REGISTERS_6_28_port, ZN => n2504);
   U2087 : INV_X1 port map( A => REGISTERS_2_28_port, ZN => n2376);
   U2088 : INV_X1 port map( A => REGISTERS_20_28_port, ZN => n2824);
   U2089 : INV_X1 port map( A => REGISTERS_18_28_port, ZN => n2760);
   U2090 : INV_X1 port map( A => REGISTERS_31_28_port, ZN => n3176);
   U2091 : INV_X1 port map( A => REGISTERS_1_29_port, ZN => n2343);
   U2092 : INV_X1 port map( A => REGISTERS_28_29_port, ZN => n3079);
   U2093 : INV_X1 port map( A => REGISTERS_6_29_port, ZN => n2503);
   U2094 : INV_X1 port map( A => REGISTERS_2_29_port, ZN => n2375);
   U2095 : INV_X1 port map( A => REGISTERS_20_29_port, ZN => n2823);
   U2096 : INV_X1 port map( A => REGISTERS_18_29_port, ZN => n2759);
   U2097 : INV_X1 port map( A => REGISTERS_31_29_port, ZN => n3175);
   U2098 : INV_X1 port map( A => REGISTERS_1_30_port, ZN => n2342);
   U2099 : INV_X1 port map( A => REGISTERS_28_30_port, ZN => n3078);
   U2100 : INV_X1 port map( A => REGISTERS_6_30_port, ZN => n2502);
   U2101 : INV_X1 port map( A => REGISTERS_2_30_port, ZN => n2374);
   U2102 : INV_X1 port map( A => REGISTERS_20_30_port, ZN => n2822);
   U2103 : INV_X1 port map( A => REGISTERS_18_30_port, ZN => n2758);
   U2104 : INV_X1 port map( A => REGISTERS_31_30_port, ZN => n3174);
   U2105 : INV_X1 port map( A => REGISTERS_1_31_port, ZN => n2341);
   U2106 : INV_X1 port map( A => REGISTERS_28_31_port, ZN => n3077);
   U2107 : INV_X1 port map( A => REGISTERS_6_31_port, ZN => n2501);
   U2108 : INV_X1 port map( A => REGISTERS_2_31_port, ZN => n2373);
   U2109 : INV_X1 port map( A => REGISTERS_20_31_port, ZN => n2821);
   U2110 : INV_X1 port map( A => REGISTERS_18_31_port, ZN => n2757);
   U2111 : INV_X1 port map( A => REGISTERS_31_31_port, ZN => n3173);
   U2112 : INV_X1 port map( A => REGISTERS_13_0_port, ZN => n2628);
   U2113 : INV_X1 port map( A => REGISTERS_12_0_port, ZN => n2596);
   U2114 : INV_X1 port map( A => REGISTERS_13_1_port, ZN => n2627);
   U2115 : INV_X1 port map( A => REGISTERS_12_1_port, ZN => n2595);
   U2116 : INV_X1 port map( A => REGISTERS_13_2_port, ZN => n2626);
   U2117 : INV_X1 port map( A => REGISTERS_12_2_port, ZN => n2594);
   U2118 : INV_X1 port map( A => REGISTERS_13_3_port, ZN => n2625);
   U2119 : INV_X1 port map( A => REGISTERS_12_3_port, ZN => n2593);
   U2120 : INV_X1 port map( A => REGISTERS_13_4_port, ZN => n2624);
   U2121 : INV_X1 port map( A => REGISTERS_12_4_port, ZN => n2592);
   U2122 : INV_X1 port map( A => REGISTERS_13_5_port, ZN => n2623);
   U2123 : INV_X1 port map( A => REGISTERS_12_5_port, ZN => n2591);
   U2124 : INV_X1 port map( A => REGISTERS_13_6_port, ZN => n2622);
   U2125 : INV_X1 port map( A => REGISTERS_12_6_port, ZN => n2590);
   U2126 : INV_X1 port map( A => REGISTERS_13_7_port, ZN => n2621);
   U2127 : INV_X1 port map( A => REGISTERS_12_7_port, ZN => n2589);
   U2128 : INV_X1 port map( A => REGISTERS_13_8_port, ZN => n2620);
   U2129 : INV_X1 port map( A => REGISTERS_12_8_port, ZN => n2588);
   U2130 : INV_X1 port map( A => REGISTERS_13_9_port, ZN => n2619);
   U2131 : INV_X1 port map( A => REGISTERS_12_9_port, ZN => n2587);
   U2132 : INV_X1 port map( A => REGISTERS_13_10_port, ZN => n2618);
   U2133 : INV_X1 port map( A => REGISTERS_12_10_port, ZN => n2586);
   U2134 : INV_X1 port map( A => REGISTERS_13_11_port, ZN => n2617);
   U2135 : INV_X1 port map( A => REGISTERS_12_11_port, ZN => n2585);
   U2136 : INV_X1 port map( A => REGISTERS_13_12_port, ZN => n2616);
   U2137 : INV_X1 port map( A => REGISTERS_12_12_port, ZN => n2584);
   U2138 : INV_X1 port map( A => REGISTERS_13_13_port, ZN => n2615);
   U2139 : INV_X1 port map( A => REGISTERS_12_13_port, ZN => n2583);
   U2140 : INV_X1 port map( A => REGISTERS_13_14_port, ZN => n2614);
   U2141 : INV_X1 port map( A => REGISTERS_12_14_port, ZN => n2582);
   U2142 : INV_X1 port map( A => REGISTERS_13_15_port, ZN => n2613);
   U2143 : INV_X1 port map( A => REGISTERS_12_15_port, ZN => n2581);
   U2144 : INV_X1 port map( A => REGISTERS_13_16_port, ZN => n2612);
   U2145 : INV_X1 port map( A => REGISTERS_12_16_port, ZN => n2580);
   U2146 : INV_X1 port map( A => REGISTERS_13_17_port, ZN => n2611);
   U2147 : INV_X1 port map( A => REGISTERS_12_17_port, ZN => n2579);
   U2148 : INV_X1 port map( A => REGISTERS_13_18_port, ZN => n2610);
   U2149 : INV_X1 port map( A => REGISTERS_12_18_port, ZN => n2578);
   U2150 : INV_X1 port map( A => REGISTERS_13_19_port, ZN => n2609);
   U2151 : INV_X1 port map( A => REGISTERS_12_19_port, ZN => n2577);
   U2152 : INV_X1 port map( A => REGISTERS_13_20_port, ZN => n2608);
   U2153 : INV_X1 port map( A => REGISTERS_12_20_port, ZN => n2576);
   U2154 : INV_X1 port map( A => REGISTERS_13_21_port, ZN => n2607);
   U2155 : INV_X1 port map( A => REGISTERS_12_21_port, ZN => n2575);
   U2156 : INV_X1 port map( A => REGISTERS_13_22_port, ZN => n2606);
   U2157 : INV_X1 port map( A => REGISTERS_12_22_port, ZN => n2574);
   U2158 : INV_X1 port map( A => REGISTERS_13_23_port, ZN => n2605);
   U2159 : INV_X1 port map( A => REGISTERS_12_23_port, ZN => n2573);
   U2160 : INV_X1 port map( A => REGISTERS_13_24_port, ZN => n2604);
   U2161 : INV_X1 port map( A => REGISTERS_12_24_port, ZN => n2572);
   U2162 : INV_X1 port map( A => REGISTERS_13_25_port, ZN => n2603);
   U2163 : INV_X1 port map( A => REGISTERS_12_25_port, ZN => n2571);
   U2164 : INV_X1 port map( A => REGISTERS_13_26_port, ZN => n2602);
   U2165 : INV_X1 port map( A => REGISTERS_12_26_port, ZN => n2570);
   U2166 : INV_X1 port map( A => REGISTERS_13_27_port, ZN => n2601);
   U2167 : INV_X1 port map( A => REGISTERS_12_27_port, ZN => n2569);
   U2168 : INV_X1 port map( A => REGISTERS_13_28_port, ZN => n2600);
   U2169 : INV_X1 port map( A => REGISTERS_12_28_port, ZN => n2568);
   U2170 : INV_X1 port map( A => REGISTERS_13_29_port, ZN => n2599);
   U2171 : INV_X1 port map( A => REGISTERS_12_29_port, ZN => n2567);
   U2172 : INV_X1 port map( A => REGISTERS_13_30_port, ZN => n2598);
   U2173 : INV_X1 port map( A => REGISTERS_12_30_port, ZN => n2566);
   U2174 : INV_X1 port map( A => REGISTERS_13_31_port, ZN => n2597);
   U2175 : INV_X1 port map( A => REGISTERS_12_31_port, ZN => n2565);
   U2176 : INV_X1 port map( A => REGISTERS_21_0_port, ZN => n2884);
   U2177 : INV_X1 port map( A => REGISTERS_21_1_port, ZN => n2883);
   U2178 : INV_X1 port map( A => REGISTERS_21_2_port, ZN => n2882);
   U2179 : INV_X1 port map( A => REGISTERS_21_3_port, ZN => n2881);
   U2180 : INV_X1 port map( A => REGISTERS_21_4_port, ZN => n2880);
   U2181 : INV_X1 port map( A => REGISTERS_21_5_port, ZN => n2879);
   U2182 : INV_X1 port map( A => REGISTERS_21_6_port, ZN => n2878);
   U2183 : INV_X1 port map( A => REGISTERS_21_7_port, ZN => n2877);
   U2184 : INV_X1 port map( A => REGISTERS_21_8_port, ZN => n2876);
   U2185 : INV_X1 port map( A => REGISTERS_21_9_port, ZN => n2875);
   U2186 : INV_X1 port map( A => REGISTERS_21_10_port, ZN => n2874);
   U2187 : INV_X1 port map( A => REGISTERS_21_11_port, ZN => n2873);
   U2188 : INV_X1 port map( A => REGISTERS_21_12_port, ZN => n2872);
   U2189 : INV_X1 port map( A => REGISTERS_21_13_port, ZN => n2871);
   U2190 : INV_X1 port map( A => REGISTERS_21_14_port, ZN => n2870);
   U2191 : INV_X1 port map( A => REGISTERS_21_15_port, ZN => n2869);
   U2192 : INV_X1 port map( A => REGISTERS_21_16_port, ZN => n2868);
   U2193 : INV_X1 port map( A => REGISTERS_21_17_port, ZN => n2867);
   U2194 : INV_X1 port map( A => REGISTERS_21_18_port, ZN => n2866);
   U2195 : INV_X1 port map( A => REGISTERS_21_19_port, ZN => n2865);
   U2196 : INV_X1 port map( A => REGISTERS_21_20_port, ZN => n2864);
   U2197 : INV_X1 port map( A => REGISTERS_21_21_port, ZN => n2863);
   U2198 : INV_X1 port map( A => REGISTERS_21_22_port, ZN => n2862);
   U2199 : INV_X1 port map( A => REGISTERS_21_23_port, ZN => n2861);
   U2200 : INV_X1 port map( A => REGISTERS_21_24_port, ZN => n2860);
   U2201 : INV_X1 port map( A => REGISTERS_21_25_port, ZN => n2859);
   U2202 : INV_X1 port map( A => REGISTERS_21_26_port, ZN => n2858);
   U2203 : INV_X1 port map( A => REGISTERS_21_27_port, ZN => n2857);
   U2204 : INV_X1 port map( A => REGISTERS_21_28_port, ZN => n2856);
   U2205 : INV_X1 port map( A => REGISTERS_21_29_port, ZN => n2855);
   U2206 : INV_X1 port map( A => REGISTERS_21_30_port, ZN => n2854);
   U2207 : INV_X1 port map( A => REGISTERS_21_31_port, ZN => n2853);
   U2208 : INV_X1 port map( A => REGISTERS_25_0_port, ZN => n3012);
   U2209 : INV_X1 port map( A => REGISTERS_3_0_port, ZN => n2436);
   U2210 : INV_X1 port map( A => REGISTERS_30_0_port, ZN => n3172);
   U2211 : INV_X1 port map( A => REGISTERS_26_0_port, ZN => n3044);
   U2212 : INV_X1 port map( A => REGISTERS_19_0_port, ZN => n2820);
   U2213 : INV_X1 port map( A => REGISTERS_16_0_port, ZN => n2724);
   U2214 : INV_X1 port map( A => REGISTERS_5_0_port, ZN => n2500);
   U2215 : INV_X1 port map( A => REGISTERS_25_1_port, ZN => n3011);
   U2216 : INV_X1 port map( A => REGISTERS_3_1_port, ZN => n2435);
   U2217 : INV_X1 port map( A => REGISTERS_30_1_port, ZN => n3171);
   U2218 : INV_X1 port map( A => REGISTERS_26_1_port, ZN => n3043);
   U2219 : INV_X1 port map( A => REGISTERS_19_1_port, ZN => n2819);
   U2220 : INV_X1 port map( A => REGISTERS_16_1_port, ZN => n2723);
   U2221 : INV_X1 port map( A => REGISTERS_5_1_port, ZN => n2499);
   U2222 : INV_X1 port map( A => REGISTERS_25_2_port, ZN => n3010);
   U2223 : INV_X1 port map( A => REGISTERS_3_2_port, ZN => n2434);
   U2224 : INV_X1 port map( A => REGISTERS_30_2_port, ZN => n3170);
   U2225 : INV_X1 port map( A => REGISTERS_26_2_port, ZN => n3042);
   U2226 : INV_X1 port map( A => REGISTERS_19_2_port, ZN => n2818);
   U2227 : INV_X1 port map( A => REGISTERS_16_2_port, ZN => n2722);
   U2228 : INV_X1 port map( A => REGISTERS_5_2_port, ZN => n2498);
   U2229 : INV_X1 port map( A => REGISTERS_25_3_port, ZN => n3009);
   U2230 : INV_X1 port map( A => REGISTERS_3_3_port, ZN => n2433);
   U2231 : INV_X1 port map( A => REGISTERS_30_3_port, ZN => n3169);
   U2232 : INV_X1 port map( A => REGISTERS_26_3_port, ZN => n3041);
   U2233 : INV_X1 port map( A => REGISTERS_19_3_port, ZN => n2817);
   U2234 : INV_X1 port map( A => REGISTERS_16_3_port, ZN => n2721);
   U2235 : INV_X1 port map( A => REGISTERS_5_3_port, ZN => n2497);
   U2236 : INV_X1 port map( A => REGISTERS_25_4_port, ZN => n3008);
   U2237 : INV_X1 port map( A => REGISTERS_3_4_port, ZN => n2432);
   U2238 : INV_X1 port map( A => REGISTERS_30_4_port, ZN => n3168);
   U2239 : INV_X1 port map( A => REGISTERS_26_4_port, ZN => n3040);
   U2240 : INV_X1 port map( A => REGISTERS_19_4_port, ZN => n2816);
   U2241 : INV_X1 port map( A => REGISTERS_16_4_port, ZN => n2720);
   U2242 : INV_X1 port map( A => REGISTERS_5_4_port, ZN => n2496);
   U2243 : INV_X1 port map( A => REGISTERS_25_5_port, ZN => n3007);
   U2244 : INV_X1 port map( A => REGISTERS_3_5_port, ZN => n2431);
   U2245 : INV_X1 port map( A => REGISTERS_30_5_port, ZN => n3167);
   U2246 : INV_X1 port map( A => REGISTERS_26_5_port, ZN => n3039);
   U2247 : INV_X1 port map( A => REGISTERS_19_5_port, ZN => n2815);
   U2248 : INV_X1 port map( A => REGISTERS_16_5_port, ZN => n2719);
   U2249 : INV_X1 port map( A => REGISTERS_5_5_port, ZN => n2495);
   U2250 : INV_X1 port map( A => REGISTERS_25_6_port, ZN => n3006);
   U2251 : INV_X1 port map( A => REGISTERS_3_6_port, ZN => n2430);
   U2252 : INV_X1 port map( A => REGISTERS_30_6_port, ZN => n3166);
   U2253 : INV_X1 port map( A => REGISTERS_26_6_port, ZN => n3038);
   U2254 : INV_X1 port map( A => REGISTERS_19_6_port, ZN => n2814);
   U2255 : INV_X1 port map( A => REGISTERS_16_6_port, ZN => n2718);
   U2256 : INV_X1 port map( A => REGISTERS_5_6_port, ZN => n2494);
   U2257 : INV_X1 port map( A => REGISTERS_25_7_port, ZN => n3005);
   U2258 : INV_X1 port map( A => REGISTERS_3_7_port, ZN => n2429);
   U2259 : INV_X1 port map( A => REGISTERS_30_7_port, ZN => n3165);
   U2260 : INV_X1 port map( A => REGISTERS_26_7_port, ZN => n3037);
   U2261 : INV_X1 port map( A => REGISTERS_19_7_port, ZN => n2813);
   U2262 : INV_X1 port map( A => REGISTERS_16_7_port, ZN => n2717);
   U2263 : INV_X1 port map( A => REGISTERS_5_7_port, ZN => n2493);
   U2264 : INV_X1 port map( A => REGISTERS_25_8_port, ZN => n3004);
   U2265 : INV_X1 port map( A => REGISTERS_3_8_port, ZN => n2428);
   U2266 : INV_X1 port map( A => REGISTERS_30_8_port, ZN => n3164);
   U2267 : INV_X1 port map( A => REGISTERS_26_8_port, ZN => n3036);
   U2268 : INV_X1 port map( A => REGISTERS_19_8_port, ZN => n2812);
   U2269 : INV_X1 port map( A => REGISTERS_16_8_port, ZN => n2716);
   U2270 : INV_X1 port map( A => REGISTERS_5_8_port, ZN => n2492);
   U2271 : INV_X1 port map( A => REGISTERS_25_9_port, ZN => n3003);
   U2272 : INV_X1 port map( A => REGISTERS_3_9_port, ZN => n2427);
   U2273 : INV_X1 port map( A => REGISTERS_30_9_port, ZN => n3163);
   U2274 : INV_X1 port map( A => REGISTERS_26_9_port, ZN => n3035);
   U2275 : INV_X1 port map( A => REGISTERS_19_9_port, ZN => n2811);
   U2276 : INV_X1 port map( A => REGISTERS_16_9_port, ZN => n2715);
   U2277 : INV_X1 port map( A => REGISTERS_5_9_port, ZN => n2491);
   U2278 : INV_X1 port map( A => REGISTERS_25_10_port, ZN => n3002);
   U2279 : INV_X1 port map( A => REGISTERS_3_10_port, ZN => n2426);
   U2280 : INV_X1 port map( A => REGISTERS_30_10_port, ZN => n3162);
   U2281 : INV_X1 port map( A => REGISTERS_26_10_port, ZN => n3034);
   U2282 : INV_X1 port map( A => REGISTERS_19_10_port, ZN => n2810);
   U2283 : INV_X1 port map( A => REGISTERS_16_10_port, ZN => n2714);
   U2284 : INV_X1 port map( A => REGISTERS_5_10_port, ZN => n2490);
   U2285 : INV_X1 port map( A => REGISTERS_25_11_port, ZN => n3001);
   U2286 : INV_X1 port map( A => REGISTERS_3_11_port, ZN => n2425);
   U2287 : INV_X1 port map( A => REGISTERS_30_11_port, ZN => n3161);
   U2288 : INV_X1 port map( A => REGISTERS_26_11_port, ZN => n3033);
   U2289 : INV_X1 port map( A => REGISTERS_19_11_port, ZN => n2809);
   U2290 : INV_X1 port map( A => REGISTERS_16_11_port, ZN => n2713);
   U2291 : INV_X1 port map( A => REGISTERS_5_11_port, ZN => n2489);
   U2292 : INV_X1 port map( A => REGISTERS_25_12_port, ZN => n3000);
   U2293 : INV_X1 port map( A => REGISTERS_3_12_port, ZN => n2424);
   U2294 : INV_X1 port map( A => REGISTERS_30_12_port, ZN => n3160);
   U2295 : INV_X1 port map( A => REGISTERS_26_12_port, ZN => n3032);
   U2296 : INV_X1 port map( A => REGISTERS_19_12_port, ZN => n2808);
   U2297 : INV_X1 port map( A => REGISTERS_16_12_port, ZN => n2712);
   U2298 : INV_X1 port map( A => REGISTERS_5_12_port, ZN => n2488);
   U2299 : INV_X1 port map( A => REGISTERS_25_13_port, ZN => n2999);
   U2300 : INV_X1 port map( A => REGISTERS_3_13_port, ZN => n2423);
   U2301 : INV_X1 port map( A => REGISTERS_30_13_port, ZN => n3159);
   U2302 : INV_X1 port map( A => REGISTERS_26_13_port, ZN => n3031);
   U2303 : INV_X1 port map( A => REGISTERS_19_13_port, ZN => n2807);
   U2304 : INV_X1 port map( A => REGISTERS_16_13_port, ZN => n2711);
   U2305 : INV_X1 port map( A => REGISTERS_5_13_port, ZN => n2487);
   U2306 : INV_X1 port map( A => REGISTERS_25_14_port, ZN => n2998);
   U2307 : INV_X1 port map( A => REGISTERS_3_14_port, ZN => n2422);
   U2308 : INV_X1 port map( A => REGISTERS_30_14_port, ZN => n3158);
   U2309 : INV_X1 port map( A => REGISTERS_26_14_port, ZN => n3030);
   U2310 : INV_X1 port map( A => REGISTERS_19_14_port, ZN => n2806);
   U2311 : INV_X1 port map( A => REGISTERS_16_14_port, ZN => n2710);
   U2312 : INV_X1 port map( A => REGISTERS_5_14_port, ZN => n2486);
   U2313 : INV_X1 port map( A => REGISTERS_25_15_port, ZN => n2997);
   U2314 : INV_X1 port map( A => REGISTERS_3_15_port, ZN => n2421);
   U2315 : INV_X1 port map( A => REGISTERS_30_15_port, ZN => n3157);
   U2316 : INV_X1 port map( A => REGISTERS_26_15_port, ZN => n3029);
   U2317 : INV_X1 port map( A => REGISTERS_19_15_port, ZN => n2805);
   U2318 : INV_X1 port map( A => REGISTERS_16_15_port, ZN => n2709);
   U2319 : INV_X1 port map( A => REGISTERS_5_15_port, ZN => n2485);
   U2320 : INV_X1 port map( A => REGISTERS_25_16_port, ZN => n2996);
   U2321 : INV_X1 port map( A => REGISTERS_3_16_port, ZN => n2420);
   U2322 : INV_X1 port map( A => REGISTERS_30_16_port, ZN => n3156);
   U2323 : INV_X1 port map( A => REGISTERS_26_16_port, ZN => n3028);
   U2324 : INV_X1 port map( A => REGISTERS_19_16_port, ZN => n2804);
   U2325 : INV_X1 port map( A => REGISTERS_16_16_port, ZN => n2708);
   U2326 : INV_X1 port map( A => REGISTERS_5_16_port, ZN => n2484);
   U2327 : INV_X1 port map( A => REGISTERS_25_17_port, ZN => n2995);
   U2328 : INV_X1 port map( A => REGISTERS_3_17_port, ZN => n2419);
   U2329 : INV_X1 port map( A => REGISTERS_30_17_port, ZN => n3155);
   U2330 : INV_X1 port map( A => REGISTERS_26_17_port, ZN => n3027);
   U2331 : INV_X1 port map( A => REGISTERS_19_17_port, ZN => n2803);
   U2332 : INV_X1 port map( A => REGISTERS_16_17_port, ZN => n2707);
   U2333 : INV_X1 port map( A => REGISTERS_5_17_port, ZN => n2483);
   U2334 : INV_X1 port map( A => REGISTERS_25_18_port, ZN => n2994);
   U2335 : INV_X1 port map( A => REGISTERS_3_18_port, ZN => n2418);
   U2336 : INV_X1 port map( A => REGISTERS_30_18_port, ZN => n3154);
   U2337 : INV_X1 port map( A => REGISTERS_26_18_port, ZN => n3026);
   U2338 : INV_X1 port map( A => REGISTERS_19_18_port, ZN => n2802);
   U2339 : INV_X1 port map( A => REGISTERS_16_18_port, ZN => n2706);
   U2340 : INV_X1 port map( A => REGISTERS_5_18_port, ZN => n2482);
   U2341 : INV_X1 port map( A => REGISTERS_25_19_port, ZN => n2993);
   U2342 : INV_X1 port map( A => REGISTERS_3_19_port, ZN => n2417);
   U2343 : INV_X1 port map( A => REGISTERS_30_19_port, ZN => n3153);
   U2344 : INV_X1 port map( A => REGISTERS_26_19_port, ZN => n3025);
   U2345 : INV_X1 port map( A => REGISTERS_19_19_port, ZN => n2801);
   U2346 : INV_X1 port map( A => REGISTERS_16_19_port, ZN => n2705);
   U2347 : INV_X1 port map( A => REGISTERS_5_19_port, ZN => n2481);
   U2348 : INV_X1 port map( A => REGISTERS_25_20_port, ZN => n2992);
   U2349 : INV_X1 port map( A => REGISTERS_3_20_port, ZN => n2416);
   U2350 : INV_X1 port map( A => REGISTERS_30_20_port, ZN => n3152);
   U2351 : INV_X1 port map( A => REGISTERS_26_20_port, ZN => n3024);
   U2352 : INV_X1 port map( A => REGISTERS_19_20_port, ZN => n2800);
   U2353 : INV_X1 port map( A => REGISTERS_16_20_port, ZN => n2704);
   U2354 : INV_X1 port map( A => REGISTERS_5_20_port, ZN => n2480);
   U2355 : INV_X1 port map( A => REGISTERS_25_21_port, ZN => n2991);
   U2356 : INV_X1 port map( A => REGISTERS_3_21_port, ZN => n2415);
   U2357 : INV_X1 port map( A => REGISTERS_30_21_port, ZN => n3151);
   U2358 : INV_X1 port map( A => REGISTERS_26_21_port, ZN => n3023);
   U2359 : INV_X1 port map( A => REGISTERS_19_21_port, ZN => n2799);
   U2360 : INV_X1 port map( A => REGISTERS_16_21_port, ZN => n2703);
   U2361 : INV_X1 port map( A => REGISTERS_5_21_port, ZN => n2479);
   U2362 : INV_X1 port map( A => REGISTERS_25_22_port, ZN => n2990);
   U2363 : INV_X1 port map( A => REGISTERS_3_22_port, ZN => n2414);
   U2364 : INV_X1 port map( A => REGISTERS_30_22_port, ZN => n3150);
   U2365 : INV_X1 port map( A => REGISTERS_26_22_port, ZN => n3022);
   U2366 : INV_X1 port map( A => REGISTERS_19_22_port, ZN => n2798);
   U2367 : INV_X1 port map( A => REGISTERS_16_22_port, ZN => n2702);
   U2368 : INV_X1 port map( A => REGISTERS_5_22_port, ZN => n2478);
   U2369 : INV_X1 port map( A => REGISTERS_25_23_port, ZN => n2989);
   U2370 : INV_X1 port map( A => REGISTERS_3_23_port, ZN => n2413);
   U2371 : INV_X1 port map( A => REGISTERS_30_23_port, ZN => n3149);
   U2372 : INV_X1 port map( A => REGISTERS_26_23_port, ZN => n3021);
   U2373 : INV_X1 port map( A => REGISTERS_19_23_port, ZN => n2797);
   U2374 : INV_X1 port map( A => REGISTERS_16_23_port, ZN => n2701);
   U2375 : INV_X1 port map( A => REGISTERS_5_23_port, ZN => n2477);
   U2376 : INV_X1 port map( A => REGISTERS_25_24_port, ZN => n2988);
   U2377 : INV_X1 port map( A => REGISTERS_3_24_port, ZN => n2412);
   U2378 : INV_X1 port map( A => REGISTERS_30_24_port, ZN => n3148);
   U2379 : INV_X1 port map( A => REGISTERS_26_24_port, ZN => n3020);
   U2380 : INV_X1 port map( A => REGISTERS_19_24_port, ZN => n2796);
   U2381 : INV_X1 port map( A => REGISTERS_16_24_port, ZN => n2700);
   U2382 : INV_X1 port map( A => REGISTERS_5_24_port, ZN => n2476);
   U2383 : INV_X1 port map( A => REGISTERS_25_25_port, ZN => n2987);
   U2384 : INV_X1 port map( A => REGISTERS_3_25_port, ZN => n2411);
   U2385 : INV_X1 port map( A => REGISTERS_30_25_port, ZN => n3147);
   U2386 : INV_X1 port map( A => REGISTERS_26_25_port, ZN => n3019);
   U2387 : INV_X1 port map( A => REGISTERS_19_25_port, ZN => n2795);
   U2388 : INV_X1 port map( A => REGISTERS_16_25_port, ZN => n2699);
   U2389 : INV_X1 port map( A => REGISTERS_5_25_port, ZN => n2475);
   U2390 : INV_X1 port map( A => REGISTERS_25_26_port, ZN => n2986);
   U2391 : INV_X1 port map( A => REGISTERS_3_26_port, ZN => n2410);
   U2392 : INV_X1 port map( A => REGISTERS_30_26_port, ZN => n3146);
   U2393 : INV_X1 port map( A => REGISTERS_26_26_port, ZN => n3018);
   U2394 : INV_X1 port map( A => REGISTERS_19_26_port, ZN => n2794);
   U2395 : INV_X1 port map( A => REGISTERS_16_26_port, ZN => n2698);
   U2396 : INV_X1 port map( A => REGISTERS_5_26_port, ZN => n2474);
   U2397 : INV_X1 port map( A => REGISTERS_25_27_port, ZN => n2985);
   U2398 : INV_X1 port map( A => REGISTERS_3_27_port, ZN => n2409);
   U2399 : INV_X1 port map( A => REGISTERS_30_27_port, ZN => n3145);
   U2400 : INV_X1 port map( A => REGISTERS_26_27_port, ZN => n3017);
   U2401 : INV_X1 port map( A => REGISTERS_19_27_port, ZN => n2793);
   U2402 : INV_X1 port map( A => REGISTERS_16_27_port, ZN => n2697);
   U2403 : INV_X1 port map( A => REGISTERS_5_27_port, ZN => n2473);
   U2404 : INV_X1 port map( A => REGISTERS_25_28_port, ZN => n2984);
   U2405 : INV_X1 port map( A => REGISTERS_3_28_port, ZN => n2408);
   U2406 : INV_X1 port map( A => REGISTERS_30_28_port, ZN => n3144);
   U2407 : INV_X1 port map( A => REGISTERS_26_28_port, ZN => n3016);
   U2408 : INV_X1 port map( A => REGISTERS_19_28_port, ZN => n2792);
   U2409 : INV_X1 port map( A => REGISTERS_16_28_port, ZN => n2696);
   U2410 : INV_X1 port map( A => REGISTERS_5_28_port, ZN => n2472);
   U2411 : INV_X1 port map( A => REGISTERS_25_29_port, ZN => n2983);
   U2412 : INV_X1 port map( A => REGISTERS_3_29_port, ZN => n2407);
   U2413 : INV_X1 port map( A => REGISTERS_30_29_port, ZN => n3143);
   U2414 : INV_X1 port map( A => REGISTERS_26_29_port, ZN => n3015);
   U2415 : INV_X1 port map( A => REGISTERS_19_29_port, ZN => n2791);
   U2416 : INV_X1 port map( A => REGISTERS_16_29_port, ZN => n2695);
   U2417 : INV_X1 port map( A => REGISTERS_5_29_port, ZN => n2471);
   U2418 : INV_X1 port map( A => REGISTERS_25_30_port, ZN => n2982);
   U2419 : INV_X1 port map( A => REGISTERS_3_30_port, ZN => n2406);
   U2420 : INV_X1 port map( A => REGISTERS_30_30_port, ZN => n3142);
   U2421 : INV_X1 port map( A => REGISTERS_26_30_port, ZN => n3014);
   U2422 : INV_X1 port map( A => REGISTERS_19_30_port, ZN => n2790);
   U2423 : INV_X1 port map( A => REGISTERS_16_30_port, ZN => n2694);
   U2424 : INV_X1 port map( A => REGISTERS_5_30_port, ZN => n2470);
   U2425 : INV_X1 port map( A => REGISTERS_25_31_port, ZN => n2981);
   U2426 : INV_X1 port map( A => REGISTERS_3_31_port, ZN => n2405);
   U2427 : INV_X1 port map( A => REGISTERS_30_31_port, ZN => n3141);
   U2428 : INV_X1 port map( A => REGISTERS_26_31_port, ZN => n3013);
   U2429 : INV_X1 port map( A => REGISTERS_19_31_port, ZN => n2789);
   U2430 : INV_X1 port map( A => REGISTERS_16_31_port, ZN => n2693);
   U2431 : INV_X1 port map( A => REGISTERS_5_31_port, ZN => n2469);
   U2432 : INV_X1 port map( A => ADD_WR(4), ZN => n3207);
   U2433 : INV_X1 port map( A => ADD_WR(3), ZN => n3208);
   U2434 : INV_X1 port map( A => CLK, ZN => n3220);
   U2435 : INV_X1 port map( A => ADD_RD2(3), ZN => n3217);
   U2436 : NOR2_X1 port map( A1 => n3216, A2 => ADD_RD2(3), ZN => n1418);
   U2437 : INV_X1 port map( A => ADD_RD2(1), ZN => n3218);
   U2438 : INV_X1 port map( A => ADD_RD1(1), ZN => n3214);
   U2439 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n3215, 
                           ZN => n1451);
   U2440 : INV_X1 port map( A => ADD_RD1(4), ZN => n3212);
   U2441 : NOR2_X1 port map( A1 => n3213, A2 => ADD_RD1(4), ZN => n1446);
   U2442 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1922);
   U2443 : INV_X1 port map( A => ADD_RD2(4), ZN => n3216);
   U2444 : NOR2_X1 port map( A1 => n3217, A2 => ADD_RD2(4), ZN => n931);
   U2445 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1407);
   U2446 : INV_X1 port map( A => ADD_RD1(0), ZN => n3215);
   U2447 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n3214, 
                           ZN => n1455);
   U2448 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n1456);
   U2449 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n3219, 
                           ZN => n936);
   U2450 : NOR3_X1 port map( A1 => n3218, A2 => ADD_RD2(2), A3 => n3219, ZN => 
                           n935);
   U2451 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n3218, 
                           ZN => n940);
   U2452 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n941);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CWBU is

   port( CLOCK : in std_logic;  ALU_OP : in std_logic_vector (0 to 4);  PSW : 
         in std_logic_vector (6 downto 0);  COND_SEL : out std_logic_vector (1 
         downto 0);  CWB_SEL : in std_logic_vector (1 downto 0);  CWB_MUW_SEL :
         out std_logic_vector (1 downto 0));

end CWBU;

architecture SYN_BEHAVIORAL of CWBU is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n4, n5, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n11, n12, n26, n27, n28, n29, n30, n31, n32, n_1533, n_1534 : 
      std_logic;

begin
   
   ALUPIPE_reg_3_inst : DFF_X1 port map( D => ALU_OP(1), CK => CLOCK, Q => n25,
                           QN => n26);
   ALUPIPE_reg_1_inst : DFF_X1 port map( D => ALU_OP(3), CK => CLOCK, Q => n11,
                           QN => n4);
   ALUPIPE_reg_4_inst : DFF_X1 port map( D => ALU_OP(0), CK => CLOCK, Q => 
                           n_1533, QN => n1);
   ALUPIPE_reg_0_inst : DFF_X1 port map( D => ALU_OP(4), CK => CLOCK, Q => 
                           n_1534, QN => n5);
   ALUPIPE_reg_2_inst : DFF_X1 port map( D => ALU_OP(2), CK => CLOCK, Q => n12,
                           QN => n24);
   U25 : NAND3_X1 port map( A1 => n32, A2 => n13, A3 => n14, ZN => 
                           CWB_MUW_SEL(1));
   U26 : NAND3_X1 port map( A1 => n25, A2 => n1, A3 => n24, ZN => n13);
   U3 : INV_X1 port map( A => CWB_SEL(1), ZN => n32);
   U4 : AOI221_X1 port map( B1 => PSW(3), B2 => n16, C1 => n5, C2 => n28, A => 
                           n22, ZN => n21);
   U5 : INV_X1 port map( A => n23, ZN => n28);
   U6 : NOR3_X1 port map( A1 => n31, A2 => n5, A3 => n11, ZN => n22);
   U7 : AOI22_X1 port map( A1 => n11, A2 => PSW(1), B1 => n4, B2 => PSW(0), ZN 
                           => n23);
   U8 : AOI221_X1 port map( B1 => n16, B2 => n30, C1 => n5, C2 => n19, A => n20
                           , ZN => n18);
   U9 : INV_X1 port map( A => PSW(3), ZN => n30);
   U10 : NOR3_X1 port map( A1 => n11, A2 => n5, A3 => PSW(2), ZN => n20);
   U11 : OAI22_X1 port map( A1 => n4, A2 => PSW(1), B1 => PSW(0), B2 => n11, ZN
                           => n19);
   U12 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n16);
   U13 : NAND4_X1 port map( A1 => n16, A2 => n1, A3 => n26, A4 => n12, ZN => 
                           n14);
   U14 : AND2_X1 port map( A1 => CWB_SEL(0), A2 => n15, ZN => CWB_MUW_SEL(0));
   U15 : OAI211_X1 port map( C1 => n16, C2 => n27, A => n1, B => n17, ZN => n15
                           );
   U16 : INV_X1 port map( A => n13, ZN => n27);
   U17 : XNOR2_X1 port map( A => n25, B => n24, ZN => n17);
   U18 : OAI22_X1 port map( A1 => n14, A2 => n29, B1 => n21, B2 => n13, ZN => 
                           COND_SEL(0));
   U19 : OAI22_X1 port map( A1 => PSW(5), A2 => n14, B1 => n18, B2 => n13, ZN 
                           => COND_SEL(1));
   U20 : INV_X1 port map( A => PSW(2), ZN => n31);
   U21 : INV_X1 port map( A => PSW(5), ZN => n29);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 is

   port( clock, rst : in std_logic;  address : in std_logic_vector (31 downto 
         0);  d_in, w_en : in std_logic;  d_out : out std_logic);

end BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0;

architecture SYN_Behavioral of BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n24, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
      n81, n82, net60602, net62447, net60531, net62449, net62444, n35, n88, n29
      , n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n83, n84, d_out_port, n91, n92,
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n_1535, n_1536, n_1537, n_1538, n_1539, 
      n_1540, n_1541, n_1542 : std_logic;

begin
   d_out <= d_out_port;
   
   BHT_reg_7_0_inst : DFFR_X1 port map( D => n68, CK => n122, RN => n97, Q => 
                           n_1535, QN => n24);
   BHT_reg_2_1_inst : DFFR_X1 port map( D => n78, CK => n122, RN => n98, Q => 
                           n_1536, QN => net60602);
   BHT_reg_1_1_inst : DFFR_X1 port map( D => n80, CK => n122, RN => n97, Q => 
                           n108, QN => net62449);
   BHT_reg_7_1_inst : DFFR_X1 port map( D => n88, CK => n122, RN => n98, Q => 
                           n_1537, QN => n67);
   BHT_reg_0_0_inst : DFFR_X1 port map( D => n81, CK => n122, RN => n98, Q => 
                           n109, QN => n64);
   BHT_reg_4_1_inst : DFFR_X1 port map( D => n74, CK => n122, RN => n97, Q => 
                           n112, QN => n62);
   BHT_reg_6_0_inst : DFFR_X1 port map( D => n69, CK => n122, RN => n97, Q => 
                           n_1538, QN => n83);
   BHT_reg_3_0_inst : DFFR_X1 port map( D => n75, CK => n122, RN => n97, Q => 
                           n_1539, QN => n65);
   BHT_reg_6_1_inst : DFFR_X1 port map( D => n70, CK => n122, RN => n97, Q => 
                           n_1540, QN => n84);
   BHT_reg_3_1_inst : DFFR_X1 port map( D => n76, CK => n122, RN => n97, Q => 
                           n_1541, QN => n61);
   BHT_reg_5_1_inst : DFFR_X1 port map( D => n72, CK => n122, RN => n97, Q => 
                           n113, QN => n35);
   BHT_reg_5_0_inst : DFFR_X1 port map( D => n71, CK => n122, RN => n97, Q => 
                           n114, QN => net62447);
   BHT_reg_2_0_inst : DFFR_X1 port map( D => n77, CK => n122, RN => n97, Q => 
                           n_1542, QN => n66);
   BHT_reg_1_0_inst : DFFR_X1 port map( D => n79, CK => n122, RN => n97, Q => 
                           n115, QN => net62444);
   U70 : NAND3_X1 port map( A1 => n119, A2 => n117, A3 => n37, ZN => n36);
   U71 : NAND3_X1 port map( A1 => address(1), A2 => n117, A3 => n39, ZN => n38)
                           ;
   U72 : NAND3_X1 port map( A1 => address(1), A2 => n117, A3 => n37, ZN => n40)
                           ;
   U73 : NAND3_X1 port map( A1 => address(2), A2 => n119, A3 => n37, ZN => n42)
                           ;
   U75 : NAND3_X1 port map( A1 => address(2), A2 => address(1), A3 => n39, ZN 
                           => n44);
   U76 : NAND3_X1 port map( A1 => address(2), A2 => n120, A3 => w_en, ZN => n47
                           );
   BHT_reg_4_0_inst : DFFR_X1 port map( D => n73, CK => n122, RN => n98, Q => 
                           n110, QN => n63);
   BHT_reg_0_1_inst : DFFR_X1 port map( D => n82, CK => n122, RN => n97, Q => 
                           n111, QN => n60);
   U3 : BUF_X1 port map( A => rst, Z => n99);
   U4 : INV_X1 port map( A => n107, ZN => d_out_port);
   U5 : INV_X1 port map( A => n99, ZN => n97);
   U6 : INV_X1 port map( A => n99, ZN => n98);
   U7 : AND3_X1 port map( A1 => w_en, A2 => n121, A3 => n43, ZN => n39);
   U8 : NAND2_X1 port map( A1 => address(1), A2 => address(0), ZN => n53);
   U9 : NOR2_X1 port map( A1 => address(0), A2 => address(1), ZN => n50);
   U10 : NOR2_X1 port map( A1 => n121, A2 => address(1), ZN => n51);
   U11 : INV_X1 port map( A => address(2), ZN => n117);
   U12 : BUF_X1 port map( A => n33, Z => n92);
   U13 : INV_X1 port map( A => n53, ZN => n120);
   U14 : OAI22_X1 port map( A1 => n56, A2 => n117, B1 => address(2), B2 => n57,
                           ZN => net60531);
   U15 : AOI221_X1 port map( B1 => n50, B2 => n112, C1 => n51, C2 => n113, A =>
                           n59, ZN => n56);
   U16 : AOI221_X1 port map( B1 => n50, B2 => n111, C1 => n51, C2 => n108, A =>
                           n58, ZN => n57);
   U17 : OR2_X1 port map( A1 => n30, A2 => n91, ZN => n88);
   U18 : AND3_X1 port map( A1 => d_in, A2 => n29, A3 => n118, ZN => n91);
   U19 : AOI21_X1 port map( B1 => n106, B2 => n118, A => n67, ZN => n30);
   U20 : OAI21_X1 port map( B1 => n24, B2 => n45, A => n46, ZN => n68);
   U21 : INV_X1 port map( A => clock, ZN => n122);
   U22 : OAI22_X1 port map( A1 => n48, A2 => n117, B1 => address(2), B2 => n49,
                           ZN => n33);
   U23 : INV_X1 port map( A => n36, ZN => n105);
   U24 : INV_X1 port map( A => n42, ZN => n103);
   U25 : INV_X1 port map( A => n40, ZN => n104);
   U26 : INV_X1 port map( A => n44, ZN => n101);
   U27 : INV_X1 port map( A => n38, ZN => n102);
   U28 : XOR2_X1 port map( A => n29, B => d_in, Z => n93);
   U29 : XOR2_X1 port map( A => n29, B => d_in, Z => n94);
   U30 : AND2_X1 port map( A1 => n117, A2 => n119, ZN => n95);
   U31 : INV_X1 port map( A => address(1), ZN => n119);
   U32 : AND2_X1 port map( A1 => n34, A2 => address(2), ZN => n96);
   U33 : NAND2_X1 port map( A1 => n34, A2 => address(2), ZN => n41);
   U34 : AND2_X1 port map( A1 => n39, A2 => n119, ZN => n34);
   U35 : NAND2_X1 port map( A1 => n95, A2 => n39, ZN => n32);
   U36 : OAI222_X1 port map( A1 => d_in, A2 => n106, B1 => n107, B2 => n33, C1 
                           => net60531, C2 => n116, ZN => n43);
   U37 : INV_X1 port map( A => n47, ZN => n118);
   U38 : INV_X1 port map( A => address(0), ZN => n121);
   U39 : INV_X1 port map( A => n32, ZN => n100);
   U40 : OAI22_X1 port map( A1 => n100, A2 => n60, B1 => n31, B2 => n32, ZN => 
                           n82);
   U41 : NAND2_X1 port map( A1 => address(1), A2 => n121, ZN => n54);
   U42 : XOR2_X1 port map( A => n29, B => d_in, Z => n31);
   U43 : INV_X1 port map( A => d_in, ZN => n116);
   U44 : AOI221_X1 port map( B1 => n50, B2 => n110, C1 => n51, C2 => n114, A =>
                           n55, ZN => n48);
   U45 : AOI21_X1 port map( B1 => d_in, B2 => d_out_port, A => n47, ZN => n45);
   U46 : OAI211_X1 port map( C1 => d_in, C2 => d_out_port, A => n106, B => n118
                           , ZN => n46);
   U47 : AND3_X1 port map( A1 => n43, A2 => address(0), A3 => w_en, ZN => n37);
   U48 : XNOR2_X1 port map( A => n106, B => d_out_port, ZN => n29);
   U49 : INV_X1 port map( A => net60531, ZN => n107);
   U50 : OAI22_X1 port map( A1 => n67, A2 => n53, B1 => n84, B2 => n54, ZN => 
                           n59);
   U51 : OAI22_X1 port map( A1 => n24, A2 => n53, B1 => n83, B2 => n54, ZN => 
                           n55);
   U52 : OAI22_X1 port map( A1 => n65, A2 => n53, B1 => n66, B2 => n54, ZN => 
                           n52);
   U53 : OAI22_X1 port map( A1 => n61, A2 => n53, B1 => net60602, B2 => n54, ZN
                           => n58);
   U54 : OAI22_X1 port map( A1 => n100, A2 => n64, B1 => n92, B2 => n32, ZN => 
                           n81);
   U55 : OAI22_X1 port map( A1 => net62444, A2 => n105, B1 => n92, B2 => n36, 
                           ZN => n79);
   U56 : OAI22_X1 port map( A1 => n66, A2 => n102, B1 => n92, B2 => n38, ZN => 
                           n77);
   U57 : OAI22_X1 port map( A1 => n65, A2 => n104, B1 => n92, B2 => n40, ZN => 
                           n75);
   U58 : OAI22_X1 port map( A1 => n96, A2 => n63, B1 => n41, B2 => n92, ZN => 
                           n73);
   U59 : OAI22_X1 port map( A1 => net62447, A2 => n103, B1 => n92, B2 => n42, 
                           ZN => n71);
   U60 : OAI22_X1 port map( A1 => n83, A2 => n101, B1 => n92, B2 => n44, ZN => 
                           n69);
   U61 : OAI22_X1 port map( A1 => n35, A2 => n103, B1 => n94, B2 => n42, ZN => 
                           n72);
   U62 : OAI22_X1 port map( A1 => n84, A2 => n101, B1 => n93, B2 => n44, ZN => 
                           n70);
   U63 : OAI22_X1 port map( A1 => n62, A2 => n96, B1 => n41, B2 => n31, ZN => 
                           n74);
   U64 : OAI22_X1 port map( A1 => n61, A2 => n104, B1 => n94, B2 => n40, ZN => 
                           n76);
   U65 : OAI22_X1 port map( A1 => net60602, A2 => n102, B1 => n93, B2 => n38, 
                           ZN => n78);
   U66 : OAI22_X1 port map( A1 => net62449, A2 => n105, B1 => n31, B2 => n36, 
                           ZN => n80);
   U67 : INV_X1 port map( A => n33, ZN => n106);
   U68 : AOI221_X1 port map( B1 => n50, B2 => n109, C1 => n51, C2 => n115, A =>
                           n52, ZN => n49);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HDU_IR_SIZE32 is

   port( clk, rst : in std_logic;  IR : in std_logic_vector (31 downto 0);  
         STALL_CODE : out std_logic_vector (1 downto 0);  IF_STALL, ID_STALL, 
         EX_STALL, MEM_STALL, WB_STALL : out std_logic);

end HDU_IR_SIZE32;

architecture SYN_behavioural of HDU_IR_SIZE32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal STALL_CODE_1_port, IF_STALL_port, EX_STALL_port, cnt_mul_30_port, 
      cnt_mul_29_port, cnt_mul_28_port, cnt_mul_27_port, cnt_mul_26_port, 
      cnt_mul_25_port, cnt_mul_24_port, cnt_mul_23_port, cnt_mul_22_port, 
      cnt_mul_21_port, cnt_mul_20_port, cnt_mul_19_port, cnt_mul_18_port, 
      cnt_mul_17_port, cnt_mul_16_port, cnt_mul_15_port, cnt_mul_14_port, 
      cnt_mul_13_port, cnt_mul_12_port, cnt_mul_11_port, cnt_mul_10_port, 
      cnt_mul_9_port, cnt_mul_8_port, cnt_mul_7_port, cnt_mul_6_port, 
      cnt_mul_5_port, cnt_mul_4_port, cnt_mul_3_port, cnt_mul_2_port, 
      cnt_mul_1_port, cnt_mul_0_port, N154, N155, N156, N157, N158, N159, N160,
      N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, 
      N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, 
      n98, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n149, n150, n151, n152, n153, 
      n155_port, n156_port, n157_port, n158_port, n159_port, n169_port, 
      n170_port, n171_port, n172_port, n173_port, n174_port, n175_port, 
      n176_port, n177_port, n178_port, n179_port, n180_port, n181_port, 
      n182_port, n183_port, n184_port, n185, n186, n187, n188, n189, n190, n191
      , n192, n193, n194, n195, n196, n197, n199, n200, n202, n93, n51, n52, 
      n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97, n100, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n154_port, n160_port, 
      STALL_CODE_0_port, n162_port, n163_port, n164_port, n165_port, n166_port,
      n167_port, n168_port, n198, n201, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555 : 
      std_logic;

begin
   STALL_CODE <= ( STALL_CODE_1_port, STALL_CODE_0_port );
   IF_STALL <= IF_STALL_port;
   ID_STALL <= IF_STALL_port;
   EX_STALL <= EX_STALL_port;
   MEM_STALL <= EX_STALL_port;
   WB_STALL <= EX_STALL_port;
   
   IR_EX_reg_31_inst : DFFR_X1 port map( D => n159_port, CK => clk, RN => 
                           n160_port, Q => n_1543, QN => n130);
   IR_EX_reg_30_inst : DFFR_X1 port map( D => n158_port, CK => clk, RN => 
                           n160_port, Q => n_1544, QN => n132);
   IR_EX_reg_29_inst : DFFR_X1 port map( D => n157_port, CK => clk, RN => 
                           n160_port, Q => n_1545, QN => n131);
   IR_EX_reg_28_inst : DFFR_X1 port map( D => n156_port, CK => clk, RN => 
                           n160_port, Q => n_1546, QN => n139);
   IR_EX_reg_27_inst : DFFR_X1 port map( D => n155_port, CK => clk, RN => 
                           n160_port, Q => n_1547, QN => n138);
   IR_EX_reg_26_inst : DFFR_X1 port map( D => n163_port, CK => clk, RN => 
                           n160_port, Q => n93, QN => n_1548);
   IR_EX_reg_20_inst : DFFR_X1 port map( D => n153, CK => clk, RN => n160_port,
                           Q => n_1549, QN => n135);
   IR_EX_reg_19_inst : DFFR_X1 port map( D => n152, CK => clk, RN => n160_port,
                           Q => n_1550, QN => n137);
   IR_EX_reg_18_inst : DFFR_X1 port map( D => n151, CK => clk, RN => n160_port,
                           Q => n_1551, QN => n136);
   IR_EX_reg_17_inst : DFFR_X1 port map( D => n150, CK => clk, RN => n160_port,
                           Q => n_1552, QN => n134);
   IR_EX_reg_16_inst : DFFR_X1 port map( D => n149, CK => clk, RN => n160_port,
                           Q => n_1553, QN => n133);
   cnt_mul_reg_1_inst : DFF_X1 port map( D => n200, CK => clk, Q => 
                           cnt_mul_1_port, QN => n100);
   cnt_mul_reg_5_inst : DFF_X1 port map( D => n194, CK => clk, Q => 
                           cnt_mul_5_port, QN => n104);
   cnt_mul_reg_4_inst : DFF_X1 port map( D => n195, CK => clk, Q => 
                           cnt_mul_4_port, QN => n103);
   cnt_mul_reg_3_inst : DFF_X1 port map( D => n196, CK => clk, Q => 
                           cnt_mul_3_port, QN => n102);
   cnt_mul_reg_2_inst : DFF_X1 port map( D => n197, CK => clk, Q => 
                           cnt_mul_2_port, QN => n101);
   cnt_mul_reg_30_inst : DFF_X1 port map( D => n169_port, CK => clk, Q => 
                           cnt_mul_30_port, QN => n129);
   cnt_mul_reg_29_inst : DFF_X1 port map( D => n170_port, CK => clk, Q => 
                           cnt_mul_29_port, QN => n128);
   cnt_mul_reg_28_inst : DFF_X1 port map( D => n171_port, CK => clk, Q => 
                           cnt_mul_28_port, QN => n127);
   cnt_mul_reg_27_inst : DFF_X1 port map( D => n172_port, CK => clk, Q => 
                           cnt_mul_27_port, QN => n126);
   cnt_mul_reg_26_inst : DFF_X1 port map( D => n173_port, CK => clk, Q => 
                           cnt_mul_26_port, QN => n125);
   cnt_mul_reg_25_inst : DFF_X1 port map( D => n174_port, CK => clk, Q => 
                           cnt_mul_25_port, QN => n124);
   cnt_mul_reg_24_inst : DFF_X1 port map( D => n175_port, CK => clk, Q => 
                           cnt_mul_24_port, QN => n123);
   cnt_mul_reg_23_inst : DFF_X1 port map( D => n176_port, CK => clk, Q => 
                           cnt_mul_23_port, QN => n122);
   cnt_mul_reg_22_inst : DFF_X1 port map( D => n177_port, CK => clk, Q => 
                           cnt_mul_22_port, QN => n121);
   cnt_mul_reg_21_inst : DFF_X1 port map( D => n178_port, CK => clk, Q => 
                           cnt_mul_21_port, QN => n120);
   cnt_mul_reg_20_inst : DFF_X1 port map( D => n179_port, CK => clk, Q => 
                           cnt_mul_20_port, QN => n119);
   cnt_mul_reg_19_inst : DFF_X1 port map( D => n180_port, CK => clk, Q => 
                           cnt_mul_19_port, QN => n118);
   cnt_mul_reg_18_inst : DFF_X1 port map( D => n181_port, CK => clk, Q => 
                           cnt_mul_18_port, QN => n117);
   cnt_mul_reg_17_inst : DFF_X1 port map( D => n182_port, CK => clk, Q => 
                           cnt_mul_17_port, QN => n116);
   cnt_mul_reg_16_inst : DFF_X1 port map( D => n183_port, CK => clk, Q => 
                           cnt_mul_16_port, QN => n115);
   cnt_mul_reg_15_inst : DFF_X1 port map( D => n184_port, CK => clk, Q => 
                           cnt_mul_15_port, QN => n114);
   cnt_mul_reg_14_inst : DFF_X1 port map( D => n185, CK => clk, Q => 
                           cnt_mul_14_port, QN => n113);
   cnt_mul_reg_13_inst : DFF_X1 port map( D => n186, CK => clk, Q => 
                           cnt_mul_13_port, QN => n112);
   cnt_mul_reg_12_inst : DFF_X1 port map( D => n187, CK => clk, Q => 
                           cnt_mul_12_port, QN => n111);
   cnt_mul_reg_11_inst : DFF_X1 port map( D => n188, CK => clk, Q => 
                           cnt_mul_11_port, QN => n110);
   cnt_mul_reg_10_inst : DFF_X1 port map( D => n189, CK => clk, Q => 
                           cnt_mul_10_port, QN => n109);
   cnt_mul_reg_9_inst : DFF_X1 port map( D => n190, CK => clk, Q => 
                           cnt_mul_9_port, QN => n108);
   cnt_mul_reg_31_inst : DFF_X1 port map( D => n164_port, CK => clk, Q => n227,
                           QN => n_1554);
   cnt_mul_reg_0_inst : DFF_X1 port map( D => n202, CK => clk, Q => 
                           cnt_mul_0_port, QN => n98);
   cnt_mul_reg_8_inst : DFF_X1 port map( D => n191, CK => clk, Q => 
                           cnt_mul_8_port, QN => n107);
   cnt_mul_reg_7_inst : DFF_X1 port map( D => n192, CK => clk, Q => 
                           cnt_mul_7_port, QN => n106);
   cnt_mul_reg_6_inst : DFF_X1 port map( D => n193, CK => clk, Q => 
                           cnt_mul_6_port, QN => n105);
   U139 : NAND3_X1 port map( A1 => n229, A2 => n228, A3 => n230, ZN => n83);
   U140 : XOR2_X1 port map( A => n136, B => IR(23), Z => n90);
   U141 : XOR2_X1 port map( A => n137, B => IR(24), Z => n88);
   r100 : HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1 port map( A(31) => n227, A(30) =>
                           cnt_mul_30_port, A(29) => cnt_mul_29_port, A(28) => 
                           cnt_mul_28_port, A(27) => cnt_mul_27_port, A(26) => 
                           cnt_mul_26_port, A(25) => cnt_mul_25_port, A(24) => 
                           cnt_mul_24_port, A(23) => cnt_mul_23_port, A(22) => 
                           cnt_mul_22_port, A(21) => cnt_mul_21_port, A(20) => 
                           cnt_mul_20_port, A(19) => cnt_mul_19_port, A(18) => 
                           cnt_mul_18_port, A(17) => cnt_mul_17_port, A(16) => 
                           cnt_mul_16_port, A(15) => cnt_mul_15_port, A(14) => 
                           cnt_mul_14_port, A(13) => cnt_mul_13_port, A(12) => 
                           cnt_mul_12_port, A(11) => cnt_mul_11_port, A(10) => 
                           cnt_mul_10_port, A(9) => cnt_mul_9_port, A(8) => 
                           cnt_mul_8_port, A(7) => cnt_mul_7_port, A(6) => 
                           cnt_mul_6_port, A(5) => cnt_mul_5_port, A(4) => 
                           cnt_mul_4_port, A(3) => cnt_mul_3_port, A(2) => 
                           cnt_mul_2_port, A(1) => cnt_mul_1_port, A(0) => 
                           cnt_mul_0_port, SUM(31) => N184, SUM(30) => N183, 
                           SUM(29) => N182, SUM(28) => N181, SUM(27) => N180, 
                           SUM(26) => N179, SUM(25) => N178, SUM(24) => N177, 
                           SUM(23) => N176, SUM(22) => N175, SUM(21) => N174, 
                           SUM(20) => N173, SUM(19) => N172, SUM(18) => N171, 
                           SUM(17) => N170, SUM(16) => N169, SUM(15) => N168, 
                           SUM(14) => N167, SUM(13) => N166, SUM(12) => N165, 
                           SUM(11) => N164, SUM(10) => N163, SUM(9) => N162, 
                           SUM(8) => N161, SUM(7) => N160, SUM(6) => N159, 
                           SUM(5) => N158, SUM(4) => N157, SUM(3) => N156, 
                           SUM(2) => N155, SUM(1) => N154, SUM(0) => n_1555);
   STALL_MUL_reg : DFF_X1 port map( D => n145, CK => clk, Q => EX_STALL_port, 
                           QN => n199);
   U3 : BUF_X1 port map( A => n140, Z => n144);
   U4 : BUF_X1 port map( A => n141, Z => n148);
   U5 : AND2_X1 port map( A1 => n54, A2 => n146, ZN => n140);
   U6 : INV_X1 port map( A => n144, ZN => n142);
   U7 : INV_X1 port map( A => n144, ZN => n143);
   U8 : INV_X1 port map( A => n148, ZN => n146);
   U9 : BUF_X1 port map( A => n140, Z => n145);
   U10 : INV_X1 port map( A => n148, ZN => n147);
   U11 : INV_X1 port map( A => rst, ZN => n160_port);
   U12 : INV_X1 port map( A => n74, ZN => STALL_CODE_0_port);
   U13 : BUF_X1 port map( A => n141, Z => n154_port);
   U14 : OR2_X1 port map( A1 => n54, A2 => n154_port, ZN => n52);
   U15 : AND2_X1 port map( A1 => n199, A2 => n57, ZN => n141);
   U16 : OAI22_X1 port map( A1 => n142, A2 => n212, B1 => n117, B2 => n147, ZN 
                           => n181_port);
   U17 : INV_X1 port map( A => N171, ZN => n212);
   U18 : OAI22_X1 port map( A1 => n143, A2 => n217, B1 => n121, B2 => n146, ZN 
                           => n177_port);
   U19 : INV_X1 port map( A => N175, ZN => n217);
   U20 : OAI22_X1 port map( A1 => n142, A2 => n204, B1 => n108, B2 => n147, ZN 
                           => n190);
   U21 : INV_X1 port map( A => N162, ZN => n204);
   U22 : OAI22_X1 port map( A1 => n142, A2 => n208, B1 => n112, B2 => n147, ZN 
                           => n186);
   U23 : INV_X1 port map( A => N166, ZN => n208);
   U24 : OAI22_X1 port map( A1 => n142, A2 => n225, B1 => n116, B2 => n147, ZN 
                           => n182_port);
   U25 : INV_X1 port map( A => N170, ZN => n225);
   U26 : OAI22_X1 port map( A1 => n143, A2 => n223, B1 => n128, B2 => n146, ZN 
                           => n170_port);
   U27 : INV_X1 port map( A => N182, ZN => n223);
   U28 : OAI22_X1 port map( A1 => n142, A2 => n201, B1 => n107, B2 => n147, ZN 
                           => n191);
   U29 : INV_X1 port map( A => N161, ZN => n201);
   U30 : OAI22_X1 port map( A1 => n142, A2 => n207, B1 => n111, B2 => n147, ZN 
                           => n187);
   U31 : INV_X1 port map( A => N165, ZN => n207);
   U32 : OAI22_X1 port map( A1 => n142, A2 => n210, B1 => n115, B2 => n147, ZN 
                           => n183_port);
   U33 : INV_X1 port map( A => N169, ZN => n210);
   U34 : OAI22_X1 port map( A1 => n143, A2 => n221, B1 => n127, B2 => n146, ZN 
                           => n171_port);
   U35 : INV_X1 port map( A => N181, ZN => n221);
   U36 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           n57);
   U37 : NOR4_X1 port map( A1 => IR(4), A2 => IR(31), A3 => IR(30), A4 => 
                           IR(29), ZN => n61);
   U38 : NOR4_X1 port map( A1 => n63, A2 => IR(7), A3 => IR(9), A4 => IR(8), ZN
                           => n62);
   U39 : OR2_X1 port map( A1 => IR(6), A2 => IR(5), ZN => n63);
   U40 : OAI22_X1 port map( A1 => n143, A2 => n214, B1 => n118, B2 => n147, ZN 
                           => n180_port);
   U41 : INV_X1 port map( A => N172, ZN => n214);
   U42 : OAI22_X1 port map( A1 => n143, A2 => n216, B1 => n122, B2 => n146, ZN 
                           => n176_port);
   U43 : INV_X1 port map( A => N176, ZN => n216);
   U44 : OAI22_X1 port map( A1 => n142, A2 => n198, B1 => n106, B2 => n147, ZN 
                           => n192);
   U45 : INV_X1 port map( A => N160, ZN => n198);
   U46 : OAI22_X1 port map( A1 => n142, A2 => n206, B1 => n110, B2 => n147, ZN 
                           => n188);
   U47 : INV_X1 port map( A => N164, ZN => n206);
   U48 : OAI22_X1 port map( A1 => n142, A2 => n211, B1 => n114, B2 => n147, ZN 
                           => n184_port);
   U49 : INV_X1 port map( A => N168, ZN => n211);
   U50 : OAI22_X1 port map( A1 => n143, A2 => n222, B1 => n126, B2 => n146, ZN 
                           => n172_port);
   U51 : INV_X1 port map( A => N180, ZN => n222);
   U52 : OAI22_X1 port map( A1 => n142, A2 => n205, B1 => n109, B2 => n147, ZN 
                           => n189);
   U53 : INV_X1 port map( A => N163, ZN => n205);
   U54 : OAI22_X1 port map( A1 => n142, A2 => n209, B1 => n113, B2 => n147, ZN 
                           => n185);
   U55 : INV_X1 port map( A => N167, ZN => n209);
   U56 : OAI22_X1 port map( A1 => n143, A2 => n213, B1 => n119, B2 => n146, ZN 
                           => n179_port);
   U57 : INV_X1 port map( A => N173, ZN => n213);
   U58 : OAI22_X1 port map( A1 => n142, A2 => n215, B1 => n120, B2 => n146, ZN 
                           => n178_port);
   U59 : INV_X1 port map( A => N174, ZN => n215);
   U60 : OAI22_X1 port map( A1 => n143, A2 => n219, B1 => n123, B2 => n146, ZN 
                           => n175_port);
   U61 : INV_X1 port map( A => N177, ZN => n219);
   U62 : OAI22_X1 port map( A1 => n142, A2 => n218, B1 => n124, B2 => n146, ZN 
                           => n174_port);
   U63 : INV_X1 port map( A => N178, ZN => n218);
   U64 : OAI22_X1 port map( A1 => n143, A2 => n220, B1 => n125, B2 => n146, ZN 
                           => n173_port);
   U65 : INV_X1 port map( A => N179, ZN => n220);
   U66 : OAI22_X1 port map( A1 => n142, A2 => n224, B1 => n129, B2 => n146, ZN 
                           => n169_port);
   U67 : INV_X1 port map( A => N183, ZN => n224);
   U68 : OAI22_X1 port map( A1 => n143, A2 => n203, B1 => n104, B2 => n147, ZN 
                           => n194);
   U69 : INV_X1 port map( A => N158, ZN => n203);
   U70 : OAI22_X1 port map( A1 => n143, A2 => n226, B1 => n103, B2 => n147, ZN 
                           => n195);
   U71 : INV_X1 port map( A => N157, ZN => n226);
   U72 : OAI22_X1 port map( A1 => n143, A2 => n167_port, B1 => n102, B2 => n147
                           , ZN => n196);
   U73 : INV_X1 port map( A => N156, ZN => n167_port);
   U74 : OAI22_X1 port map( A1 => n143, A2 => n168_port, B1 => n105, B2 => n147
                           , ZN => n193);
   U75 : INV_X1 port map( A => N159, ZN => n168_port);
   U76 : OAI22_X1 port map( A1 => n143, A2 => n166_port, B1 => n101, B2 => n147
                           , ZN => n197);
   U77 : INV_X1 port map( A => N155, ZN => n166_port);
   U78 : NAND4_X1 port map( A1 => n131, A2 => n132, A3 => n75, A4 => n162_port,
                           ZN => n74);
   U79 : INV_X1 port map( A => n76, ZN => n162_port);
   U80 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n130, ZN => n75);
   U81 : AOI21_X1 port map( B1 => n93, B2 => n139, A => n138, ZN => n76);
   U82 : OR3_X1 port map( A1 => IR(29), A2 => IR(31), A3 => n96, ZN => n89);
   U83 : XNOR2_X1 port map( A => n133, B => n236, ZN => n80);
   U84 : NOR3_X1 port map( A1 => n85, A2 => n86, A3 => n87, ZN => n81);
   U85 : INV_X1 port map( A => IR(16), ZN => n236);
   U86 : INV_X1 port map( A => IR(31), ZN => n228);
   U87 : INV_X1 port map( A => IR(29), ZN => n230);
   U88 : INV_X1 port map( A => IR(30), ZN => n229);
   U89 : INV_X1 port map( A => n55, ZN => n164_port);
   U90 : AOI22_X1 port map( A1 => n145, A2 => N184, B1 => n227, B2 => n154_port
                           , ZN => n55);
   U91 : OAI21_X1 port map( B1 => n58, B2 => n227, A => n57, ZN => n54);
   U92 : NOR4_X1 port map( A1 => n64, A2 => n65, A3 => n66, A4 => n67, ZN => 
                           n58);
   U93 : NAND4_X1 port map( A1 => n120, A2 => n119, A3 => n118, A4 => n117, ZN 
                           => n66);
   U94 : NAND4_X1 port map( A1 => n124, A2 => n123, A3 => n122, A4 => n121, ZN 
                           => n67);
   U95 : OAI221_X1 port map( B1 => n154_port, B2 => n165_port, C1 => n100, C2 
                           => n147, A => n52, ZN => n200);
   U96 : INV_X1 port map( A => N154, ZN => n165_port);
   U97 : NAND4_X1 port map( A1 => n98, A2 => n129, A3 => n100, A4 => n68, ZN =>
                           n65);
   U98 : AND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN 
                           => n68);
   U99 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n64);
   U100 : AND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN 
                           => n69);
   U101 : AND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN 
                           => n70);
   U102 : AND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN 
                           => n71);
   U103 : AND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN 
                           => n72);
   U104 : NOR2_X1 port map( A1 => n199, A2 => STALL_CODE_0_port, ZN => 
                           STALL_CODE_1_port);
   U105 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => n202);
   U106 : XNOR2_X1 port map( A => n154_port, B => n98, ZN => n51);
   U107 : INV_X1 port map( A => n73, ZN => n163_port);
   U108 : OAI22_X1 port map( A1 => n133, A2 => n199, B1 => n236, B2 => 
                           EX_STALL_port, ZN => n149);
   U109 : OAI22_X1 port map( A1 => n134, A2 => n199, B1 => n235, B2 => 
                           EX_STALL_port, ZN => n150);
   U110 : OAI22_X1 port map( A1 => n136, A2 => n199, B1 => n234, B2 => 
                           EX_STALL_port, ZN => n151);
   U111 : OAI22_X1 port map( A1 => n137, A2 => n199, B1 => n233, B2 => 
                           EX_STALL_port, ZN => n152);
   U112 : OAI22_X1 port map( A1 => n135, A2 => n199, B1 => n232, B2 => 
                           EX_STALL_port, ZN => n153);
   U113 : OAI22_X1 port map( A1 => n138, A2 => n199, B1 => n238, B2 => 
                           EX_STALL_port, ZN => n155_port);
   U114 : OAI22_X1 port map( A1 => n139, A2 => n199, B1 => n237, B2 => 
                           EX_STALL_port, ZN => n156_port);
   U115 : OAI22_X1 port map( A1 => n131, A2 => n199, B1 => EX_STALL_port, B2 =>
                           n230, ZN => n157_port);
   U116 : OAI22_X1 port map( A1 => n132, A2 => n199, B1 => EX_STALL_port, B2 =>
                           n229, ZN => n158_port);
   U117 : OAI22_X1 port map( A1 => n130, A2 => n199, B1 => EX_STALL_port, B2 =>
                           n228, ZN => n159_port);
   U118 : NAND4_X1 port map( A1 => n88, A2 => n89, A3 => n90, A4 => n91, ZN => 
                           n77);
   U119 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           n78);
   U120 : NOR3_X1 port map( A1 => n83, A2 => IR(27), A3 => n84, ZN => n82);
   U121 : INV_X1 port map( A => IR(27), ZN => n238);
   U122 : INV_X1 port map( A => IR(19), ZN => n233);
   U123 : XNOR2_X1 port map( A => IR(19), B => n137, ZN => n86);
   U124 : INV_X1 port map( A => IR(17), ZN => n235);
   U125 : XNOR2_X1 port map( A => IR(17), B => n134, ZN => n85);
   U126 : XNOR2_X1 port map( A => n134, B => IR(22), ZN => n92);
   U127 : INV_X1 port map( A => IR(20), ZN => n232);
   U128 : XNOR2_X1 port map( A => IR(20), B => n135, ZN => n84);
   U129 : XNOR2_X1 port map( A => n133, B => IR(21), ZN => n94);
   U130 : AOI22_X1 port map( A1 => n237, A2 => IR(27), B1 => n238, B2 => n97, 
                           ZN => n96);
   U131 : OAI22_X1 port map( A1 => n79, A2 => IR(30), B1 => n237, B2 => n231, 
                           ZN => n97);
   U132 : INV_X1 port map( A => IR(18), ZN => n234);
   U133 : XNOR2_X1 port map( A => IR(18), B => n136, ZN => n87);
   U134 : AND4_X1 port map( A1 => IR(3), A2 => IR(2), A3 => IR(1), A4 => IR(26)
                           , ZN => n59);
   U135 : AOI22_X1 port map( A1 => EX_STALL_port, A2 => n93, B1 => IR(26), B2 
                           => n199, ZN => n73);
   U136 : INV_X1 port map( A => IR(26), ZN => n231);
   U137 : NOR4_X1 port map( A1 => IR(28), A2 => IR(27), A3 => IR(10), A4 => 
                           IR(0), ZN => n60);
   U138 : NOR2_X1 port map( A1 => IR(28), A2 => IR(26), ZN => n79);
   U142 : INV_X1 port map( A => IR(28), ZN => n237);
   U143 : NOR3_X1 port map( A1 => n92, A2 => n94, A3 => n95, ZN => n91);
   U144 : XNOR2_X1 port map( A => n135, B => IR(25), ZN => n95);
   U145 : NAND2_X1 port map( A1 => n199, A2 => n74, ZN => IF_STALL_port);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWDU_IR_SIZE32 is

   port( CLOCK, RESET, EN : in std_logic;  IR : in std_logic_vector (31 downto 
         0);  FWD_A, FWD_B : out std_logic_vector (1 downto 0);  FWD_B2 : out 
         std_logic;  ZDU_SEL : out std_logic_vector (1 downto 0));

end FWDU_IR_SIZE32;

architecture SYN_BEHAVIORAL of FWDU_IR_SIZE32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n106, n107, n108, n109, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n173, n175, n2, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n172, n174, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562,
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582 : std_logic;

begin
   
   IR_EX_reg_31_inst : DFFR_X1 port map( D => n175, CK => CLOCK, RN => n200, Q 
                           => n_1556, QN => n2);
   IR_EX_reg_30_inst : DFFR_X1 port map( D => n173, CK => CLOCK, RN => n200, Q 
                           => n193, QN => n174);
   IR_EX_reg_29_inst : DFFR_X1 port map( D => n203, CK => CLOCK, RN => n200, Q 
                           => n189, QN => n177);
   IR_EX_reg_28_inst : DFFR_X1 port map( D => n171, CK => CLOCK, RN => n200, Q 
                           => n190, QN => n123);
   IR_EX_reg_27_inst : DFFR_X1 port map( D => n170, CK => CLOCK, RN => n200, Q 
                           => n_1557, QN => n124);
   IR_EX_reg_26_inst : DFFR_X1 port map( D => n169, CK => CLOCK, RN => n200, Q 
                           => n192, QN => n119);
   IR_EX_reg_20_inst : DFFR_X1 port map( D => n168, CK => CLOCK, RN => n200, Q 
                           => n_1558, QN => n172);
   IR_EX_reg_19_inst : DFFR_X1 port map( D => n167, CK => CLOCK, RN => n200, Q 
                           => n_1559, QN => n134);
   IR_EX_reg_18_inst : DFFR_X1 port map( D => n166, CK => CLOCK, RN => n200, Q 
                           => n_1560, QN => n132);
   IR_EX_reg_17_inst : DFFR_X1 port map( D => n165, CK => CLOCK, RN => n200, Q 
                           => n_1561, QN => n130);
   IR_EX_reg_16_inst : DFFR_X1 port map( D => n164, CK => CLOCK, RN => n200, Q 
                           => n_1562, QN => n131);
   IR_EX_reg_15_inst : DFFR_X1 port map( D => n163, CK => CLOCK, RN => n201, Q 
                           => n_1563, QN => n135);
   IR_EX_reg_14_inst : DFFR_X1 port map( D => n162, CK => CLOCK, RN => n201, Q 
                           => n_1564, QN => n133);
   IR_EX_reg_13_inst : DFFR_X1 port map( D => n161, CK => CLOCK, RN => n201, Q 
                           => n_1565, QN => n129);
   IR_EX_reg_12_inst : DFFR_X1 port map( D => n160, CK => CLOCK, RN => n201, Q 
                           => n_1566, QN => n127);
   IR_EX_reg_11_inst : DFFR_X1 port map( D => n159, CK => CLOCK, RN => n201, Q 
                           => n_1567, QN => n128);
   IR_MEM_reg_31_inst : DFFR_X1 port map( D => n158, CK => CLOCK, RN => n201, Q
                           => n_1568, QN => n120);
   IR_MEM_reg_30_inst : DFFR_X1 port map( D => n157, CK => CLOCK, RN => n201, Q
                           => n_1569, QN => n215);
   IR_MEM_reg_29_inst : DFFR_X1 port map( D => n156, CK => CLOCK, RN => n201, Q
                           => n_1570, QN => n188);
   IR_MEM_reg_28_inst : DFFR_X1 port map( D => n155, CK => CLOCK, RN => n201, Q
                           => n191, QN => n122);
   IR_MEM_reg_27_inst : DFFR_X1 port map( D => n154, CK => CLOCK, RN => n201, Q
                           => n_1571, QN => n121);
   IR_MEM_reg_20_inst : DFFR_X1 port map( D => n153, CK => CLOCK, RN => n201, Q
                           => n_1572, QN => n185);
   IR_MEM_reg_19_inst : DFFR_X1 port map( D => n152, CK => CLOCK, RN => n201, Q
                           => n_1573, QN => n187);
   IR_MEM_reg_18_inst : DFFR_X1 port map( D => n151, CK => CLOCK, RN => n201, Q
                           => n_1574, QN => n183);
   IR_MEM_reg_17_inst : DFFR_X1 port map( D => n150, CK => CLOCK, RN => n200, Q
                           => n_1575, QN => n181);
   IR_MEM_reg_16_inst : DFFR_X1 port map( D => n149, CK => CLOCK, RN => n200, Q
                           => n_1576, QN => n182);
   IR_MEM_reg_15_inst : DFFR_X1 port map( D => n148, CK => CLOCK, RN => n200, Q
                           => n_1577, QN => n184);
   IR_MEM_reg_14_inst : DFFR_X1 port map( D => n147, CK => CLOCK, RN => n200, Q
                           => n_1578, QN => n186);
   IR_MEM_reg_13_inst : DFFR_X1 port map( D => n146, CK => CLOCK, RN => n200, Q
                           => n_1579, QN => n180);
   IR_MEM_reg_12_inst : DFFR_X1 port map( D => n145, CK => CLOCK, RN => n200, Q
                           => n_1580, QN => n178);
   IR_MEM_reg_11_inst : DFFR_X1 port map( D => n144, CK => CLOCK, RN => n200, Q
                           => n_1581, QN => n179);
   FWD_B2_tmp2_reg : DFF_X1 port map( D => n143, CK => CLOCK, Q => n_1582, QN 
                           => n117);
   FWD_B2_reg : DFF_X1 port map( D => n142, CK => CLOCK, Q => FWD_B2, QN => 
                           n118);
   FWD_A_reg_1_inst : DFF_X1 port map( D => n141, CK => CLOCK, Q => FWD_A(1), 
                           QN => n109);
   FWD_A_reg_0_inst : DFF_X1 port map( D => n140, CK => CLOCK, Q => FWD_A(0), 
                           QN => n108);
   FWD_B_reg_1_inst : DFF_X1 port map( D => n139, CK => CLOCK, Q => FWD_B(1), 
                           QN => n107);
   FWD_B_reg_0_inst : DFF_X1 port map( D => n138, CK => CLOCK, Q => FWD_B(0), 
                           QN => n106);
   ZDU_SEL_reg_1_inst : DFF_X1 port map( D => n137, CK => CLOCK, Q => 
                           ZDU_SEL(1), QN => n125);
   ZDU_SEL_reg_0_inst : DFF_X1 port map( D => n136, CK => CLOCK, Q => 
                           ZDU_SEL(0), QN => n126);
   U131 : NAND3_X1 port map( A1 => n206, A2 => n54, A3 => n204, ZN => n53);
   U132 : XOR2_X1 port map( A => n65, B => IR(18), Z => n64);
   U133 : XOR2_X1 port map( A => n66, B => IR(20), Z => n63);
   U134 : NAND3_X1 port map( A1 => n67, A2 => n68, A3 => n69, ZN => n62);
   U135 : XOR2_X1 port map( A => n222, B => n70, Z => n69);
   U136 : XOR2_X1 port map( A => n223, B => n71, Z => n68);
   U137 : XOR2_X1 port map( A => n220, B => n72, Z => n67);
   U138 : NAND3_X1 port map( A1 => n51, A2 => n224, A3 => n73, ZN => n55);
   U139 : NAND3_X1 port map( A1 => n59, A2 => n40, A3 => n74, ZN => n73);
   U140 : XOR2_X1 port map( A => n82, B => IR(17), Z => n81);
   U141 : XOR2_X1 port map( A => n83, B => IR(20), Z => n80);
   U142 : XOR2_X1 port map( A => n223, B => n84, Z => n78);
   U143 : XOR2_X1 port map( A => n220, B => n85, Z => n77);
   U144 : XOR2_X1 port map( A => n221, B => n86, Z => n76);
   U145 : XOR2_X1 port map( A => n66, B => IR(25), Z => n98);
   U146 : XOR2_X1 port map( A => n72, B => IR(24), Z => n97);
   U147 : XOR2_X1 port map( A => n86, B => IR(23), Z => n115);
   U148 : XOR2_X1 port map( A => n82, B => IR(22), Z => n114);
   U149 : XOR2_X1 port map( A => IR(25), B => n207, Z => n112);
   U150 : XOR2_X1 port map( A => IR(24), B => n208, Z => n110);
   U2 : BUF_X1 port map( A => n198, Z => n196);
   U3 : INV_X1 port map( A => n44, ZN => n205);
   U4 : NAND2_X1 port map( A1 => n195, A2 => n200, ZN => n44);
   U5 : INV_X1 port map( A => n196, ZN => n195);
   U6 : BUF_X1 port map( A => n202, Z => n200);
   U7 : BUF_X1 port map( A => n202, Z => n201);
   U8 : INV_X1 port map( A => n197, ZN => n194);
   U9 : BUF_X1 port map( A => n198, Z => n197);
   U10 : INV_X1 port map( A => RESET, ZN => n202);
   U11 : INV_X1 port map( A => n51, ZN => n214);
   U12 : BUF_X1 port map( A => n199, Z => n198);
   U13 : INV_X1 port map( A => EN, ZN => n199);
   U14 : INV_X1 port map( A => n105, ZN => n209);
   U15 : AND4_X1 port map( A1 => n76, A2 => n77, A3 => n78, A4 => n79, ZN => 
                           n40);
   U16 : AND2_X1 port map( A1 => n40, A2 => n61, ZN => n58);
   U17 : INV_X1 port map( A => n50, ZN => n206);
   U18 : INV_X1 port map( A => n83, ZN => n207);
   U19 : INV_X1 port map( A => n85, ZN => n208);
   U20 : INV_X1 port map( A => n96, ZN => n213);
   U21 : INV_X1 port map( A => n72, ZN => n212);
   U22 : INV_X1 port map( A => n54, ZN => n210);
   U23 : OAI211_X1 port map( C1 => n57, C2 => n58, A => n204, B => n59, ZN => 
                           n56);
   U24 : NOR3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n57);
   U25 : OAI211_X1 port map( C1 => n210, C2 => n50, A => n51, B => n52, ZN => 
                           n45);
   U26 : NAND4_X1 port map( A1 => n204, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           n46);
   U27 : NAND4_X1 port map( A1 => n88, A2 => n87, A3 => n50, A4 => n52, ZN => 
                           n93);
   U28 : NAND4_X1 port map( A1 => n95, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           n94);
   U29 : NAND4_X1 port map( A1 => n95, A2 => n206, A3 => n88, A4 => n87, ZN => 
                           n99);
   U30 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n224, A4 => n217, ZN =>
                           n38);
   U31 : INV_X1 port map( A => n32, ZN => n203);
   U32 : OAI22_X1 port map( A1 => n131, A2 => n197, B1 => n182, B2 => EN, ZN =>
                           n149);
   U33 : OAI22_X1 port map( A1 => n129, A2 => n196, B1 => n180, B2 => n194, ZN 
                           => n146);
   U34 : OAI22_X1 port map( A1 => n133, A2 => n196, B1 => n186, B2 => EN, ZN =>
                           n147);
   U35 : OAI22_X1 port map( A1 => n124, A2 => n197, B1 => n121, B2 => n194, ZN 
                           => n154);
   U36 : OAI22_X1 port map( A1 => n123, A2 => n197, B1 => n122, B2 => n194, ZN 
                           => n155);
   U37 : OAI22_X1 port map( A1 => n130, A2 => n197, B1 => n181, B2 => n194, ZN 
                           => n150);
   U38 : OAI22_X1 port map( A1 => n128, A2 => n197, B1 => n179, B2 => EN, ZN =>
                           n144);
   U39 : OAI22_X1 port map( A1 => n132, A2 => n197, B1 => n183, B2 => n194, ZN 
                           => n151);
   U40 : OAI22_X1 port map( A1 => n177, A2 => n197, B1 => n188, B2 => n194, ZN 
                           => n156);
   U41 : OAI22_X1 port map( A1 => n2, A2 => n197, B1 => n120, B2 => n194, ZN =>
                           n158);
   U42 : OAI22_X1 port map( A1 => n135, A2 => n197, B1 => n184, B2 => EN, ZN =>
                           n148);
   U43 : OAI22_X1 port map( A1 => n134, A2 => n197, B1 => n187, B2 => n194, ZN 
                           => n152);
   U44 : OAI22_X1 port map( A1 => n172, A2 => n197, B1 => n185, B2 => n194, ZN 
                           => n153);
   U45 : OAI22_X1 port map( A1 => n174, A2 => n197, B1 => EN, B2 => n215, ZN =>
                           n157);
   U46 : OAI22_X1 port map( A1 => n199, A2 => n223, B1 => n131, B2 => n195, ZN 
                           => n164);
   U47 : OAI22_X1 port map( A1 => n198, A2 => n222, B1 => n130, B2 => n194, ZN 
                           => n165);
   U48 : OAI22_X1 port map( A1 => n198, A2 => n221, B1 => n132, B2 => n194, ZN 
                           => n166);
   U49 : OAI22_X1 port map( A1 => n199, A2 => n219, B1 => n172, B2 => n194, ZN 
                           => n168);
   U50 : OAI22_X1 port map( A1 => n199, A2 => n218, B1 => n119, B2 => n194, ZN 
                           => n169);
   U51 : OAI22_X1 port map( A1 => n199, A2 => n225, B1 => n124, B2 => n194, ZN 
                           => n170);
   U52 : OAI22_X1 port map( A1 => n199, A2 => n224, B1 => n123, B2 => n194, ZN 
                           => n171);
   U53 : OAI22_X1 port map( A1 => n199, A2 => n217, B1 => n174, B2 => n194, ZN 
                           => n173);
   U54 : OAI22_X1 port map( A1 => n199, A2 => n216, B1 => n2, B2 => n195, ZN =>
                           n175);
   U55 : INV_X1 port map( A => IR(31), ZN => n216);
   U56 : OAI21_X1 port map( B1 => n128, B2 => EN, A => n37, ZN => n159);
   U57 : NAND2_X1 port map( A1 => IR(11), A2 => n194, ZN => n37);
   U58 : OAI21_X1 port map( B1 => n129, B2 => EN, A => n35, ZN => n161);
   U59 : NAND2_X1 port map( A1 => IR(13), A2 => n194, ZN => n35);
   U60 : OAI21_X1 port map( B1 => n127, B2 => EN, A => n36, ZN => n160);
   U61 : NAND2_X1 port map( A1 => IR(12), A2 => n194, ZN => n36);
   U62 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n33, ZN => n163);
   U63 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n34, ZN => n162);
   U64 : NAND2_X1 port map( A1 => IR(14), A2 => n194, ZN => n34);
   U65 : OAI22_X1 port map( A1 => n196, A2 => n220, B1 => n134, B2 => n194, ZN 
                           => n167);
   U66 : NAND4_X1 port map( A1 => n123, A2 => n124, A3 => n116, A4 => n174, ZN 
                           => n105);
   U67 : AND2_X1 port map( A1 => n2, A2 => n177, ZN => n116);
   U68 : OAI22_X1 port map( A1 => n127, A2 => n105, B1 => n130, B2 => n209, ZN 
                           => n82);
   U69 : NOR2_X1 port map( A1 => n80, A2 => n81, ZN => n79);
   U70 : OAI22_X1 port map( A1 => n135, A2 => n105, B1 => n172, B2 => n209, ZN 
                           => n83);
   U71 : OAI22_X1 port map( A1 => n129, A2 => n105, B1 => n132, B2 => n209, ZN 
                           => n86);
   U72 : NAND4_X1 port map( A1 => n110, A2 => n111, A3 => n112, A4 => n113, ZN 
                           => n50);
   U73 : NOR2_X1 port map( A1 => n114, A2 => n115, ZN => n113);
   U74 : OAI22_X1 port map( A1 => n133, A2 => n105, B1 => n134, B2 => n209, ZN 
                           => n85);
   U75 : OAI211_X1 port map( C1 => n103, C2 => n104, A => n208, B => n207, ZN 
                           => n88);
   U76 : AND4_X1 port map( A1 => n105, A2 => n132, A3 => n131, A4 => n130, ZN 
                           => n103);
   U77 : AND4_X1 port map( A1 => n209, A2 => n129, A3 => n128, A4 => n127, ZN 
                           => n104);
   U78 : NAND4_X1 port map( A1 => n121, A2 => n215, A3 => n122, A4 => n102, ZN 
                           => n96);
   U79 : AND2_X1 port map( A1 => n188, A2 => n120, ZN => n102);
   U80 : OAI22_X1 port map( A1 => n186, A2 => n96, B1 => n187, B2 => n213, ZN 
                           => n72);
   U81 : OAI211_X1 port map( C1 => n100, C2 => n101, A => n212, B => n211, ZN 
                           => n87);
   U82 : AND4_X1 port map( A1 => n96, A2 => n183, A3 => n182, A4 => n181, ZN =>
                           n100);
   U83 : AND4_X1 port map( A1 => n213, A2 => n180, A3 => n179, A4 => n178, ZN 
                           => n101);
   U84 : INV_X1 port map( A => n66, ZN => n211);
   U85 : OAI22_X1 port map( A1 => n184, A2 => n96, B1 => n185, B2 => n213, ZN 
                           => n66);
   U86 : OAI22_X1 port map( A1 => n128, A2 => n105, B1 => n131, B2 => n209, ZN 
                           => n84);
   U87 : NOR2_X1 port map( A1 => n97, A2 => n98, ZN => n52);
   U88 : OAI22_X1 port map( A1 => n180, A2 => n96, B1 => n183, B2 => n213, ZN 
                           => n65);
   U89 : OAI22_X1 port map( A1 => n179, A2 => n96, B1 => n182, B2 => n213, ZN 
                           => n71);
   U90 : OAI22_X1 port map( A1 => n178, A2 => n96, B1 => n181, B2 => n213, ZN 
                           => n70);
   U91 : XNOR2_X1 port map( A => n65, B => IR(23), ZN => n47);
   U92 : OAI211_X1 port map( C1 => n89, C2 => n90, A => n2, B => n177, ZN => 
                           n54);
   U93 : AND3_X1 port map( A1 => n124, A2 => n190, A3 => n174, ZN => n89);
   U94 : NOR2_X1 port map( A1 => n124, A2 => n190, ZN => n90);
   U95 : INV_X1 port map( A => IR(16), ZN => n223);
   U96 : OAI211_X1 port map( C1 => n91, C2 => n92, A => n188, B => n120, ZN => 
                           n51);
   U97 : AND3_X1 port map( A1 => n121, A2 => n191, A3 => n215, ZN => n91);
   U98 : NOR2_X1 port map( A1 => n121, A2 => n191, ZN => n92);
   U99 : NOR4_X1 port map( A1 => n193, A2 => n189, A3 => n75, A4 => n2, ZN => 
                           n61);
   U100 : AOI22_X1 port map( A1 => n192, A2 => n123, B1 => n124, B2 => n119, ZN
                           => n75);
   U101 : NAND4_X1 port map( A1 => n220, A2 => n219, A3 => n221, A4 => n43, ZN 
                           => n42);
   U102 : INV_X1 port map( A => IR(30), ZN => n217);
   U103 : OAI22_X1 port map( A1 => n127, A2 => n197, B1 => n178, B2 => EN, ZN 
                           => n145);
   U104 : INV_X1 port map( A => IR(27), ZN => n225);
   U105 : NAND2_X1 port map( A1 => IR(27), A2 => n218, ZN => n41);
   U106 : NOR4_X1 port map( A1 => IR(27), A2 => IR(29), A3 => IR(30), A4 => 
                           IR(31), ZN => n59);
   U107 : INV_X1 port map( A => IR(19), ZN => n220);
   U108 : NOR2_X1 port map( A1 => IR(17), A2 => IR(16), ZN => n43);
   U109 : INV_X1 port map( A => IR(17), ZN => n222);
   U110 : XNOR2_X1 port map( A => n70, B => IR(22), ZN => n48);
   U111 : AOI22_X1 port map( A1 => n194, A2 => IR(29), B1 => n189, B2 => n197, 
                           ZN => n32);
   U112 : INV_X1 port map( A => IR(20), ZN => n219);
   U113 : XNOR2_X1 port map( A => n71, B => IR(21), ZN => n49);
   U114 : XNOR2_X1 port map( A => IR(21), B => n84, ZN => n111);
   U115 : INV_X1 port map( A => IR(18), ZN => n221);
   U116 : INV_X1 port map( A => IR(26), ZN => n218);
   U117 : INV_X1 port map( A => IR(28), ZN => n224);
   U118 : AOI211_X1 port map( C1 => n61, C2 => n218, A => IR(28), B => n210, ZN
                           => n74);
   U119 : OAI21_X1 port map( B1 => n108, B2 => n205, A => n53, ZN => n140);
   U120 : OAI21_X1 port map( B1 => n126, B2 => n205, A => n99, ZN => n136);
   U121 : OAI22_X1 port map( A1 => n117, A2 => n205, B1 => n38, B2 => n39, ZN 
                           => n143);
   U122 : OAI22_X1 port map( A1 => n107, A2 => n205, B1 => n55, B2 => n56, ZN 
                           => n139);
   U123 : OAI22_X1 port map( A1 => n125, A2 => n205, B1 => n93, B2 => n94, ZN 
                           => n137);
   U124 : OAI22_X1 port map( A1 => n106, A2 => n205, B1 => n60, B2 => n73, ZN 
                           => n138);
   U125 : OAI22_X1 port map( A1 => n117, A2 => n44, B1 => n118, B2 => n205, ZN 
                           => n142);
   U126 : OAI22_X1 port map( A1 => n45, A2 => n46, B1 => n109, B2 => n205, ZN 
                           => n141);
   U127 : NAND4_X1 port map( A1 => n205, A2 => n40, A3 => IR(29), A4 => IR(31),
                           ZN => n39);
   U128 : INV_X1 port map( A => n60, ZN => n204);
   U129 : AND3_X1 port map( A1 => n205, A2 => IR(28), A3 => n59, ZN => n95);
   U130 : OAI221_X1 port map( B1 => n214, B2 => n87, C1 => n210, C2 => n88, A 
                           => n205, ZN => n60);
   U151 : NAND2_X1 port map( A1 => IR(15), A2 => n194, ZN => n33);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( CLOCK : in std_logic;  AluOpcode : in std_logic_vector (0 to 4);  A, B
         : in std_logic_vector (31 downto 0);  Cin : in std_logic;  ALU_out : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic;  COND : out
         std_logic_vector (5 downto 0));

end ALU_NBIT32;

architecture SYN_BEHAVIORAL of ALU_NBIT32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX4to1_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUL
      port( CLOCK : in std_logic;  A, B : in std_logic_vector (15 downto 0);  Y
            : out std_logic_vector (31 downto 0));
   end component;
   
   component CMP_NBIT32
      port( SUM : in std_logic_vector (31 downto 0);  Cout : in std_logic;  
            A_L_B, A_LE_B, A_G_B, A_GE_B, A_E_B, A_NE_B : out std_logic);
   end component;
   
   component LOGIC_NBIT32_N_SELECTOR4
      port( S : in std_logic_vector (3 downto 0);  A, B : in std_logic_vector 
            (31 downto 0);  O : out std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER
      port( data_in : in std_logic_vector (31 downto 0);  R : in 
            std_logic_vector (4 downto 0);  conf : in std_logic_vector (1 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component AND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal Cout_port, cin_internal, en_adder, A_adder_31_port, A_adder_30_port, 
      A_adder_29_port, A_adder_28_port, A_adder_27_port, A_adder_26_port, 
      A_adder_25_port, A_adder_24_port, A_adder_23_port, A_adder_22_port, 
      A_adder_21_port, A_adder_20_port, A_adder_19_port, A_adder_18_port, 
      A_adder_17_port, A_adder_16_port, A_adder_15_port, A_adder_14_port, 
      A_adder_13_port, A_adder_12_port, A_adder_11_port, A_adder_10_port, 
      A_adder_9_port, A_adder_8_port, A_adder_7_port, A_adder_6_port, 
      A_adder_5_port, A_adder_4_port, A_adder_3_port, A_adder_2_port, 
      A_adder_1_port, A_adder_0_port, B_adder_31_port, B_adder_30_port, 
      B_adder_29_port, B_adder_28_port, B_adder_27_port, B_adder_26_port, 
      B_adder_25_port, B_adder_24_port, B_adder_23_port, B_adder_22_port, 
      B_adder_21_port, B_adder_20_port, B_adder_19_port, B_adder_18_port, 
      B_adder_17_port, B_adder_16_port, B_adder_15_port, B_adder_14_port, 
      B_adder_13_port, B_adder_12_port, B_adder_11_port, B_adder_10_port, 
      B_adder_9_port, B_adder_8_port, B_adder_7_port, B_adder_6_port, 
      B_adder_5_port, B_adder_4_port, B_adder_3_port, B_adder_2_port, 
      B_adder_1_port, B_adder_0_port, en_logic, A_logic_31_port, 
      A_logic_30_port, A_logic_29_port, A_logic_28_port, A_logic_27_port, 
      A_logic_26_port, A_logic_25_port, A_logic_24_port, A_logic_23_port, 
      A_logic_22_port, A_logic_21_port, A_logic_20_port, A_logic_19_port, 
      A_logic_18_port, A_logic_17_port, A_logic_16_port, A_logic_15_port, 
      A_logic_14_port, A_logic_13_port, A_logic_12_port, A_logic_11_port, 
      A_logic_10_port, A_logic_9_port, A_logic_8_port, A_logic_7_port, 
      A_logic_6_port, A_logic_5_port, A_logic_4_port, A_logic_3_port, 
      A_logic_2_port, A_logic_1_port, A_logic_0_port, B_logic_31_port, 
      B_logic_30_port, B_logic_29_port, B_logic_28_port, B_logic_27_port, 
      B_logic_26_port, B_logic_25_port, B_logic_24_port, B_logic_23_port, 
      B_logic_22_port, B_logic_21_port, B_logic_20_port, B_logic_19_port, 
      B_logic_18_port, B_logic_17_port, B_logic_16_port, B_logic_15_port, 
      B_logic_14_port, B_logic_13_port, B_logic_12_port, B_logic_11_port, 
      B_logic_10_port, B_logic_9_port, B_logic_8_port, B_logic_7_port, 
      B_logic_6_port, B_logic_5_port, B_logic_4_port, B_logic_3_port, 
      B_logic_2_port, B_logic_1_port, B_logic_0_port, en_shifter, 
      A_shifter_31_port, A_shifter_30_port, A_shifter_29_port, 
      A_shifter_28_port, A_shifter_27_port, A_shifter_26_port, 
      A_shifter_25_port, A_shifter_24_port, A_shifter_23_port, 
      A_shifter_22_port, A_shifter_21_port, A_shifter_20_port, 
      A_shifter_19_port, A_shifter_18_port, A_shifter_17_port, 
      A_shifter_16_port, A_shifter_15_port, A_shifter_14_port, 
      A_shifter_13_port, A_shifter_12_port, A_shifter_11_port, 
      A_shifter_10_port, A_shifter_9_port, A_shifter_8_port, A_shifter_7_port, 
      A_shifter_6_port, A_shifter_5_port, A_shifter_4_port, A_shifter_3_port, 
      A_shifter_2_port, A_shifter_1_port, A_shifter_0_port, B_shifter_4_port, 
      B_shifter_3_port, B_shifter_2_port, B_shifter_1_port, B_shifter_0_port, 
      in_cmp_31_port, in_cmp_30_port, in_cmp_29_port, in_cmp_28_port, 
      in_cmp_27_port, in_cmp_26_port, in_cmp_25_port, in_cmp_24_port, 
      in_cmp_23_port, in_cmp_22_port, in_cmp_21_port, in_cmp_20_port, 
      in_cmp_19_port, in_cmp_18_port, in_cmp_17_port, in_cmp_16_port, 
      in_cmp_15_port, in_cmp_14_port, in_cmp_13_port, in_cmp_12_port, 
      in_cmp_11_port, in_cmp_10_port, in_cmp_9_port, in_cmp_8_port, 
      in_cmp_7_port, in_cmp_6_port, in_cmp_5_port, in_cmp_4_port, in_cmp_3_port
      , in_cmp_2_port, in_cmp_1_port, in_cmp_0_port, out_adder_31_port, 
      out_adder_30_port, out_adder_29_port, out_adder_28_port, 
      out_adder_27_port, out_adder_26_port, out_adder_25_port, 
      out_adder_24_port, out_adder_23_port, out_adder_22_port, 
      out_adder_21_port, out_adder_20_port, out_adder_19_port, 
      out_adder_18_port, out_adder_17_port, out_adder_16_port, 
      out_adder_15_port, out_adder_14_port, out_adder_13_port, 
      out_adder_12_port, out_adder_11_port, out_adder_10_port, out_adder_9_port
      , out_adder_8_port, out_adder_7_port, out_adder_6_port, out_adder_5_port,
      out_adder_4_port, out_adder_3_port, out_adder_2_port, out_adder_1_port, 
      out_adder_0_port, A_mul_15_port, A_mul_14_port, A_mul_13_port, 
      A_mul_12_port, A_mul_11_port, A_mul_10_port, A_mul_9_port, A_mul_8_port, 
      A_mul_7_port, A_mul_6_port, A_mul_5_port, A_mul_4_port, A_mul_3_port, 
      A_mul_2_port, A_mul_1_port, A_mul_0_port, B_mul_15_port, B_mul_14_port, 
      B_mul_13_port, B_mul_12_port, B_mul_11_port, B_mul_10_port, B_mul_9_port,
      B_mul_8_port, B_mul_7_port, B_mul_6_port, B_mul_5_port, B_mul_4_port, 
      B_mul_3_port, B_mul_2_port, B_mul_1_port, B_mul_0_port, conf_1_port, 
      conf_0_port, out_shifter_31_port, out_shifter_30_port, 
      out_shifter_29_port, out_shifter_28_port, out_shifter_27_port, 
      out_shifter_26_port, out_shifter_25_port, out_shifter_24_port, 
      out_shifter_23_port, out_shifter_22_port, out_shifter_21_port, 
      out_shifter_20_port, out_shifter_19_port, out_shifter_18_port, 
      out_shifter_17_port, out_shifter_16_port, out_shifter_15_port, 
      out_shifter_14_port, out_shifter_13_port, out_shifter_12_port, 
      out_shifter_11_port, out_shifter_10_port, out_shifter_9_port, 
      out_shifter_8_port, out_shifter_7_port, out_shifter_6_port, 
      out_shifter_5_port, out_shifter_4_port, out_shifter_3_port, 
      out_shifter_2_port, out_shifter_1_port, out_shifter_0_port, 
      logic_sel_3_port, logic_sel_2_port, logic_sel_1_port, logic_sel_0_port, 
      out_logic_31_port, out_logic_30_port, out_logic_29_port, 
      out_logic_28_port, out_logic_27_port, out_logic_26_port, 
      out_logic_25_port, out_logic_24_port, out_logic_23_port, 
      out_logic_22_port, out_logic_21_port, out_logic_20_port, 
      out_logic_19_port, out_logic_18_port, out_logic_17_port, 
      out_logic_16_port, out_logic_15_port, out_logic_14_port, 
      out_logic_13_port, out_logic_12_port, out_logic_11_port, 
      out_logic_10_port, out_logic_9_port, out_logic_8_port, out_logic_7_port, 
      out_logic_6_port, out_logic_5_port, out_logic_4_port, out_logic_3_port, 
      out_logic_2_port, out_logic_1_port, out_logic_0_port, out_mul_31_port, 
      out_mul_30_port, out_mul_29_port, out_mul_28_port, out_mul_27_port, 
      out_mul_26_port, out_mul_25_port, out_mul_24_port, out_mul_23_port, 
      out_mul_22_port, out_mul_21_port, out_mul_20_port, out_mul_19_port, 
      out_mul_18_port, out_mul_17_port, out_mul_16_port, out_mul_15_port, 
      out_mul_14_port, out_mul_13_port, out_mul_12_port, out_mul_11_port, 
      out_mul_10_port, out_mul_9_port, out_mul_8_port, out_mul_7_port, 
      out_mul_6_port, out_mul_5_port, out_mul_4_port, out_mul_3_port, 
      out_mul_2_port, out_mul_1_port, out_mul_0_port, mux_out_1_port, 
      mux_out_0_port, N88, N89, N90, N91, N92, N93, n1, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88_port, 
      n89_port, n90_port, n91_port, n92_port, n93_port, n94, n95, n96, n97 : 
      std_logic;

begin
   Cout <= Cout_port;
   
   conf_reg_1_inst : DLH_X1 port map( G => N91, D => N93, Q => conf_1_port);
   conf_reg_0_inst : DLH_X1 port map( G => N91, D => N92, Q => conf_0_port);
   logic_sel_reg_3_inst : DLH_X1 port map( G => n78, D => N90, Q => 
                           logic_sel_3_port);
   logic_sel_reg_2_inst : DLH_X1 port map( G => n78, D => N89, Q => 
                           logic_sel_2_port);
   logic_sel_reg_1_inst : DLH_X1 port map( G => n78, D => N89, Q => 
                           logic_sel_1_port);
   logic_sel_reg_0_inst : DLH_X1 port map( G => n78, D => N88, Q => 
                           logic_sel_0_port);
   U39 : NAND3_X1 port map( A1 => n19, A2 => n93_port, A3 => n20, ZN => n16);
   U40 : NAND3_X1 port map( A1 => n17, A2 => AluOpcode(1), A3 => AluOpcode(4), 
                           ZN => n26);
   U41 : NAND3_X1 port map( A1 => n97, A2 => n93_port, A3 => AluOpcode(2), ZN 
                           => n12);
   ADDER_A_i_0 : AND2_0 port map( A => A(0), B => n87, Y => A_adder_0_port);
   ADDER_B_i_0 : AND2_228 port map( A => B(0), B => n82, Y => B_adder_0_port);
   ADDER_A_i_1 : AND2_227 port map( A => A(1), B => n82, Y => A_adder_1_port);
   ADDER_B_i_1 : AND2_226 port map( A => B(1), B => n82, Y => B_adder_1_port);
   ADDER_A_i_2 : AND2_225 port map( A => A(2), B => n82, Y => A_adder_2_port);
   ADDER_B_i_2 : AND2_224 port map( A => B(2), B => n82, Y => B_adder_2_port);
   ADDER_A_i_3 : AND2_223 port map( A => A(3), B => n82, Y => A_adder_3_port);
   ADDER_B_i_3 : AND2_222 port map( A => B(3), B => n82, Y => B_adder_3_port);
   ADDER_A_i_4 : AND2_221 port map( A => A(4), B => n82, Y => A_adder_4_port);
   ADDER_B_i_4 : AND2_220 port map( A => B(4), B => n82, Y => B_adder_4_port);
   ADDER_A_i_5 : AND2_219 port map( A => A(5), B => n82, Y => A_adder_5_port);
   ADDER_B_i_5 : AND2_218 port map( A => B(5), B => n82, Y => B_adder_5_port);
   ADDER_A_i_6 : AND2_217 port map( A => A(6), B => n82, Y => A_adder_6_port);
   ADDER_B_i_6 : AND2_216 port map( A => B(6), B => n83, Y => B_adder_6_port);
   ADDER_A_i_7 : AND2_215 port map( A => A(7), B => n83, Y => A_adder_7_port);
   ADDER_B_i_7 : AND2_214 port map( A => B(7), B => n83, Y => B_adder_7_port);
   ADDER_A_i_8 : AND2_213 port map( A => A(8), B => n83, Y => A_adder_8_port);
   ADDER_B_i_8 : AND2_212 port map( A => B(8), B => n83, Y => B_adder_8_port);
   ADDER_A_i_9 : AND2_211 port map( A => A(9), B => n83, Y => A_adder_9_port);
   ADDER_B_i_9 : AND2_210 port map( A => B(9), B => n83, Y => B_adder_9_port);
   ADDER_A_i_10 : AND2_209 port map( A => A(10), B => n83, Y => A_adder_10_port
                           );
   ADDER_B_i_10 : AND2_208 port map( A => B(10), B => n83, Y => B_adder_10_port
                           );
   ADDER_A_i_11 : AND2_207 port map( A => A(11), B => n83, Y => A_adder_11_port
                           );
   ADDER_B_i_11 : AND2_206 port map( A => B(11), B => n83, Y => B_adder_11_port
                           );
   ADDER_A_i_12 : AND2_205 port map( A => A(12), B => n83, Y => A_adder_12_port
                           );
   ADDER_B_i_12 : AND2_204 port map( A => B(12), B => n84, Y => B_adder_12_port
                           );
   ADDER_A_i_13 : AND2_203 port map( A => A(13), B => n84, Y => A_adder_13_port
                           );
   ADDER_B_i_13 : AND2_202 port map( A => B(13), B => n84, Y => B_adder_13_port
                           );
   ADDER_A_i_14 : AND2_201 port map( A => A(14), B => n84, Y => A_adder_14_port
                           );
   ADDER_B_i_14 : AND2_200 port map( A => B(14), B => n84, Y => B_adder_14_port
                           );
   ADDER_A_i_15 : AND2_199 port map( A => A(15), B => n84, Y => A_adder_15_port
                           );
   ADDER_B_i_15 : AND2_198 port map( A => B(15), B => n84, Y => B_adder_15_port
                           );
   ADDER_A_i_16 : AND2_197 port map( A => A(16), B => n84, Y => A_adder_16_port
                           );
   ADDER_B_i_16 : AND2_196 port map( A => B(16), B => n84, Y => B_adder_16_port
                           );
   ADDER_A_i_17 : AND2_195 port map( A => A(17), B => n84, Y => A_adder_17_port
                           );
   ADDER_B_i_17 : AND2_194 port map( A => B(17), B => n84, Y => B_adder_17_port
                           );
   ADDER_A_i_18 : AND2_193 port map( A => A(18), B => n84, Y => A_adder_18_port
                           );
   ADDER_B_i_18 : AND2_192 port map( A => B(18), B => n85, Y => B_adder_18_port
                           );
   ADDER_A_i_19 : AND2_191 port map( A => A(19), B => n85, Y => A_adder_19_port
                           );
   ADDER_B_i_19 : AND2_190 port map( A => B(19), B => n85, Y => B_adder_19_port
                           );
   ADDER_A_i_20 : AND2_189 port map( A => A(20), B => n85, Y => A_adder_20_port
                           );
   ADDER_B_i_20 : AND2_188 port map( A => B(20), B => n85, Y => B_adder_20_port
                           );
   ADDER_A_i_21 : AND2_187 port map( A => A(21), B => n85, Y => A_adder_21_port
                           );
   ADDER_B_i_21 : AND2_186 port map( A => B(21), B => n85, Y => B_adder_21_port
                           );
   ADDER_A_i_22 : AND2_185 port map( A => A(22), B => n85, Y => A_adder_22_port
                           );
   ADDER_B_i_22 : AND2_184 port map( A => B(22), B => n85, Y => B_adder_22_port
                           );
   ADDER_A_i_23 : AND2_183 port map( A => A(23), B => n85, Y => A_adder_23_port
                           );
   ADDER_B_i_23 : AND2_182 port map( A => B(23), B => n85, Y => B_adder_23_port
                           );
   ADDER_A_i_24 : AND2_181 port map( A => A(24), B => n85, Y => A_adder_24_port
                           );
   ADDER_B_i_24 : AND2_180 port map( A => B(24), B => n86, Y => B_adder_24_port
                           );
   ADDER_A_i_25 : AND2_179 port map( A => A(25), B => n86, Y => A_adder_25_port
                           );
   ADDER_B_i_25 : AND2_178 port map( A => B(25), B => n86, Y => B_adder_25_port
                           );
   ADDER_A_i_26 : AND2_177 port map( A => A(26), B => n86, Y => A_adder_26_port
                           );
   ADDER_B_i_26 : AND2_176 port map( A => B(26), B => n86, Y => B_adder_26_port
                           );
   ADDER_A_i_27 : AND2_175 port map( A => A(27), B => n86, Y => A_adder_27_port
                           );
   ADDER_B_i_27 : AND2_174 port map( A => B(27), B => n86, Y => B_adder_27_port
                           );
   ADDER_A_i_28 : AND2_173 port map( A => A(28), B => n86, Y => A_adder_28_port
                           );
   ADDER_B_i_28 : AND2_172 port map( A => B(28), B => n86, Y => B_adder_28_port
                           );
   ADDER_A_i_29 : AND2_171 port map( A => A(29), B => n86, Y => A_adder_29_port
                           );
   ADDER_B_i_29 : AND2_170 port map( A => B(29), B => n86, Y => B_adder_29_port
                           );
   ADDER_A_i_30 : AND2_169 port map( A => A(30), B => n86, Y => A_adder_30_port
                           );
   ADDER_B_i_30 : AND2_168 port map( A => B(30), B => n87, Y => B_adder_30_port
                           );
   ADDER_A_i_31 : AND2_167 port map( A => A(31), B => n87, Y => A_adder_31_port
                           );
   ADDER_B_i_31 : AND2_166 port map( A => B(31), B => n87, Y => B_adder_31_port
                           );
   LOGIC_A_i_0 : AND2_165 port map( A => A(0), B => n73, Y => A_logic_0_port);
   LOGIC_B_i_0 : AND2_164 port map( A => B(0), B => n73, Y => B_logic_0_port);
   LOGIC_A_i_1 : AND2_163 port map( A => A(1), B => n73, Y => A_logic_1_port);
   LOGIC_B_i_1 : AND2_162 port map( A => B(1), B => n73, Y => B_logic_1_port);
   LOGIC_A_i_2 : AND2_161 port map( A => A(2), B => n73, Y => A_logic_2_port);
   LOGIC_B_i_2 : AND2_160 port map( A => B(2), B => n73, Y => B_logic_2_port);
   LOGIC_A_i_3 : AND2_159 port map( A => A(3), B => n73, Y => A_logic_3_port);
   LOGIC_B_i_3 : AND2_158 port map( A => B(3), B => n73, Y => B_logic_3_port);
   LOGIC_A_i_4 : AND2_157 port map( A => A(4), B => n73, Y => A_logic_4_port);
   LOGIC_B_i_4 : AND2_156 port map( A => B(4), B => n73, Y => B_logic_4_port);
   LOGIC_A_i_5 : AND2_155 port map( A => A(5), B => n73, Y => A_logic_5_port);
   LOGIC_B_i_5 : AND2_154 port map( A => B(5), B => n73, Y => B_logic_5_port);
   LOGIC_A_i_6 : AND2_153 port map( A => A(6), B => n74, Y => A_logic_6_port);
   LOGIC_B_i_6 : AND2_152 port map( A => B(6), B => n74, Y => B_logic_6_port);
   LOGIC_A_i_7 : AND2_151 port map( A => A(7), B => n74, Y => A_logic_7_port);
   LOGIC_B_i_7 : AND2_150 port map( A => B(7), B => n74, Y => B_logic_7_port);
   LOGIC_A_i_8 : AND2_149 port map( A => A(8), B => n74, Y => A_logic_8_port);
   LOGIC_B_i_8 : AND2_148 port map( A => B(8), B => n74, Y => B_logic_8_port);
   LOGIC_A_i_9 : AND2_147 port map( A => A(9), B => n74, Y => A_logic_9_port);
   LOGIC_B_i_9 : AND2_146 port map( A => B(9), B => n74, Y => B_logic_9_port);
   LOGIC_A_i_10 : AND2_145 port map( A => A(10), B => n74, Y => A_logic_10_port
                           );
   LOGIC_B_i_10 : AND2_144 port map( A => B(10), B => n74, Y => B_logic_10_port
                           );
   LOGIC_A_i_11 : AND2_143 port map( A => A(11), B => n74, Y => A_logic_11_port
                           );
   LOGIC_B_i_11 : AND2_142 port map( A => B(11), B => n74, Y => B_logic_11_port
                           );
   LOGIC_A_i_12 : AND2_141 port map( A => A(12), B => n75, Y => A_logic_12_port
                           );
   LOGIC_B_i_12 : AND2_140 port map( A => B(12), B => n75, Y => B_logic_12_port
                           );
   LOGIC_A_i_13 : AND2_139 port map( A => A(13), B => n75, Y => A_logic_13_port
                           );
   LOGIC_B_i_13 : AND2_138 port map( A => B(13), B => n75, Y => B_logic_13_port
                           );
   LOGIC_A_i_14 : AND2_137 port map( A => A(14), B => n75, Y => A_logic_14_port
                           );
   LOGIC_B_i_14 : AND2_136 port map( A => B(14), B => n75, Y => B_logic_14_port
                           );
   LOGIC_A_i_15 : AND2_135 port map( A => A(15), B => n75, Y => A_logic_15_port
                           );
   LOGIC_B_i_15 : AND2_134 port map( A => B(15), B => n75, Y => B_logic_15_port
                           );
   LOGIC_A_i_16 : AND2_133 port map( A => A(16), B => n75, Y => A_logic_16_port
                           );
   LOGIC_B_i_16 : AND2_132 port map( A => B(16), B => n75, Y => B_logic_16_port
                           );
   LOGIC_A_i_17 : AND2_131 port map( A => A(17), B => n75, Y => A_logic_17_port
                           );
   LOGIC_B_i_17 : AND2_130 port map( A => B(17), B => n75, Y => B_logic_17_port
                           );
   LOGIC_A_i_18 : AND2_129 port map( A => A(18), B => n76, Y => A_logic_18_port
                           );
   LOGIC_B_i_18 : AND2_128 port map( A => B(18), B => n76, Y => B_logic_18_port
                           );
   LOGIC_A_i_19 : AND2_127 port map( A => A(19), B => n76, Y => A_logic_19_port
                           );
   LOGIC_B_i_19 : AND2_126 port map( A => B(19), B => n76, Y => B_logic_19_port
                           );
   LOGIC_A_i_20 : AND2_125 port map( A => A(20), B => n76, Y => A_logic_20_port
                           );
   LOGIC_B_i_20 : AND2_124 port map( A => B(20), B => n76, Y => B_logic_20_port
                           );
   LOGIC_A_i_21 : AND2_123 port map( A => A(21), B => n76, Y => A_logic_21_port
                           );
   LOGIC_B_i_21 : AND2_122 port map( A => B(21), B => n76, Y => B_logic_21_port
                           );
   LOGIC_A_i_22 : AND2_121 port map( A => A(22), B => n76, Y => A_logic_22_port
                           );
   LOGIC_B_i_22 : AND2_120 port map( A => B(22), B => n76, Y => B_logic_22_port
                           );
   LOGIC_A_i_23 : AND2_119 port map( A => A(23), B => n76, Y => A_logic_23_port
                           );
   LOGIC_B_i_23 : AND2_118 port map( A => B(23), B => n76, Y => B_logic_23_port
                           );
   LOGIC_A_i_24 : AND2_117 port map( A => A(24), B => n77, Y => A_logic_24_port
                           );
   LOGIC_B_i_24 : AND2_116 port map( A => B(24), B => n77, Y => B_logic_24_port
                           );
   LOGIC_A_i_25 : AND2_115 port map( A => A(25), B => n77, Y => A_logic_25_port
                           );
   LOGIC_B_i_25 : AND2_114 port map( A => B(25), B => n77, Y => B_logic_25_port
                           );
   LOGIC_A_i_26 : AND2_113 port map( A => A(26), B => n77, Y => A_logic_26_port
                           );
   LOGIC_B_i_26 : AND2_112 port map( A => B(26), B => n77, Y => B_logic_26_port
                           );
   LOGIC_A_i_27 : AND2_111 port map( A => A(27), B => n77, Y => A_logic_27_port
                           );
   LOGIC_B_i_27 : AND2_110 port map( A => B(27), B => n77, Y => B_logic_27_port
                           );
   LOGIC_A_i_28 : AND2_109 port map( A => A(28), B => n77, Y => A_logic_28_port
                           );
   LOGIC_B_i_28 : AND2_108 port map( A => B(28), B => n77, Y => B_logic_28_port
                           );
   LOGIC_A_i_29 : AND2_107 port map( A => A(29), B => n77, Y => A_logic_29_port
                           );
   LOGIC_B_i_29 : AND2_106 port map( A => B(29), B => n77, Y => B_logic_29_port
                           );
   LOGIC_A_i_30 : AND2_105 port map( A => A(30), B => n78, Y => A_logic_30_port
                           );
   LOGIC_B_i_30 : AND2_104 port map( A => B(30), B => n78, Y => B_logic_30_port
                           );
   LOGIC_A_i_31 : AND2_103 port map( A => A(31), B => n78, Y => A_logic_31_port
                           );
   LOGIC_B_i_31 : AND2_102 port map( A => B(31), B => n78, Y => B_logic_31_port
                           );
   SHIFTER_A_i_0 : AND2_101 port map( A => A(0), B => n66, Y => 
                           A_shifter_0_port);
   SHIFTER_A_i_1 : AND2_100 port map( A => A(1), B => n66, Y => 
                           A_shifter_1_port);
   SHIFTER_A_i_2 : AND2_99 port map( A => A(2), B => n66, Y => A_shifter_2_port
                           );
   SHIFTER_A_i_3 : AND2_98 port map( A => A(3), B => n66, Y => A_shifter_3_port
                           );
   SHIFTER_A_i_4 : AND2_97 port map( A => A(4), B => n66, Y => A_shifter_4_port
                           );
   SHIFTER_A_i_5 : AND2_96 port map( A => A(5), B => n66, Y => A_shifter_5_port
                           );
   SHIFTER_A_i_6 : AND2_95 port map( A => A(6), B => n66, Y => A_shifter_6_port
                           );
   SHIFTER_A_i_7 : AND2_94 port map( A => A(7), B => n66, Y => A_shifter_7_port
                           );
   SHIFTER_A_i_8 : AND2_93 port map( A => A(8), B => n66, Y => A_shifter_8_port
                           );
   SHIFTER_A_i_9 : AND2_92 port map( A => A(9), B => n66, Y => A_shifter_9_port
                           );
   SHIFTER_A_i_10 : AND2_91 port map( A => A(10), B => n66, Y => 
                           A_shifter_10_port);
   SHIFTER_A_i_11 : AND2_90 port map( A => A(11), B => n66, Y => 
                           A_shifter_11_port);
   SHIFTER_A_i_12 : AND2_89 port map( A => A(12), B => n67, Y => 
                           A_shifter_12_port);
   SHIFTER_A_i_13 : AND2_88 port map( A => A(13), B => n67, Y => 
                           A_shifter_13_port);
   SHIFTER_A_i_14 : AND2_87 port map( A => A(14), B => n67, Y => 
                           A_shifter_14_port);
   SHIFTER_A_i_15 : AND2_86 port map( A => A(15), B => n67, Y => 
                           A_shifter_15_port);
   SHIFTER_A_i_16 : AND2_85 port map( A => A(16), B => n67, Y => 
                           A_shifter_16_port);
   SHIFTER_A_i_17 : AND2_84 port map( A => A(17), B => n67, Y => 
                           A_shifter_17_port);
   SHIFTER_A_i_18 : AND2_83 port map( A => A(18), B => n67, Y => 
                           A_shifter_18_port);
   SHIFTER_A_i_19 : AND2_82 port map( A => A(19), B => n67, Y => 
                           A_shifter_19_port);
   SHIFTER_A_i_20 : AND2_81 port map( A => A(20), B => n67, Y => 
                           A_shifter_20_port);
   SHIFTER_A_i_21 : AND2_80 port map( A => A(21), B => n67, Y => 
                           A_shifter_21_port);
   SHIFTER_A_i_22 : AND2_79 port map( A => A(22), B => n67, Y => 
                           A_shifter_22_port);
   SHIFTER_A_i_23 : AND2_78 port map( A => A(23), B => n67, Y => 
                           A_shifter_23_port);
   SHIFTER_A_i_24 : AND2_77 port map( A => A(24), B => n68, Y => 
                           A_shifter_24_port);
   SHIFTER_A_i_25 : AND2_76 port map( A => A(25), B => n68, Y => 
                           A_shifter_25_port);
   SHIFTER_A_i_26 : AND2_75 port map( A => A(26), B => n68, Y => 
                           A_shifter_26_port);
   SHIFTER_A_i_27 : AND2_74 port map( A => A(27), B => n68, Y => 
                           A_shifter_27_port);
   SHIFTER_A_i_28 : AND2_73 port map( A => A(28), B => n68, Y => 
                           A_shifter_28_port);
   SHIFTER_A_i_29 : AND2_72 port map( A => A(29), B => n68, Y => 
                           A_shifter_29_port);
   SHIFTER_A_i_30 : AND2_71 port map( A => A(30), B => n68, Y => 
                           A_shifter_30_port);
   SHIFTER_A_i_31 : AND2_70 port map( A => A(31), B => n68, Y => 
                           A_shifter_31_port);
   SHIFTER_B_i_0 : AND2_69 port map( A => B(0), B => n68, Y => B_shifter_0_port
                           );
   SHIFTER_B_i_1 : AND2_68 port map( A => B(1), B => n68, Y => B_shifter_1_port
                           );
   SHIFTER_B_i_2 : AND2_67 port map( A => B(2), B => n68, Y => B_shifter_2_port
                           );
   SHIFTER_B_i_3 : AND2_66 port map( A => B(3), B => n68, Y => B_shifter_3_port
                           );
   SHIFTER_B_i_4 : AND2_65 port map( A => B(4), B => n69, Y => B_shifter_4_port
                           );
   SUM_i_0 : AND2_64 port map( A => out_adder_0_port, B => n61, Y => 
                           in_cmp_0_port);
   SUM_i_1 : AND2_63 port map( A => out_adder_1_port, B => n61, Y => 
                           in_cmp_1_port);
   SUM_i_2 : AND2_62 port map( A => out_adder_2_port, B => n61, Y => 
                           in_cmp_2_port);
   SUM_i_3 : AND2_61 port map( A => out_adder_3_port, B => n61, Y => 
                           in_cmp_3_port);
   SUM_i_4 : AND2_60 port map( A => out_adder_4_port, B => n61, Y => 
                           in_cmp_4_port);
   SUM_i_5 : AND2_59 port map( A => out_adder_5_port, B => n61, Y => 
                           in_cmp_5_port);
   SUM_i_6 : AND2_58 port map( A => out_adder_6_port, B => n61, Y => 
                           in_cmp_6_port);
   SUM_i_7 : AND2_57 port map( A => out_adder_7_port, B => n61, Y => 
                           in_cmp_7_port);
   SUM_i_8 : AND2_56 port map( A => out_adder_8_port, B => n61, Y => 
                           in_cmp_8_port);
   SUM_i_9 : AND2_55 port map( A => out_adder_9_port, B => n61, Y => 
                           in_cmp_9_port);
   SUM_i_10 : AND2_54 port map( A => out_adder_10_port, B => n61, Y => 
                           in_cmp_10_port);
   SUM_i_11 : AND2_53 port map( A => out_adder_11_port, B => n61, Y => 
                           in_cmp_11_port);
   SUM_i_12 : AND2_52 port map( A => out_adder_12_port, B => n61, Y => 
                           in_cmp_12_port);
   SUM_i_13 : AND2_51 port map( A => out_adder_13_port, B => n61, Y => 
                           in_cmp_13_port);
   SUM_i_14 : AND2_50 port map( A => out_adder_14_port, B => n61, Y => 
                           in_cmp_14_port);
   SUM_i_15 : AND2_49 port map( A => out_adder_15_port, B => n61, Y => 
                           in_cmp_15_port);
   SUM_i_16 : AND2_48 port map( A => out_adder_16_port, B => n61, Y => 
                           in_cmp_16_port);
   SUM_i_17 : AND2_47 port map( A => out_adder_17_port, B => n60, Y => 
                           in_cmp_17_port);
   SUM_i_18 : AND2_46 port map( A => out_adder_18_port, B => n60, Y => 
                           in_cmp_18_port);
   SUM_i_19 : AND2_45 port map( A => out_adder_19_port, B => n60, Y => 
                           in_cmp_19_port);
   SUM_i_20 : AND2_44 port map( A => out_adder_20_port, B => n60, Y => 
                           in_cmp_20_port);
   SUM_i_21 : AND2_43 port map( A => out_adder_21_port, B => n60, Y => 
                           in_cmp_21_port);
   SUM_i_22 : AND2_42 port map( A => out_adder_22_port, B => n60, Y => 
                           in_cmp_22_port);
   SUM_i_23 : AND2_41 port map( A => out_adder_23_port, B => n60, Y => 
                           in_cmp_23_port);
   SUM_i_24 : AND2_40 port map( A => out_adder_24_port, B => n60, Y => 
                           in_cmp_24_port);
   SUM_i_25 : AND2_39 port map( A => out_adder_25_port, B => n60, Y => 
                           in_cmp_25_port);
   SUM_i_26 : AND2_38 port map( A => out_adder_26_port, B => n60, Y => 
                           in_cmp_26_port);
   SUM_i_27 : AND2_37 port map( A => out_adder_27_port, B => n60, Y => 
                           in_cmp_27_port);
   SUM_i_28 : AND2_36 port map( A => out_adder_28_port, B => n60, Y => 
                           in_cmp_28_port);
   SUM_i_29 : AND2_35 port map( A => out_adder_29_port, B => n60, Y => 
                           in_cmp_29_port);
   SUM_i_30 : AND2_34 port map( A => out_adder_30_port, B => n60, Y => 
                           in_cmp_30_port);
   SUM_i_31 : AND2_33 port map( A => out_adder_31_port, B => n60, Y => 
                           in_cmp_31_port);
   MUL_A_i_0 : AND2_32 port map( A => A(0), B => n62, Y => A_mul_0_port);
   MUL_B_i_0 : AND2_31 port map( A => B(0), B => n64, Y => B_mul_0_port);
   MUL_A_i_1 : AND2_30 port map( A => A(1), B => n64, Y => A_mul_1_port);
   MUL_B_i_1 : AND2_29 port map( A => B(1), B => n64, Y => B_mul_1_port);
   MUL_A_i_2 : AND2_28 port map( A => A(2), B => n64, Y => A_mul_2_port);
   MUL_B_i_2 : AND2_27 port map( A => B(2), B => n64, Y => B_mul_2_port);
   MUL_A_i_3 : AND2_26 port map( A => A(3), B => n64, Y => A_mul_3_port);
   MUL_B_i_3 : AND2_25 port map( A => B(3), B => n64, Y => B_mul_3_port);
   MUL_A_i_4 : AND2_24 port map( A => A(4), B => n64, Y => A_mul_4_port);
   MUL_B_i_4 : AND2_23 port map( A => B(4), B => n63, Y => B_mul_4_port);
   MUL_A_i_5 : AND2_22 port map( A => A(5), B => n63, Y => A_mul_5_port);
   MUL_B_i_5 : AND2_21 port map( A => B(5), B => n63, Y => B_mul_5_port);
   MUL_A_i_6 : AND2_20 port map( A => A(6), B => n63, Y => A_mul_6_port);
   MUL_B_i_6 : AND2_19 port map( A => B(6), B => n63, Y => B_mul_6_port);
   MUL_A_i_7 : AND2_18 port map( A => A(7), B => n63, Y => A_mul_7_port);
   MUL_B_i_7 : AND2_17 port map( A => B(7), B => n63, Y => B_mul_7_port);
   MUL_A_i_8 : AND2_16 port map( A => A(8), B => n63, Y => A_mul_8_port);
   MUL_B_i_8 : AND2_15 port map( A => B(8), B => n63, Y => B_mul_8_port);
   MUL_A_i_9 : AND2_14 port map( A => A(9), B => n63, Y => A_mul_9_port);
   MUL_B_i_9 : AND2_13 port map( A => B(9), B => n63, Y => B_mul_9_port);
   MUL_A_i_10 : AND2_12 port map( A => A(10), B => n62, Y => A_mul_10_port);
   MUL_B_i_10 : AND2_11 port map( A => B(10), B => n62, Y => B_mul_10_port);
   MUL_A_i_11 : AND2_10 port map( A => A(11), B => n62, Y => A_mul_11_port);
   MUL_B_i_11 : AND2_9 port map( A => B(11), B => n62, Y => B_mul_11_port);
   MUL_A_i_12 : AND2_8 port map( A => A(12), B => n62, Y => A_mul_12_port);
   MUL_B_i_12 : AND2_7 port map( A => B(12), B => n63, Y => B_mul_12_port);
   MUL_A_i_13 : AND2_6 port map( A => A(13), B => n62, Y => A_mul_13_port);
   MUL_B_i_13 : AND2_5 port map( A => B(13), B => n62, Y => B_mul_13_port);
   MUL_A_i_14 : AND2_4 port map( A => A(14), B => n62, Y => A_mul_14_port);
   MUL_B_i_14 : AND2_3 port map( A => B(14), B => n62, Y => B_mul_14_port);
   MUL_A_i_15 : AND2_2 port map( A => A(15), B => n62, Y => A_mul_15_port);
   MUL_B_i_15 : AND2_1 port map( A => B(15), B => n62, Y => B_mul_15_port);
   ADD : ADDER_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A_adder_31_port, 
                           A(30) => A_adder_30_port, A(29) => A_adder_29_port, 
                           A(28) => A_adder_28_port, A(27) => A_adder_27_port, 
                           A(26) => A_adder_26_port, A(25) => A_adder_25_port, 
                           A(24) => A_adder_24_port, A(23) => A_adder_23_port, 
                           A(22) => A_adder_22_port, A(21) => A_adder_21_port, 
                           A(20) => A_adder_20_port, A(19) => A_adder_19_port, 
                           A(18) => A_adder_18_port, A(17) => A_adder_17_port, 
                           A(16) => A_adder_16_port, A(15) => A_adder_15_port, 
                           A(14) => A_adder_14_port, A(13) => A_adder_13_port, 
                           A(12) => A_adder_12_port, A(11) => A_adder_11_port, 
                           A(10) => A_adder_10_port, A(9) => A_adder_9_port, 
                           A(8) => A_adder_8_port, A(7) => A_adder_7_port, A(6)
                           => A_adder_6_port, A(5) => A_adder_5_port, A(4) => 
                           A_adder_4_port, A(3) => A_adder_3_port, A(2) => 
                           A_adder_2_port, A(1) => A_adder_1_port, A(0) => 
                           A_adder_0_port, B(31) => B_adder_31_port, B(30) => 
                           B_adder_30_port, B(29) => B_adder_29_port, B(28) => 
                           B_adder_28_port, B(27) => B_adder_27_port, B(26) => 
                           B_adder_26_port, B(25) => B_adder_25_port, B(24) => 
                           B_adder_24_port, B(23) => B_adder_23_port, B(22) => 
                           B_adder_22_port, B(21) => B_adder_21_port, B(20) => 
                           B_adder_20_port, B(19) => B_adder_19_port, B(18) => 
                           B_adder_18_port, B(17) => B_adder_17_port, B(16) => 
                           B_adder_16_port, B(15) => B_adder_15_port, B(14) => 
                           B_adder_14_port, B(13) => B_adder_13_port, B(12) => 
                           B_adder_12_port, B(11) => B_adder_11_port, B(10) => 
                           B_adder_10_port, B(9) => B_adder_9_port, B(8) => 
                           B_adder_8_port, B(7) => B_adder_7_port, B(6) => 
                           B_adder_6_port, B(5) => B_adder_5_port, B(4) => 
                           B_adder_4_port, B(3) => B_adder_3_port, B(2) => 
                           B_adder_2_port, B(1) => B_adder_1_port, B(0) => 
                           B_adder_0_port, ADD_SUB => n91_port, Cin => 
                           cin_internal, S(31) => out_adder_31_port, S(30) => 
                           out_adder_30_port, S(29) => out_adder_29_port, S(28)
                           => out_adder_28_port, S(27) => out_adder_27_port, 
                           S(26) => out_adder_26_port, S(25) => 
                           out_adder_25_port, S(24) => out_adder_24_port, S(23)
                           => out_adder_23_port, S(22) => out_adder_22_port, 
                           S(21) => out_adder_21_port, S(20) => 
                           out_adder_20_port, S(19) => out_adder_19_port, S(18)
                           => out_adder_18_port, S(17) => out_adder_17_port, 
                           S(16) => out_adder_16_port, S(15) => 
                           out_adder_15_port, S(14) => out_adder_14_port, S(13)
                           => out_adder_13_port, S(12) => out_adder_12_port, 
                           S(11) => out_adder_11_port, S(10) => 
                           out_adder_10_port, S(9) => out_adder_9_port, S(8) =>
                           out_adder_8_port, S(7) => out_adder_7_port, S(6) => 
                           out_adder_6_port, S(5) => out_adder_5_port, S(4) => 
                           out_adder_4_port, S(3) => out_adder_3_port, S(2) => 
                           out_adder_2_port, S(1) => out_adder_1_port, S(0) => 
                           out_adder_0_port, Cout => Cout_port);
   SHIFT : SHIFTER port map( data_in(31) => A_shifter_31_port, data_in(30) => 
                           A_shifter_30_port, data_in(29) => A_shifter_29_port,
                           data_in(28) => A_shifter_28_port, data_in(27) => 
                           A_shifter_27_port, data_in(26) => A_shifter_26_port,
                           data_in(25) => A_shifter_25_port, data_in(24) => 
                           A_shifter_24_port, data_in(23) => A_shifter_23_port,
                           data_in(22) => A_shifter_22_port, data_in(21) => 
                           A_shifter_21_port, data_in(20) => A_shifter_20_port,
                           data_in(19) => A_shifter_19_port, data_in(18) => 
                           A_shifter_18_port, data_in(17) => A_shifter_17_port,
                           data_in(16) => A_shifter_16_port, data_in(15) => 
                           A_shifter_15_port, data_in(14) => A_shifter_14_port,
                           data_in(13) => A_shifter_13_port, data_in(12) => 
                           A_shifter_12_port, data_in(11) => A_shifter_11_port,
                           data_in(10) => A_shifter_10_port, data_in(9) => 
                           A_shifter_9_port, data_in(8) => A_shifter_8_port, 
                           data_in(7) => A_shifter_7_port, data_in(6) => 
                           A_shifter_6_port, data_in(5) => A_shifter_5_port, 
                           data_in(4) => A_shifter_4_port, data_in(3) => 
                           A_shifter_3_port, data_in(2) => A_shifter_2_port, 
                           data_in(1) => A_shifter_1_port, data_in(0) => 
                           A_shifter_0_port, R(4) => B_shifter_4_port, R(3) => 
                           B_shifter_3_port, R(2) => B_shifter_2_port, R(1) => 
                           B_shifter_1_port, R(0) => B_shifter_0_port, conf(1) 
                           => conf_1_port, conf(0) => conf_0_port, data_out(31)
                           => out_shifter_31_port, data_out(30) => 
                           out_shifter_30_port, data_out(29) => 
                           out_shifter_29_port, data_out(28) => 
                           out_shifter_28_port, data_out(27) => 
                           out_shifter_27_port, data_out(26) => 
                           out_shifter_26_port, data_out(25) => 
                           out_shifter_25_port, data_out(24) => 
                           out_shifter_24_port, data_out(23) => 
                           out_shifter_23_port, data_out(22) => 
                           out_shifter_22_port, data_out(21) => 
                           out_shifter_21_port, data_out(20) => 
                           out_shifter_20_port, data_out(19) => 
                           out_shifter_19_port, data_out(18) => 
                           out_shifter_18_port, data_out(17) => 
                           out_shifter_17_port, data_out(16) => 
                           out_shifter_16_port, data_out(15) => 
                           out_shifter_15_port, data_out(14) => 
                           out_shifter_14_port, data_out(13) => 
                           out_shifter_13_port, data_out(12) => 
                           out_shifter_12_port, data_out(11) => 
                           out_shifter_11_port, data_out(10) => 
                           out_shifter_10_port, data_out(9) => 
                           out_shifter_9_port, data_out(8) => 
                           out_shifter_8_port, data_out(7) => 
                           out_shifter_7_port, data_out(6) => 
                           out_shifter_6_port, data_out(5) => 
                           out_shifter_5_port, data_out(4) => 
                           out_shifter_4_port, data_out(3) => 
                           out_shifter_3_port, data_out(2) => 
                           out_shifter_2_port, data_out(1) => 
                           out_shifter_1_port, data_out(0) => 
                           out_shifter_0_port);
   LOGICALS : LOGIC_NBIT32_N_SELECTOR4 port map( S(3) => logic_sel_3_port, S(2)
                           => logic_sel_2_port, S(1) => logic_sel_1_port, S(0) 
                           => logic_sel_0_port, A(31) => A_logic_31_port, A(30)
                           => A_logic_30_port, A(29) => A_logic_29_port, A(28) 
                           => A_logic_28_port, A(27) => A_logic_27_port, A(26) 
                           => A_logic_26_port, A(25) => A_logic_25_port, A(24) 
                           => A_logic_24_port, A(23) => A_logic_23_port, A(22) 
                           => A_logic_22_port, A(21) => A_logic_21_port, A(20) 
                           => A_logic_20_port, A(19) => A_logic_19_port, A(18) 
                           => A_logic_18_port, A(17) => A_logic_17_port, A(16) 
                           => A_logic_16_port, A(15) => A_logic_15_port, A(14) 
                           => A_logic_14_port, A(13) => A_logic_13_port, A(12) 
                           => A_logic_12_port, A(11) => A_logic_11_port, A(10) 
                           => A_logic_10_port, A(9) => A_logic_9_port, A(8) => 
                           A_logic_8_port, A(7) => A_logic_7_port, A(6) => 
                           A_logic_6_port, A(5) => A_logic_5_port, A(4) => 
                           A_logic_4_port, A(3) => A_logic_3_port, A(2) => 
                           A_logic_2_port, A(1) => A_logic_1_port, A(0) => 
                           A_logic_0_port, B(31) => B_logic_31_port, B(30) => 
                           B_logic_30_port, B(29) => B_logic_29_port, B(28) => 
                           B_logic_28_port, B(27) => B_logic_27_port, B(26) => 
                           B_logic_26_port, B(25) => B_logic_25_port, B(24) => 
                           B_logic_24_port, B(23) => B_logic_23_port, B(22) => 
                           B_logic_22_port, B(21) => B_logic_21_port, B(20) => 
                           B_logic_20_port, B(19) => B_logic_19_port, B(18) => 
                           B_logic_18_port, B(17) => B_logic_17_port, B(16) => 
                           B_logic_16_port, B(15) => B_logic_15_port, B(14) => 
                           B_logic_14_port, B(13) => B_logic_13_port, B(12) => 
                           B_logic_12_port, B(11) => B_logic_11_port, B(10) => 
                           B_logic_10_port, B(9) => B_logic_9_port, B(8) => 
                           B_logic_8_port, B(7) => B_logic_7_port, B(6) => 
                           B_logic_6_port, B(5) => B_logic_5_port, B(4) => 
                           B_logic_4_port, B(3) => B_logic_3_port, B(2) => 
                           B_logic_2_port, B(1) => B_logic_1_port, B(0) => 
                           B_logic_0_port, O(31) => out_logic_31_port, O(30) =>
                           out_logic_30_port, O(29) => out_logic_29_port, O(28)
                           => out_logic_28_port, O(27) => out_logic_27_port, 
                           O(26) => out_logic_26_port, O(25) => 
                           out_logic_25_port, O(24) => out_logic_24_port, O(23)
                           => out_logic_23_port, O(22) => out_logic_22_port, 
                           O(21) => out_logic_21_port, O(20) => 
                           out_logic_20_port, O(19) => out_logic_19_port, O(18)
                           => out_logic_18_port, O(17) => out_logic_17_port, 
                           O(16) => out_logic_16_port, O(15) => 
                           out_logic_15_port, O(14) => out_logic_14_port, O(13)
                           => out_logic_13_port, O(12) => out_logic_12_port, 
                           O(11) => out_logic_11_port, O(10) => 
                           out_logic_10_port, O(9) => out_logic_9_port, O(8) =>
                           out_logic_8_port, O(7) => out_logic_7_port, O(6) => 
                           out_logic_6_port, O(5) => out_logic_5_port, O(4) => 
                           out_logic_4_port, O(3) => out_logic_3_port, O(2) => 
                           out_logic_2_port, O(1) => out_logic_1_port, O(0) => 
                           out_logic_0_port);
   COMPARATOR : CMP_NBIT32 port map( SUM(31) => in_cmp_31_port, SUM(30) => 
                           in_cmp_30_port, SUM(29) => in_cmp_29_port, SUM(28) 
                           => in_cmp_28_port, SUM(27) => in_cmp_27_port, 
                           SUM(26) => in_cmp_26_port, SUM(25) => in_cmp_25_port
                           , SUM(24) => in_cmp_24_port, SUM(23) => 
                           in_cmp_23_port, SUM(22) => in_cmp_22_port, SUM(21) 
                           => in_cmp_21_port, SUM(20) => in_cmp_20_port, 
                           SUM(19) => in_cmp_19_port, SUM(18) => in_cmp_18_port
                           , SUM(17) => in_cmp_17_port, SUM(16) => 
                           in_cmp_16_port, SUM(15) => in_cmp_15_port, SUM(14) 
                           => in_cmp_14_port, SUM(13) => in_cmp_13_port, 
                           SUM(12) => in_cmp_12_port, SUM(11) => in_cmp_11_port
                           , SUM(10) => in_cmp_10_port, SUM(9) => in_cmp_9_port
                           , SUM(8) => in_cmp_8_port, SUM(7) => in_cmp_7_port, 
                           SUM(6) => in_cmp_6_port, SUM(5) => in_cmp_5_port, 
                           SUM(4) => in_cmp_4_port, SUM(3) => in_cmp_3_port, 
                           SUM(2) => in_cmp_2_port, SUM(1) => in_cmp_1_port, 
                           SUM(0) => in_cmp_0_port, Cout => Cout_port, A_L_B =>
                           COND(0), A_LE_B => COND(1), A_G_B => COND(2), A_GE_B
                           => COND(3), A_E_B => COND(4), A_NE_B => COND(5));
   MULTIPLIER : MUL port map( CLOCK => CLOCK, A(15) => A_mul_15_port, A(14) => 
                           A_mul_14_port, A(13) => A_mul_13_port, A(12) => 
                           A_mul_12_port, A(11) => A_mul_11_port, A(10) => 
                           A_mul_10_port, A(9) => A_mul_9_port, A(8) => 
                           A_mul_8_port, A(7) => A_mul_7_port, A(6) => 
                           A_mul_6_port, A(5) => A_mul_5_port, A(4) => 
                           A_mul_4_port, A(3) => A_mul_3_port, A(2) => 
                           A_mul_2_port, A(1) => A_mul_1_port, A(0) => 
                           A_mul_0_port, B(15) => B_mul_15_port, B(14) => 
                           B_mul_14_port, B(13) => B_mul_13_port, B(12) => 
                           B_mul_12_port, B(11) => B_mul_11_port, B(10) => 
                           B_mul_10_port, B(9) => B_mul_9_port, B(8) => 
                           B_mul_8_port, B(7) => B_mul_7_port, B(6) => 
                           B_mul_6_port, B(5) => B_mul_5_port, B(4) => 
                           B_mul_4_port, B(3) => B_mul_3_port, B(2) => 
                           B_mul_2_port, B(1) => B_mul_1_port, B(0) => 
                           B_mul_0_port, Y(31) => out_mul_31_port, Y(30) => 
                           out_mul_30_port, Y(29) => out_mul_29_port, Y(28) => 
                           out_mul_28_port, Y(27) => out_mul_27_port, Y(26) => 
                           out_mul_26_port, Y(25) => out_mul_25_port, Y(24) => 
                           out_mul_24_port, Y(23) => out_mul_23_port, Y(22) => 
                           out_mul_22_port, Y(21) => out_mul_21_port, Y(20) => 
                           out_mul_20_port, Y(19) => out_mul_19_port, Y(18) => 
                           out_mul_18_port, Y(17) => out_mul_17_port, Y(16) => 
                           out_mul_16_port, Y(15) => out_mul_15_port, Y(14) => 
                           out_mul_14_port, Y(13) => out_mul_13_port, Y(12) => 
                           out_mul_12_port, Y(11) => out_mul_11_port, Y(10) => 
                           out_mul_10_port, Y(9) => out_mul_9_port, Y(8) => 
                           out_mul_8_port, Y(7) => out_mul_7_port, Y(6) => 
                           out_mul_6_port, Y(5) => out_mul_5_port, Y(4) => 
                           out_mul_4_port, Y(3) => out_mul_3_port, Y(2) => 
                           out_mul_2_port, Y(1) => out_mul_1_port, Y(0) => 
                           out_mul_0_port);
   OUTPUT_SEL : MUX4to1_NBIT32_1 port map( A(31) => out_adder_31_port, A(30) =>
                           out_adder_30_port, A(29) => out_adder_29_port, A(28)
                           => out_adder_28_port, A(27) => out_adder_27_port, 
                           A(26) => out_adder_26_port, A(25) => 
                           out_adder_25_port, A(24) => out_adder_24_port, A(23)
                           => out_adder_23_port, A(22) => out_adder_22_port, 
                           A(21) => out_adder_21_port, A(20) => 
                           out_adder_20_port, A(19) => out_adder_19_port, A(18)
                           => out_adder_18_port, A(17) => out_adder_17_port, 
                           A(16) => out_adder_16_port, A(15) => 
                           out_adder_15_port, A(14) => out_adder_14_port, A(13)
                           => out_adder_13_port, A(12) => out_adder_12_port, 
                           A(11) => out_adder_11_port, A(10) => 
                           out_adder_10_port, A(9) => out_adder_9_port, A(8) =>
                           out_adder_8_port, A(7) => out_adder_7_port, A(6) => 
                           out_adder_6_port, A(5) => out_adder_5_port, A(4) => 
                           out_adder_4_port, A(3) => out_adder_3_port, A(2) => 
                           out_adder_2_port, A(1) => out_adder_1_port, A(0) => 
                           out_adder_0_port, B(31) => out_logic_31_port, B(30) 
                           => out_logic_30_port, B(29) => out_logic_29_port, 
                           B(28) => out_logic_28_port, B(27) => 
                           out_logic_27_port, B(26) => out_logic_26_port, B(25)
                           => out_logic_25_port, B(24) => out_logic_24_port, 
                           B(23) => out_logic_23_port, B(22) => 
                           out_logic_22_port, B(21) => out_logic_21_port, B(20)
                           => out_logic_20_port, B(19) => out_logic_19_port, 
                           B(18) => out_logic_18_port, B(17) => 
                           out_logic_17_port, B(16) => out_logic_16_port, B(15)
                           => out_logic_15_port, B(14) => out_logic_14_port, 
                           B(13) => out_logic_13_port, B(12) => 
                           out_logic_12_port, B(11) => out_logic_11_port, B(10)
                           => out_logic_10_port, B(9) => out_logic_9_port, B(8)
                           => out_logic_8_port, B(7) => out_logic_7_port, B(6) 
                           => out_logic_6_port, B(5) => out_logic_5_port, B(4) 
                           => out_logic_4_port, B(3) => out_logic_3_port, B(2) 
                           => out_logic_2_port, B(1) => out_logic_1_port, B(0) 
                           => out_logic_0_port, C(31) => out_shifter_31_port, 
                           C(30) => out_shifter_30_port, C(29) => 
                           out_shifter_29_port, C(28) => out_shifter_28_port, 
                           C(27) => out_shifter_27_port, C(26) => 
                           out_shifter_26_port, C(25) => out_shifter_25_port, 
                           C(24) => out_shifter_24_port, C(23) => 
                           out_shifter_23_port, C(22) => out_shifter_22_port, 
                           C(21) => out_shifter_21_port, C(20) => 
                           out_shifter_20_port, C(19) => out_shifter_19_port, 
                           C(18) => out_shifter_18_port, C(17) => 
                           out_shifter_17_port, C(16) => out_shifter_16_port, 
                           C(15) => out_shifter_15_port, C(14) => 
                           out_shifter_14_port, C(13) => out_shifter_13_port, 
                           C(12) => out_shifter_12_port, C(11) => 
                           out_shifter_11_port, C(10) => out_shifter_10_port, 
                           C(9) => out_shifter_9_port, C(8) => 
                           out_shifter_8_port, C(7) => out_shifter_7_port, C(6)
                           => out_shifter_6_port, C(5) => out_shifter_5_port, 
                           C(4) => out_shifter_4_port, C(3) => 
                           out_shifter_3_port, C(2) => out_shifter_2_port, C(1)
                           => out_shifter_1_port, C(0) => out_shifter_0_port, 
                           D(31) => out_mul_31_port, D(30) => out_mul_30_port, 
                           D(29) => out_mul_29_port, D(28) => out_mul_28_port, 
                           D(27) => out_mul_27_port, D(26) => out_mul_26_port, 
                           D(25) => out_mul_25_port, D(24) => out_mul_24_port, 
                           D(23) => out_mul_23_port, D(22) => out_mul_22_port, 
                           D(21) => out_mul_21_port, D(20) => out_mul_20_port, 
                           D(19) => out_mul_19_port, D(18) => out_mul_18_port, 
                           D(17) => out_mul_17_port, D(16) => out_mul_16_port, 
                           D(15) => out_mul_15_port, D(14) => out_mul_14_port, 
                           D(13) => out_mul_13_port, D(12) => out_mul_12_port, 
                           D(11) => out_mul_11_port, D(10) => out_mul_10_port, 
                           D(9) => out_mul_9_port, D(8) => out_mul_8_port, D(7)
                           => out_mul_7_port, D(6) => out_mul_6_port, D(5) => 
                           out_mul_5_port, D(4) => out_mul_4_port, D(3) => 
                           out_mul_3_port, D(2) => out_mul_2_port, D(1) => 
                           out_mul_1_port, D(0) => out_mul_0_port, SEL(1) => 
                           mux_out_1_port, SEL(0) => mux_out_0_port, Y(31) => 
                           ALU_out(31), Y(30) => ALU_out(30), Y(29) => 
                           ALU_out(29), Y(28) => ALU_out(28), Y(27) => 
                           ALU_out(27), Y(26) => ALU_out(26), Y(25) => 
                           ALU_out(25), Y(24) => ALU_out(24), Y(23) => 
                           ALU_out(23), Y(22) => ALU_out(22), Y(21) => 
                           ALU_out(21), Y(20) => ALU_out(20), Y(19) => 
                           ALU_out(19), Y(18) => ALU_out(18), Y(17) => 
                           ALU_out(17), Y(16) => ALU_out(16), Y(15) => 
                           ALU_out(15), Y(14) => ALU_out(14), Y(13) => 
                           ALU_out(13), Y(12) => ALU_out(12), Y(11) => 
                           ALU_out(11), Y(10) => ALU_out(10), Y(9) => 
                           ALU_out(9), Y(8) => ALU_out(8), Y(7) => ALU_out(7), 
                           Y(6) => ALU_out(6), Y(5) => ALU_out(5), Y(4) => 
                           ALU_out(4), Y(3) => ALU_out(3), Y(2) => ALU_out(2), 
                           Y(1) => ALU_out(1), Y(0) => ALU_out(0));
   U3 : BUF_X1 port map( A => n72, Z => n70);
   U4 : BUF_X1 port map( A => en_logic, Z => n80);
   U5 : BUF_X1 port map( A => en_logic, Z => n79);
   U6 : BUF_X1 port map( A => n81, Z => n88_port);
   U7 : BUF_X1 port map( A => n81, Z => n89_port);
   U8 : BUF_X1 port map( A => n1, Z => n65);
   U9 : BUF_X1 port map( A => n70, Z => n68);
   U10 : BUF_X1 port map( A => n70, Z => n67);
   U11 : BUF_X1 port map( A => n70, Z => n69);
   U12 : OR2_X1 port map( A1 => n64, A2 => n69, ZN => mux_out_1_port);
   U13 : OR2_X1 port map( A1 => n78, A2 => n64, ZN => mux_out_0_port);
   U14 : INV_X1 port map( A => n10, ZN => n91_port);
   U15 : BUF_X1 port map( A => n80, Z => n73);
   U16 : BUF_X1 port map( A => n80, Z => n74);
   U17 : BUF_X1 port map( A => n80, Z => n75);
   U18 : BUF_X1 port map( A => n79, Z => n76);
   U19 : BUF_X1 port map( A => n79, Z => n77);
   U20 : BUF_X1 port map( A => n89_port, Z => n83);
   U21 : BUF_X1 port map( A => n88_port, Z => n85);
   U22 : BUF_X1 port map( A => n89_port, Z => n82);
   U23 : BUF_X1 port map( A => n89_port, Z => n84);
   U24 : BUF_X1 port map( A => n88_port, Z => n86);
   U25 : BUF_X1 port map( A => n71, Z => n66);
   U26 : BUF_X1 port map( A => n72, Z => n71);
   U27 : BUF_X1 port map( A => n79, Z => n78);
   U28 : BUF_X1 port map( A => n88_port, Z => n87);
   U29 : AOI21_X1 port map( B1 => n96, B2 => n17, A => n60, ZN => n10);
   U30 : NOR3_X1 port map( A1 => n12, A2 => n94, A3 => n96, ZN => N92);
   U31 : INV_X1 port map( A => n13, ZN => n95);
   U32 : NAND2_X1 port map( A1 => n20, A2 => n96, ZN => n21);
   U33 : BUF_X1 port map( A => en_shifter, Z => n72);
   U34 : NOR2_X1 port map( A1 => n12, A2 => n13, ZN => en_shifter);
   U35 : BUF_X1 port map( A => n92_port, Z => n61);
   U36 : BUF_X1 port map( A => n92_port, Z => n60);
   U37 : BUF_X1 port map( A => n65, Z => n63);
   U38 : BUF_X1 port map( A => n65, Z => n62);
   U42 : BUF_X1 port map( A => n65, Z => n64);
   U43 : OAI221_X1 port map( B1 => n11, B2 => n21, C1 => n95, C2 => n12, A => 
                           n26, ZN => N89);
   U44 : OR3_X1 port map( A1 => N88, A2 => N89, A3 => n14, ZN => en_logic);
   U45 : AND3_X1 port map( A1 => AluOpcode(3), A2 => n15, A3 => n13, ZN => n14)
                           ;
   U46 : NOR2_X1 port map( A1 => n96, A2 => AluOpcode(1), ZN => n13);
   U47 : NOR2_X1 port map( A1 => AluOpcode(2), A2 => AluOpcode(1), ZN => n20);
   U48 : NOR2_X1 port map( A1 => AluOpcode(2), A2 => AluOpcode(0), ZN => n15);
   U49 : AOI211_X1 port map( C1 => n15, C2 => n97, A => n24, B => n95, ZN => 
                           N90);
   U50 : NAND2_X1 port map( A1 => n25, A2 => n11, ZN => n24);
   U51 : OAI21_X1 port map( B1 => AluOpcode(3), B2 => AluOpcode(0), A => 
                           AluOpcode(2), ZN => n25);
   U52 : OAI22_X1 port map( A1 => n20, A2 => n93_port, B1 => AluOpcode(3), B2 
                           => n22, ZN => N91);
   U53 : AOI22_X1 port map( A1 => n23, A2 => n96, B1 => AluOpcode(2), B2 => 
                           AluOpcode(1), ZN => n22);
   U54 : NOR2_X1 port map( A1 => AluOpcode(0), A2 => AluOpcode(1), ZN => n23);
   U55 : NOR4_X1 port map( A1 => n90_port, A2 => n21, A3 => n97, A4 => 
                           AluOpcode(0), ZN => cin_internal);
   U56 : INV_X1 port map( A => Cin, ZN => n90_port);
   U57 : AOI21_X1 port map( B1 => n27, B2 => n21, A => n93_port, ZN => N88);
   U58 : OR3_X1 port map( A1 => n95, A2 => AluOpcode(2), A3 => AluOpcode(3), ZN
                           => n27);
   U59 : INV_X1 port map( A => AluOpcode(4), ZN => n96);
   U60 : NOR3_X1 port map( A1 => n12, A2 => AluOpcode(1), A3 => AluOpcode(4), 
                           ZN => N93);
   U61 : NAND2_X1 port map( A1 => AluOpcode(0), A2 => AluOpcode(3), ZN => n11);
   U62 : INV_X1 port map( A => AluOpcode(3), ZN => n97);
   U63 : INV_X1 port map( A => AluOpcode(0), ZN => n93_port);
   U64 : INV_X1 port map( A => AluOpcode(1), ZN => n94);
   U65 : AND3_X1 port map( A1 => AluOpcode(3), A2 => n93_port, A3 => 
                           AluOpcode(2), ZN => n17);
   U66 : NOR3_X1 port map( A1 => n11, A2 => AluOpcode(2), A3 => n95, ZN => n1);
   U67 : BUF_X1 port map( A => en_adder, Z => n81);
   U68 : NAND2_X1 port map( A1 => n16, A2 => n10, ZN => en_adder);
   U69 : XNOR2_X1 port map( A => n97, B => AluOpcode(4), ZN => n19);
   U70 : INV_X1 port map( A => n18, ZN => n92_port);
   U71 : AOI22_X1 port map( A1 => n94, A2 => n17, B1 => n15, B2 => AluOpcode(1)
                           , ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT5 is

   port( A, B, C : in std_logic_vector (4 downto 0);  SEL : in std_logic_vector
         (1 downto 0);  Y : out std_logic_vector (4 downto 0));

end MUX3to1_NBIT5;

architecture SYN_Behavioral of MUX3to1_NBIT5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n7, n8, n9, n10, n11, n12_port, n13, n14, n15, n16, n17, n18, 
      n19, n20 : std_logic;

begin
   
   Y_reg_4_inst : DLH_X1 port map( G => N12, D => n15, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => N12, D => n16, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => N12, D => n17, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => n18, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => n19, Q => Y(0));
   U3 : NOR2_X1 port map( A1 => n20, A2 => SEL(1), ZN => n9);
   U4 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n8);
   U5 : AND2_X1 port map( A1 => SEL(1), A2 => n20, ZN => n10);
   U6 : NAND2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => N12);
   U7 : INV_X1 port map( A => SEL(0), ZN => n20);
   U8 : INV_X1 port map( A => n14, ZN => n19);
   U9 : AOI222_X1 port map( A1 => A(0), A2 => n8, B1 => B(0), B2 => n9, C1 => 
                           C(0), C2 => n10, ZN => n14);
   U10 : INV_X1 port map( A => n13, ZN => n18);
   U11 : AOI222_X1 port map( A1 => A(1), A2 => n8, B1 => B(1), B2 => n9, C1 => 
                           C(1), C2 => n10, ZN => n13);
   U12 : INV_X1 port map( A => n12_port, ZN => n17);
   U13 : AOI222_X1 port map( A1 => A(2), A2 => n8, B1 => B(2), B2 => n9, C1 => 
                           C(2), C2 => n10, ZN => n12_port);
   U14 : INV_X1 port map( A => n11, ZN => n16);
   U15 : AOI222_X1 port map( A1 => A(3), A2 => n8, B1 => B(3), B2 => n9, C1 => 
                           C(3), C2 => n10, ZN => n11);
   U16 : INV_X1 port map( A => n7, ZN => n15);
   U17 : AOI222_X1 port map( A1 => A(4), A2 => n8, B1 => B(4), B2 => n9, C1 => 
                           C(4), C2 => n10, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_1;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n105, n106, n107, n108, n109, n110, n111, n112 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n108, Z => n112);
   U2 : BUF_X1 port map( A => n108, Z => n111);
   U3 : BUF_X1 port map( A => SEL, Z => n108);
   U4 : INV_X1 port map( A => n111, ZN => n109);
   U5 : INV_X1 port map( A => n111, ZN => n110);
   U6 : BUF_X1 port map( A => n112, Z => n105);
   U7 : BUF_X1 port map( A => n112, Z => n106);
   U8 : BUF_X1 port map( A => n112, Z => n107);
   U9 : INV_X1 port map( A => n65, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n109, B1 => B(0), B2 => n105, ZN 
                           => n65);
   U11 : INV_X1 port map( A => n64, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n109, B1 => B(1), B2 => n105, ZN 
                           => n64);
   U13 : INV_X1 port map( A => n63, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => n109, B1 => B(2), B2 => n105, ZN 
                           => n63);
   U15 : INV_X1 port map( A => n62, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n109, B1 => B(3), B2 => n105, ZN 
                           => n62);
   U17 : INV_X1 port map( A => n61, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n109, B1 => B(4), B2 => n105, ZN 
                           => n61);
   U19 : INV_X1 port map( A => n60, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n109, B1 => B(5), B2 => n105, ZN 
                           => n60);
   U21 : INV_X1 port map( A => n59, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n109, B1 => B(6), B2 => n105, ZN 
                           => n59);
   U23 : INV_X1 port map( A => n58, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n109, B1 => B(7), B2 => n105, ZN 
                           => n58);
   U25 : INV_X1 port map( A => n57, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n109, B1 => B(8), B2 => n105, ZN 
                           => n57);
   U27 : INV_X1 port map( A => n56, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n109, B1 => B(9), B2 => n105, ZN 
                           => n56);
   U29 : INV_X1 port map( A => n55, ZN => Y(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n109, B1 => B(10), B2 => n105, 
                           ZN => n55);
   U31 : INV_X1 port map( A => n54, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => A(11), A2 => n109, B1 => B(11), B2 => n105, 
                           ZN => n54);
   U33 : INV_X1 port map( A => n53, ZN => Y(12));
   U34 : AOI22_X1 port map( A1 => A(12), A2 => n110, B1 => B(12), B2 => n106, 
                           ZN => n53);
   U35 : INV_X1 port map( A => n52, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n110, B1 => B(13), B2 => n106, 
                           ZN => n52);
   U37 : INV_X1 port map( A => n51, ZN => Y(14));
   U38 : AOI22_X1 port map( A1 => A(14), A2 => n110, B1 => B(14), B2 => n106, 
                           ZN => n51);
   U39 : INV_X1 port map( A => n50, ZN => Y(15));
   U40 : AOI22_X1 port map( A1 => A(15), A2 => n110, B1 => B(15), B2 => n106, 
                           ZN => n50);
   U41 : INV_X1 port map( A => n49, ZN => Y(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n110, B1 => B(16), B2 => n106, 
                           ZN => n49);
   U43 : INV_X1 port map( A => n48, ZN => Y(17));
   U44 : AOI22_X1 port map( A1 => A(17), A2 => n110, B1 => B(17), B2 => n106, 
                           ZN => n48);
   U45 : INV_X1 port map( A => n47, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n110, B1 => B(18), B2 => n106, 
                           ZN => n47);
   U47 : INV_X1 port map( A => n46, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n110, B1 => B(19), B2 => n106, 
                           ZN => n46);
   U49 : INV_X1 port map( A => n45, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n110, B1 => B(20), B2 => n106, 
                           ZN => n45);
   U51 : INV_X1 port map( A => n44, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n110, B1 => B(21), B2 => n106, 
                           ZN => n44);
   U53 : INV_X1 port map( A => n43, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n110, B1 => B(22), B2 => n106, 
                           ZN => n43);
   U55 : INV_X1 port map( A => n42, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n110, B1 => B(23), B2 => n106, 
                           ZN => n42);
   U57 : INV_X1 port map( A => n41, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A(24), A2 => n110, B1 => B(24), B2 => n107, 
                           ZN => n41);
   U59 : INV_X1 port map( A => n40, ZN => Y(25));
   U60 : AOI22_X1 port map( A1 => A(25), A2 => n110, B1 => B(25), B2 => n107, 
                           ZN => n40);
   U61 : INV_X1 port map( A => n39, ZN => Y(26));
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n109, B1 => B(26), B2 => n107, 
                           ZN => n39);
   U63 : INV_X1 port map( A => n38, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n110, B1 => B(27), B2 => n107, 
                           ZN => n38);
   U65 : INV_X1 port map( A => n37, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n109, B1 => B(28), B2 => n107, 
                           ZN => n37);
   U67 : INV_X1 port map( A => n36, ZN => Y(29));
   U68 : AOI22_X1 port map( A1 => A(29), A2 => n110, B1 => B(29), B2 => n107, 
                           ZN => n36);
   U69 : INV_X1 port map( A => n35, ZN => Y(30));
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n109, B1 => B(30), B2 => n107, 
                           ZN => n35);
   U71 : INV_X1 port map( A => n34, ZN => Y(31));
   U72 : AOI22_X1 port map( A1 => A(31), A2 => n109, B1 => n107, B2 => B(31), 
                           ZN => n34);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX4to1_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX4to1_NBIT32_0;

architecture SYN_Behavioral of MUX4to1_NBIT32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102 : std_logic
      ;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n93);
   U2 : BUF_X1 port map( A => n7, Z => n89);
   U3 : BUF_X1 port map( A => n4, Z => n98);
   U4 : BUF_X1 port map( A => n5, Z => n94);
   U5 : BUF_X1 port map( A => n93, Z => n90);
   U6 : BUF_X1 port map( A => n93, Z => n91);
   U7 : BUF_X1 port map( A => n98, Z => n99);
   U8 : BUF_X1 port map( A => n98, Z => n100);
   U9 : BUF_X1 port map( A => n89, Z => n86);
   U10 : BUF_X1 port map( A => n89, Z => n87);
   U11 : BUF_X1 port map( A => n94, Z => n95);
   U12 : BUF_X1 port map( A => n94, Z => n96);
   U13 : BUF_X1 port map( A => n93, Z => n92);
   U14 : BUF_X1 port map( A => n98, Z => n101);
   U15 : BUF_X1 port map( A => n89, Z => n88);
   U16 : BUF_X1 port map( A => n94, Z => n97);
   U17 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(16));
   U18 : AOI22_X1 port map( A1 => A(16), A2 => n90, B1 => B(16), B2 => n86, ZN 
                           => n54);
   U19 : AOI22_X1 port map( A1 => C(16), A2 => n99, B1 => D(16), B2 => n95, ZN 
                           => n55);
   U20 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(17));
   U21 : AOI22_X1 port map( A1 => A(17), A2 => n90, B1 => B(17), B2 => n86, ZN 
                           => n52);
   U22 : AOI22_X1 port map( A1 => C(17), A2 => n99, B1 => D(17), B2 => n95, ZN 
                           => n53);
   U23 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(18));
   U24 : AOI22_X1 port map( A1 => A(18), A2 => n90, B1 => B(18), B2 => n86, ZN 
                           => n50);
   U25 : AOI22_X1 port map( A1 => C(18), A2 => n99, B1 => D(18), B2 => n95, ZN 
                           => n51);
   U26 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(19));
   U27 : AOI22_X1 port map( A1 => A(19), A2 => n90, B1 => B(19), B2 => n86, ZN 
                           => n48);
   U28 : AOI22_X1 port map( A1 => C(19), A2 => n99, B1 => D(19), B2 => n95, ZN 
                           => n49);
   U29 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(20));
   U30 : AOI22_X1 port map( A1 => A(20), A2 => n91, B1 => B(20), B2 => n87, ZN 
                           => n44);
   U31 : AOI22_X1 port map( A1 => C(20), A2 => n100, B1 => D(20), B2 => n96, ZN
                           => n45);
   U32 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(21));
   U33 : AOI22_X1 port map( A1 => A(21), A2 => n91, B1 => B(21), B2 => n87, ZN 
                           => n42);
   U34 : AOI22_X1 port map( A1 => C(21), A2 => n100, B1 => D(21), B2 => n96, ZN
                           => n43);
   U35 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(22));
   U36 : AOI22_X1 port map( A1 => A(22), A2 => n91, B1 => B(22), B2 => n87, ZN 
                           => n40);
   U37 : AOI22_X1 port map( A1 => C(22), A2 => n100, B1 => D(22), B2 => n96, ZN
                           => n41);
   U38 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(23));
   U39 : AOI22_X1 port map( A1 => A(23), A2 => n91, B1 => B(23), B2 => n87, ZN 
                           => n38);
   U40 : AOI22_X1 port map( A1 => C(23), A2 => n100, B1 => D(23), B2 => n96, ZN
                           => n39);
   U41 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(24));
   U42 : AOI22_X1 port map( A1 => A(24), A2 => n91, B1 => B(24), B2 => n87, ZN 
                           => n36);
   U43 : AOI22_X1 port map( A1 => C(24), A2 => n100, B1 => D(24), B2 => n96, ZN
                           => n37);
   U44 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(25));
   U45 : AOI22_X1 port map( A1 => A(25), A2 => n91, B1 => B(25), B2 => n87, ZN 
                           => n34);
   U46 : AOI22_X1 port map( A1 => C(25), A2 => n100, B1 => D(25), B2 => n96, ZN
                           => n35);
   U47 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(26));
   U48 : AOI22_X1 port map( A1 => A(26), A2 => n91, B1 => B(26), B2 => n87, ZN 
                           => n32);
   U49 : AOI22_X1 port map( A1 => C(26), A2 => n100, B1 => D(26), B2 => n96, ZN
                           => n33);
   U50 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(27));
   U51 : AOI22_X1 port map( A1 => A(27), A2 => n91, B1 => B(27), B2 => n87, ZN 
                           => n30);
   U52 : AOI22_X1 port map( A1 => C(27), A2 => n100, B1 => D(27), B2 => n96, ZN
                           => n31);
   U53 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(28));
   U54 : AOI22_X1 port map( A1 => A(28), A2 => n91, B1 => B(28), B2 => n87, ZN 
                           => n28);
   U55 : AOI22_X1 port map( A1 => C(28), A2 => n100, B1 => D(28), B2 => n96, ZN
                           => n29);
   U56 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(29));
   U57 : AOI22_X1 port map( A1 => A(29), A2 => n91, B1 => B(29), B2 => n87, ZN 
                           => n26);
   U58 : AOI22_X1 port map( A1 => C(29), A2 => n100, B1 => D(29), B2 => n96, ZN
                           => n27);
   U59 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(30));
   U60 : AOI22_X1 port map( A1 => A(30), A2 => n91, B1 => B(30), B2 => n87, ZN 
                           => n22);
   U61 : AOI22_X1 port map( A1 => C(30), A2 => n100, B1 => D(30), B2 => n96, ZN
                           => n23);
   U62 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(31));
   U63 : AOI22_X1 port map( A1 => A(31), A2 => n92, B1 => B(31), B2 => n88, ZN 
                           => n20);
   U64 : AOI22_X1 port map( A1 => C(31), A2 => n101, B1 => D(31), B2 => n97, ZN
                           => n21);
   U65 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(0));
   U66 : AOI22_X1 port map( A1 => C(0), A2 => n99, B1 => D(0), B2 => n95, ZN =>
                           n69);
   U67 : AOI22_X1 port map( A1 => A(0), A2 => n90, B1 => B(0), B2 => n86, ZN =>
                           n68);
   U68 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(1));
   U69 : AOI22_X1 port map( A1 => C(1), A2 => n99, B1 => D(1), B2 => n95, ZN =>
                           n47);
   U70 : AOI22_X1 port map( A1 => A(1), A2 => n90, B1 => B(1), B2 => n86, ZN =>
                           n46);
   U71 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(2));
   U72 : AOI22_X1 port map( A1 => C(2), A2 => n100, B1 => D(2), B2 => n96, ZN 
                           => n25);
   U73 : AOI22_X1 port map( A1 => A(2), A2 => n91, B1 => B(2), B2 => n87, ZN =>
                           n24);
   U74 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(3));
   U75 : AOI22_X1 port map( A1 => C(3), A2 => n101, B1 => D(3), B2 => n97, ZN 
                           => n19);
   U76 : AOI22_X1 port map( A1 => A(3), A2 => n92, B1 => B(3), B2 => n88, ZN =>
                           n18);
   U77 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(4));
   U78 : AOI22_X1 port map( A1 => C(4), A2 => n101, B1 => D(4), B2 => n97, ZN 
                           => n17);
   U79 : AOI22_X1 port map( A1 => A(4), A2 => n92, B1 => B(4), B2 => n88, ZN =>
                           n16);
   U80 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(5));
   U81 : AOI22_X1 port map( A1 => C(5), A2 => n101, B1 => D(5), B2 => n97, ZN 
                           => n15);
   U82 : AOI22_X1 port map( A1 => A(5), A2 => n92, B1 => B(5), B2 => n88, ZN =>
                           n14);
   U83 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(6));
   U84 : AOI22_X1 port map( A1 => C(6), A2 => n101, B1 => D(6), B2 => n97, ZN 
                           => n13);
   U85 : AOI22_X1 port map( A1 => A(6), A2 => n92, B1 => B(6), B2 => n88, ZN =>
                           n12);
   U86 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(7));
   U87 : AOI22_X1 port map( A1 => C(7), A2 => n101, B1 => D(7), B2 => n97, ZN 
                           => n11);
   U88 : AOI22_X1 port map( A1 => A(7), A2 => n92, B1 => B(7), B2 => n88, ZN =>
                           n10);
   U89 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(8));
   U90 : AOI22_X1 port map( A1 => C(8), A2 => n101, B1 => D(8), B2 => n97, ZN 
                           => n9);
   U91 : AOI22_X1 port map( A1 => A(8), A2 => n92, B1 => B(8), B2 => n88, ZN =>
                           n8);
   U92 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(9));
   U93 : AOI22_X1 port map( A1 => C(9), A2 => n101, B1 => D(9), B2 => n97, ZN 
                           => n3);
   U94 : AOI22_X1 port map( A1 => A(9), A2 => n92, B1 => B(9), B2 => n88, ZN =>
                           n2);
   U95 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(10));
   U96 : AOI22_X1 port map( A1 => C(10), A2 => n99, B1 => D(10), B2 => n95, ZN 
                           => n67);
   U97 : AOI22_X1 port map( A1 => A(10), A2 => n90, B1 => B(10), B2 => n86, ZN 
                           => n66);
   U98 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(11));
   U99 : AOI22_X1 port map( A1 => C(11), A2 => n99, B1 => D(11), B2 => n95, ZN 
                           => n65);
   U100 : AOI22_X1 port map( A1 => A(11), A2 => n90, B1 => B(11), B2 => n86, ZN
                           => n64);
   U101 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(12));
   U102 : AOI22_X1 port map( A1 => C(12), A2 => n99, B1 => D(12), B2 => n95, ZN
                           => n63);
   U103 : AOI22_X1 port map( A1 => A(12), A2 => n90, B1 => B(12), B2 => n86, ZN
                           => n62);
   U104 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(13));
   U105 : AOI22_X1 port map( A1 => C(13), A2 => n99, B1 => D(13), B2 => n95, ZN
                           => n61);
   U106 : AOI22_X1 port map( A1 => A(13), A2 => n90, B1 => B(13), B2 => n86, ZN
                           => n60);
   U107 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(14));
   U108 : AOI22_X1 port map( A1 => C(14), A2 => n99, B1 => D(14), B2 => n95, ZN
                           => n59);
   U109 : AOI22_X1 port map( A1 => A(14), A2 => n90, B1 => B(14), B2 => n86, ZN
                           => n58);
   U110 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(15));
   U111 : AOI22_X1 port map( A1 => C(15), A2 => n99, B1 => D(15), B2 => n95, ZN
                           => n57);
   U112 : AOI22_X1 port map( A1 => A(15), A2 => n90, B1 => B(15), B2 => n86, ZN
                           => n56);
   U113 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n6);
   U114 : NOR2_X1 port map( A1 => n102, A2 => SEL(1), ZN => n7);
   U115 : INV_X1 port map( A => SEL(0), ZN => n102);
   U116 : AND2_X1 port map( A1 => SEL(1), A2 => n102, ZN => n4);
   U117 : AND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n5);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT2 is

   port( A, B, C, SEL : in std_logic_vector (1 downto 0);  Y : out 
         std_logic_vector (1 downto 0));

end MUX3to1_NBIT2;

architecture SYN_Behavioral of MUX3to1_NBIT2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, N13, N14, n2, n3, n4, n5, n6 : std_logic;

begin
   
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => N14, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => N13, Q => Y(0));
   U9 : NAND3_X1 port map( A1 => C(1), A2 => n6, A3 => SEL(1), ZN => n3);
   U10 : NAND3_X1 port map( A1 => SEL(1), A2 => n6, A3 => C(0), ZN => n5);
   U3 : INV_X1 port map( A => SEL(0), ZN => n6);
   U4 : NAND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => N12);
   U5 : OAI21_X1 port map( B1 => SEL(1), B2 => n4, A => n5, ZN => N13);
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n6, B1 => B(0), B2 => SEL(0), ZN 
                           => n4);
   U7 : OAI21_X1 port map( B1 => SEL(1), B2 => n2, A => n3, ZN => N14);
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n6, B1 => SEL(0), B2 => B(1), ZN 
                           => n2);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_3;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n105, n106, n107, n108, n109, n110, n111, n112 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n108, Z => n111);
   U2 : BUF_X1 port map( A => n108, Z => n112);
   U3 : INV_X1 port map( A => n111, ZN => n109);
   U4 : INV_X1 port map( A => n111, ZN => n110);
   U5 : BUF_X1 port map( A => n112, Z => n105);
   U6 : BUF_X1 port map( A => n112, Z => n106);
   U7 : BUF_X1 port map( A => n112, Z => n107);
   U8 : INV_X1 port map( A => n65, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n109, B1 => B(0), B2 => n105, ZN 
                           => n65);
   U10 : INV_X1 port map( A => n64, ZN => Y(1));
   U11 : AOI22_X1 port map( A1 => A(1), A2 => n109, B1 => B(1), B2 => n105, ZN 
                           => n64);
   U12 : INV_X1 port map( A => n63, ZN => Y(2));
   U13 : AOI22_X1 port map( A1 => A(2), A2 => n109, B1 => B(2), B2 => n105, ZN 
                           => n63);
   U14 : INV_X1 port map( A => n62, ZN => Y(3));
   U15 : AOI22_X1 port map( A1 => A(3), A2 => n109, B1 => B(3), B2 => n105, ZN 
                           => n62);
   U16 : INV_X1 port map( A => n61, ZN => Y(4));
   U17 : AOI22_X1 port map( A1 => A(4), A2 => n109, B1 => B(4), B2 => n105, ZN 
                           => n61);
   U18 : INV_X1 port map( A => n60, ZN => Y(5));
   U19 : AOI22_X1 port map( A1 => A(5), A2 => n109, B1 => B(5), B2 => n105, ZN 
                           => n60);
   U20 : INV_X1 port map( A => n59, ZN => Y(6));
   U21 : AOI22_X1 port map( A1 => A(6), A2 => n109, B1 => B(6), B2 => n105, ZN 
                           => n59);
   U22 : INV_X1 port map( A => n58, ZN => Y(7));
   U23 : AOI22_X1 port map( A1 => A(7), A2 => n109, B1 => B(7), B2 => n105, ZN 
                           => n58);
   U24 : INV_X1 port map( A => n57, ZN => Y(8));
   U25 : AOI22_X1 port map( A1 => A(8), A2 => n109, B1 => B(8), B2 => n105, ZN 
                           => n57);
   U26 : INV_X1 port map( A => n56, ZN => Y(9));
   U27 : AOI22_X1 port map( A1 => A(9), A2 => n109, B1 => B(9), B2 => n105, ZN 
                           => n56);
   U28 : INV_X1 port map( A => n55, ZN => Y(10));
   U29 : AOI22_X1 port map( A1 => A(10), A2 => n109, B1 => B(10), B2 => n105, 
                           ZN => n55);
   U30 : INV_X1 port map( A => n54, ZN => Y(11));
   U31 : AOI22_X1 port map( A1 => A(11), A2 => n109, B1 => B(11), B2 => n105, 
                           ZN => n54);
   U32 : INV_X1 port map( A => n53, ZN => Y(12));
   U33 : AOI22_X1 port map( A1 => A(12), A2 => n110, B1 => B(12), B2 => n106, 
                           ZN => n53);
   U34 : INV_X1 port map( A => n52, ZN => Y(13));
   U35 : AOI22_X1 port map( A1 => A(13), A2 => n110, B1 => B(13), B2 => n106, 
                           ZN => n52);
   U36 : INV_X1 port map( A => n51, ZN => Y(14));
   U37 : AOI22_X1 port map( A1 => A(14), A2 => n110, B1 => B(14), B2 => n106, 
                           ZN => n51);
   U38 : INV_X1 port map( A => n50, ZN => Y(15));
   U39 : AOI22_X1 port map( A1 => A(15), A2 => n110, B1 => B(15), B2 => n106, 
                           ZN => n50);
   U40 : INV_X1 port map( A => n49, ZN => Y(16));
   U41 : AOI22_X1 port map( A1 => A(16), A2 => n110, B1 => B(16), B2 => n106, 
                           ZN => n49);
   U42 : INV_X1 port map( A => n48, ZN => Y(17));
   U43 : AOI22_X1 port map( A1 => A(17), A2 => n110, B1 => B(17), B2 => n106, 
                           ZN => n48);
   U44 : INV_X1 port map( A => n47, ZN => Y(18));
   U45 : AOI22_X1 port map( A1 => A(18), A2 => n110, B1 => B(18), B2 => n106, 
                           ZN => n47);
   U46 : INV_X1 port map( A => n46, ZN => Y(19));
   U47 : AOI22_X1 port map( A1 => A(19), A2 => n110, B1 => B(19), B2 => n106, 
                           ZN => n46);
   U48 : INV_X1 port map( A => n45, ZN => Y(20));
   U49 : AOI22_X1 port map( A1 => A(20), A2 => n110, B1 => B(20), B2 => n106, 
                           ZN => n45);
   U50 : INV_X1 port map( A => n44, ZN => Y(21));
   U51 : AOI22_X1 port map( A1 => A(21), A2 => n110, B1 => B(21), B2 => n106, 
                           ZN => n44);
   U52 : INV_X1 port map( A => n43, ZN => Y(22));
   U53 : AOI22_X1 port map( A1 => A(22), A2 => n110, B1 => B(22), B2 => n106, 
                           ZN => n43);
   U54 : INV_X1 port map( A => n42, ZN => Y(23));
   U55 : AOI22_X1 port map( A1 => A(23), A2 => n110, B1 => B(23), B2 => n106, 
                           ZN => n42);
   U56 : INV_X1 port map( A => n41, ZN => Y(24));
   U57 : AOI22_X1 port map( A1 => A(24), A2 => n109, B1 => B(24), B2 => n107, 
                           ZN => n41);
   U58 : INV_X1 port map( A => n40, ZN => Y(25));
   U59 : AOI22_X1 port map( A1 => A(25), A2 => n110, B1 => B(25), B2 => n107, 
                           ZN => n40);
   U60 : INV_X1 port map( A => n39, ZN => Y(26));
   U61 : AOI22_X1 port map( A1 => A(26), A2 => n109, B1 => B(26), B2 => n107, 
                           ZN => n39);
   U62 : INV_X1 port map( A => n38, ZN => Y(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n110, B1 => B(27), B2 => n107, 
                           ZN => n38);
   U64 : INV_X1 port map( A => n37, ZN => Y(28));
   U65 : AOI22_X1 port map( A1 => A(28), A2 => n109, B1 => B(28), B2 => n107, 
                           ZN => n37);
   U66 : INV_X1 port map( A => n36, ZN => Y(29));
   U67 : AOI22_X1 port map( A1 => A(29), A2 => n110, B1 => B(29), B2 => n107, 
                           ZN => n36);
   U68 : INV_X1 port map( A => n35, ZN => Y(30));
   U69 : AOI22_X1 port map( A1 => A(30), A2 => n109, B1 => B(30), B2 => n107, 
                           ZN => n35);
   U70 : INV_X1 port map( A => n34, ZN => Y(31));
   U71 : AOI22_X1 port map( A1 => A(31), A2 => n110, B1 => n107, B2 => B(31), 
                           ZN => n34);
   U72 : BUF_X1 port map( A => SEL, Z => n108);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_0 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_0;

architecture SYN_Behavioral of MUX5to1_NBIT32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n118, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n118, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n118, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n118, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n118, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n118, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n118, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n118, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n118, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n118, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n117, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n119, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n119, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n119, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n119, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n119, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n119, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n119, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n119, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n119, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n119, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n118, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n117, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n117, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n117, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n117, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n117, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n117, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n117, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n117, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n117, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n117, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n120);
   U4 : BUF_X1 port map( A => n6, Z => n112);
   U5 : BUF_X1 port map( A => n7, Z => n108);
   U6 : BUF_X1 port map( A => n5, Z => n116);
   U7 : BUF_X1 port map( A => n8, Z => n104);
   U8 : BUF_X1 port map( A => n9, Z => n97);
   U9 : BUF_X1 port map( A => n120, Z => n117);
   U10 : BUF_X1 port map( A => n120, Z => n118);
   U11 : BUF_X1 port map( A => n120, Z => n119);
   U12 : OR4_X1 port map( A1 => n103, A2 => n100, A3 => n115, A4 => n72, ZN => 
                           N25);
   U13 : OR2_X1 port map( A1 => n107, A2 => n111, ZN => n72);
   U14 : BUF_X1 port map( A => n104, Z => n102);
   U15 : BUF_X1 port map( A => n104, Z => n101);
   U16 : BUF_X1 port map( A => n97, Z => n99);
   U17 : BUF_X1 port map( A => n97, Z => n98);
   U18 : BUF_X1 port map( A => n112, Z => n110);
   U19 : BUF_X1 port map( A => n112, Z => n109);
   U20 : BUF_X1 port map( A => n108, Z => n106);
   U21 : BUF_X1 port map( A => n108, Z => n105);
   U22 : BUF_X1 port map( A => n116, Z => n114);
   U23 : BUF_X1 port map( A => n116, Z => n113);
   U24 : BUF_X1 port map( A => n104, Z => n103);
   U25 : BUF_X1 port map( A => n97, Z => n100);
   U26 : BUF_X1 port map( A => n112, Z => n111);
   U27 : BUF_X1 port map( A => n108, Z => n107);
   U28 : BUF_X1 port map( A => n116, Z => n115);
   U29 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n122, ZN => n6);
   U30 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n121, ZN => n7);
   U31 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n5);
   U32 : NOR3_X1 port map( A1 => n122, A2 => SEL(2), A3 => n121, ZN => n8);
   U33 : AND3_X1 port map( A1 => n121, A2 => n122, A3 => SEL(2), ZN => n9);
   U34 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U35 : AOI22_X1 port map( A1 => D(0), A2 => n103, B1 => E(0), B2 => n100, ZN 
                           => n70);
   U36 : AOI222_X1 port map( A1 => A(0), A2 => n115, B1 => C(0), B2 => n111, C1
                           => B(0), C2 => n107, ZN => n71);
   U37 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U38 : AOI22_X1 port map( A1 => D(1), A2 => n103, B1 => E(1), B2 => n100, ZN 
                           => n68);
   U39 : AOI222_X1 port map( A1 => A(1), A2 => n115, B1 => C(1), B2 => n111, C1
                           => B(1), C2 => n107, ZN => n69);
   U40 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U41 : AOI22_X1 port map( A1 => D(2), A2 => n103, B1 => E(2), B2 => n100, ZN 
                           => n66);
   U42 : AOI222_X1 port map( A1 => A(2), A2 => n115, B1 => C(2), B2 => n111, C1
                           => B(2), C2 => n107, ZN => n67);
   U43 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U44 : AOI22_X1 port map( A1 => D(3), A2 => n103, B1 => E(3), B2 => n100, ZN 
                           => n64);
   U45 : AOI222_X1 port map( A1 => A(3), A2 => n115, B1 => C(3), B2 => n111, C1
                           => B(3), C2 => n107, ZN => n65);
   U46 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U47 : AOI22_X1 port map( A1 => D(4), A2 => n103, B1 => E(4), B2 => n100, ZN 
                           => n62);
   U48 : AOI222_X1 port map( A1 => A(4), A2 => n115, B1 => C(4), B2 => n111, C1
                           => B(4), C2 => n107, ZN => n63);
   U49 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U50 : AOI22_X1 port map( A1 => D(5), A2 => n103, B1 => E(5), B2 => n100, ZN 
                           => n60);
   U51 : AOI222_X1 port map( A1 => A(5), A2 => n115, B1 => C(5), B2 => n111, C1
                           => B(5), C2 => n107, ZN => n61);
   U52 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U53 : AOI22_X1 port map( A1 => D(6), A2 => n103, B1 => E(6), B2 => n100, ZN 
                           => n58);
   U54 : AOI222_X1 port map( A1 => A(6), A2 => n115, B1 => C(6), B2 => n111, C1
                           => B(6), C2 => n107, ZN => n59);
   U55 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U56 : AOI22_X1 port map( A1 => D(7), A2 => n103, B1 => E(7), B2 => n100, ZN 
                           => n56_port);
   U57 : AOI222_X1 port map( A1 => A(7), A2 => n115, B1 => C(7), B2 => n111, C1
                           => B(7), C2 => n107, ZN => n57_port);
   U58 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U59 : AOI22_X1 port map( A1 => D(8), A2 => n102, B1 => E(8), B2 => n99, ZN 
                           => n54_port);
   U60 : AOI222_X1 port map( A1 => A(8), A2 => n114, B1 => C(8), B2 => n110, C1
                           => B(8), C2 => n106, ZN => n55_port);
   U61 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U62 : AOI22_X1 port map( A1 => D(9), A2 => n102, B1 => E(9), B2 => n99, ZN 
                           => n52_port);
   U63 : AOI222_X1 port map( A1 => A(9), A2 => n114, B1 => C(9), B2 => n110, C1
                           => B(9), C2 => n106, ZN => n53_port);
   U64 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U65 : AOI22_X1 port map( A1 => D(10), A2 => n102, B1 => E(10), B2 => n99, ZN
                           => n50_port);
   U66 : AOI222_X1 port map( A1 => A(10), A2 => n114, B1 => C(10), B2 => n110, 
                           C1 => B(10), C2 => n106, ZN => n51_port);
   U67 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U68 : AOI22_X1 port map( A1 => D(11), A2 => n102, B1 => E(11), B2 => n99, ZN
                           => n48_port);
   U69 : AOI222_X1 port map( A1 => A(11), A2 => n114, B1 => C(11), B2 => n110, 
                           C1 => B(11), C2 => n106, ZN => n49_port);
   U70 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U71 : AOI22_X1 port map( A1 => D(12), A2 => n102, B1 => E(12), B2 => n99, ZN
                           => n46_port);
   U72 : AOI222_X1 port map( A1 => A(12), A2 => n114, B1 => C(12), B2 => n110, 
                           C1 => B(12), C2 => n106, ZN => n47_port);
   U73 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U74 : AOI22_X1 port map( A1 => D(13), A2 => n102, B1 => E(13), B2 => n99, ZN
                           => n44_port);
   U75 : AOI222_X1 port map( A1 => A(13), A2 => n114, B1 => C(13), B2 => n110, 
                           C1 => B(13), C2 => n106, ZN => n45_port);
   U76 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U77 : AOI22_X1 port map( A1 => D(14), A2 => n102, B1 => E(14), B2 => n99, ZN
                           => n42_port);
   U78 : AOI222_X1 port map( A1 => A(14), A2 => n114, B1 => C(14), B2 => n110, 
                           C1 => B(14), C2 => n106, ZN => n43_port);
   U79 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U80 : AOI22_X1 port map( A1 => D(15), A2 => n102, B1 => E(15), B2 => n99, ZN
                           => n40_port);
   U81 : AOI222_X1 port map( A1 => A(15), A2 => n114, B1 => C(15), B2 => n110, 
                           C1 => B(15), C2 => n106, ZN => n41_port);
   U82 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U83 : AOI22_X1 port map( A1 => D(16), A2 => n102, B1 => E(16), B2 => n99, ZN
                           => n38_port);
   U84 : AOI222_X1 port map( A1 => A(16), A2 => n114, B1 => C(16), B2 => n110, 
                           C1 => B(16), C2 => n106, ZN => n39_port);
   U85 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U86 : AOI22_X1 port map( A1 => D(17), A2 => n102, B1 => E(17), B2 => n99, ZN
                           => n36_port);
   U87 : AOI222_X1 port map( A1 => A(17), A2 => n114, B1 => C(17), B2 => n110, 
                           C1 => B(17), C2 => n106, ZN => n37_port);
   U88 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U89 : AOI22_X1 port map( A1 => D(18), A2 => n102, B1 => E(18), B2 => n99, ZN
                           => n34_port);
   U90 : AOI222_X1 port map( A1 => A(18), A2 => n114, B1 => C(18), B2 => n110, 
                           C1 => B(18), C2 => n106, ZN => n35_port);
   U91 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U92 : AOI22_X1 port map( A1 => D(19), A2 => n102, B1 => E(19), B2 => n99, ZN
                           => n32_port);
   U93 : AOI222_X1 port map( A1 => A(19), A2 => n114, B1 => C(19), B2 => n110, 
                           C1 => B(19), C2 => n106, ZN => n33_port);
   U94 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U95 : AOI22_X1 port map( A1 => D(20), A2 => n101, B1 => E(20), B2 => n98, ZN
                           => n30_port);
   U96 : AOI222_X1 port map( A1 => A(20), A2 => n113, B1 => C(20), B2 => n109, 
                           C1 => B(20), C2 => n105, ZN => n31_port);
   U97 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U98 : AOI22_X1 port map( A1 => D(21), A2 => n101, B1 => E(21), B2 => n98, ZN
                           => n28_port);
   U99 : AOI222_X1 port map( A1 => A(21), A2 => n113, B1 => C(21), B2 => n109, 
                           C1 => B(21), C2 => n105, ZN => n29_port);
   U100 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U101 : AOI22_X1 port map( A1 => D(22), A2 => n101, B1 => E(22), B2 => n98, 
                           ZN => n26_port);
   U102 : AOI222_X1 port map( A1 => A(22), A2 => n113, B1 => C(22), B2 => n109,
                           C1 => B(22), C2 => n105, ZN => n27_port);
   U103 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U104 : AOI22_X1 port map( A1 => D(23), A2 => n101, B1 => E(23), B2 => n98, 
                           ZN => n24);
   U105 : AOI222_X1 port map( A1 => A(23), A2 => n113, B1 => C(23), B2 => n109,
                           C1 => B(23), C2 => n105, ZN => n25_port);
   U106 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U107 : AOI22_X1 port map( A1 => D(24), A2 => n101, B1 => E(24), B2 => n98, 
                           ZN => n22);
   U108 : AOI222_X1 port map( A1 => A(24), A2 => n113, B1 => C(24), B2 => n109,
                           C1 => B(24), C2 => n105, ZN => n23);
   U109 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U110 : AOI22_X1 port map( A1 => D(25), A2 => n101, B1 => E(25), B2 => n98, 
                           ZN => n20);
   U111 : AOI222_X1 port map( A1 => A(25), A2 => n113, B1 => C(25), B2 => n109,
                           C1 => B(25), C2 => n105, ZN => n21);
   U112 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U113 : AOI22_X1 port map( A1 => D(26), A2 => n101, B1 => E(26), B2 => n98, 
                           ZN => n18);
   U114 : AOI222_X1 port map( A1 => A(26), A2 => n113, B1 => C(26), B2 => n109,
                           C1 => B(26), C2 => n105, ZN => n19);
   U115 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U116 : AOI22_X1 port map( A1 => D(27), A2 => n101, B1 => E(27), B2 => n98, 
                           ZN => n16);
   U117 : AOI222_X1 port map( A1 => A(27), A2 => n113, B1 => C(27), B2 => n109,
                           C1 => B(27), C2 => n105, ZN => n17);
   U118 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U119 : AOI22_X1 port map( A1 => D(28), A2 => n101, B1 => E(28), B2 => n98, 
                           ZN => n14);
   U120 : AOI222_X1 port map( A1 => A(28), A2 => n113, B1 => C(28), B2 => n109,
                           C1 => B(28), C2 => n105, ZN => n15);
   U121 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U122 : AOI22_X1 port map( A1 => D(29), A2 => n101, B1 => E(29), B2 => n98, 
                           ZN => n12);
   U123 : AOI222_X1 port map( A1 => A(29), A2 => n113, B1 => C(29), B2 => n109,
                           C1 => B(29), C2 => n105, ZN => n13);
   U124 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U125 : AOI22_X1 port map( A1 => D(30), A2 => n101, B1 => E(30), B2 => n98, 
                           ZN => n10);
   U126 : AOI222_X1 port map( A1 => A(30), A2 => n113, B1 => C(30), B2 => n109,
                           C1 => B(30), C2 => n105, ZN => n11);
   U127 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U128 : AOI22_X1 port map( A1 => D(31), A2 => n101, B1 => E(31), B2 => n98, 
                           ZN => n3);
   U129 : AOI222_X1 port map( A1 => A(31), A2 => n113, B1 => C(31), B2 => n109,
                           C1 => B(31), C2 => n105, ZN => n4);
   U130 : INV_X1 port map( A => SEL(0), ZN => n121);
   U131 : INV_X1 port map( A => SEL(1), ZN => n122);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_4;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n105, n106, n107, n108, n109, n110, n111, n112 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n108, Z => n111);
   U2 : BUF_X1 port map( A => n108, Z => n112);
   U3 : INV_X1 port map( A => n111, ZN => n109);
   U4 : INV_X1 port map( A => n111, ZN => n110);
   U5 : BUF_X1 port map( A => n112, Z => n105);
   U6 : BUF_X1 port map( A => n112, Z => n106);
   U7 : BUF_X1 port map( A => n112, Z => n107);
   U8 : INV_X1 port map( A => n65, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n109, B1 => B(0), B2 => n105, ZN 
                           => n65);
   U10 : INV_X1 port map( A => n64, ZN => Y(1));
   U11 : AOI22_X1 port map( A1 => A(1), A2 => n109, B1 => B(1), B2 => n105, ZN 
                           => n64);
   U12 : INV_X1 port map( A => n63, ZN => Y(2));
   U13 : AOI22_X1 port map( A1 => A(2), A2 => n109, B1 => B(2), B2 => n105, ZN 
                           => n63);
   U14 : INV_X1 port map( A => n62, ZN => Y(3));
   U15 : AOI22_X1 port map( A1 => A(3), A2 => n109, B1 => B(3), B2 => n105, ZN 
                           => n62);
   U16 : INV_X1 port map( A => n61, ZN => Y(4));
   U17 : AOI22_X1 port map( A1 => A(4), A2 => n109, B1 => B(4), B2 => n105, ZN 
                           => n61);
   U18 : INV_X1 port map( A => n60, ZN => Y(5));
   U19 : AOI22_X1 port map( A1 => A(5), A2 => n109, B1 => B(5), B2 => n105, ZN 
                           => n60);
   U20 : INV_X1 port map( A => n59, ZN => Y(6));
   U21 : AOI22_X1 port map( A1 => A(6), A2 => n109, B1 => B(6), B2 => n105, ZN 
                           => n59);
   U22 : INV_X1 port map( A => n58, ZN => Y(7));
   U23 : AOI22_X1 port map( A1 => A(7), A2 => n109, B1 => B(7), B2 => n105, ZN 
                           => n58);
   U24 : INV_X1 port map( A => n57, ZN => Y(8));
   U25 : AOI22_X1 port map( A1 => A(8), A2 => n109, B1 => B(8), B2 => n105, ZN 
                           => n57);
   U26 : INV_X1 port map( A => n56, ZN => Y(9));
   U27 : AOI22_X1 port map( A1 => A(9), A2 => n109, B1 => B(9), B2 => n105, ZN 
                           => n56);
   U28 : INV_X1 port map( A => n55, ZN => Y(10));
   U29 : AOI22_X1 port map( A1 => A(10), A2 => n109, B1 => B(10), B2 => n105, 
                           ZN => n55);
   U30 : INV_X1 port map( A => n54, ZN => Y(11));
   U31 : AOI22_X1 port map( A1 => A(11), A2 => n109, B1 => B(11), B2 => n105, 
                           ZN => n54);
   U32 : INV_X1 port map( A => n53, ZN => Y(12));
   U33 : AOI22_X1 port map( A1 => A(12), A2 => n110, B1 => B(12), B2 => n106, 
                           ZN => n53);
   U34 : INV_X1 port map( A => n52, ZN => Y(13));
   U35 : AOI22_X1 port map( A1 => A(13), A2 => n110, B1 => B(13), B2 => n106, 
                           ZN => n52);
   U36 : INV_X1 port map( A => n51, ZN => Y(14));
   U37 : AOI22_X1 port map( A1 => A(14), A2 => n110, B1 => B(14), B2 => n106, 
                           ZN => n51);
   U38 : INV_X1 port map( A => n50, ZN => Y(15));
   U39 : AOI22_X1 port map( A1 => A(15), A2 => n110, B1 => B(15), B2 => n106, 
                           ZN => n50);
   U40 : INV_X1 port map( A => n49, ZN => Y(16));
   U41 : AOI22_X1 port map( A1 => A(16), A2 => n110, B1 => B(16), B2 => n106, 
                           ZN => n49);
   U42 : INV_X1 port map( A => n48, ZN => Y(17));
   U43 : AOI22_X1 port map( A1 => A(17), A2 => n110, B1 => B(17), B2 => n106, 
                           ZN => n48);
   U44 : INV_X1 port map( A => n47, ZN => Y(18));
   U45 : AOI22_X1 port map( A1 => A(18), A2 => n110, B1 => B(18), B2 => n106, 
                           ZN => n47);
   U46 : INV_X1 port map( A => n46, ZN => Y(19));
   U47 : AOI22_X1 port map( A1 => A(19), A2 => n110, B1 => B(19), B2 => n106, 
                           ZN => n46);
   U48 : INV_X1 port map( A => n45, ZN => Y(20));
   U49 : AOI22_X1 port map( A1 => A(20), A2 => n110, B1 => B(20), B2 => n106, 
                           ZN => n45);
   U50 : INV_X1 port map( A => n44, ZN => Y(21));
   U51 : AOI22_X1 port map( A1 => A(21), A2 => n110, B1 => B(21), B2 => n106, 
                           ZN => n44);
   U52 : INV_X1 port map( A => n43, ZN => Y(22));
   U53 : AOI22_X1 port map( A1 => A(22), A2 => n110, B1 => B(22), B2 => n106, 
                           ZN => n43);
   U54 : INV_X1 port map( A => n42, ZN => Y(23));
   U55 : AOI22_X1 port map( A1 => A(23), A2 => n110, B1 => B(23), B2 => n106, 
                           ZN => n42);
   U56 : INV_X1 port map( A => n41, ZN => Y(24));
   U57 : AOI22_X1 port map( A1 => A(24), A2 => n109, B1 => B(24), B2 => n107, 
                           ZN => n41);
   U58 : INV_X1 port map( A => n40, ZN => Y(25));
   U59 : AOI22_X1 port map( A1 => A(25), A2 => n110, B1 => B(25), B2 => n107, 
                           ZN => n40);
   U60 : INV_X1 port map( A => n39, ZN => Y(26));
   U61 : AOI22_X1 port map( A1 => A(26), A2 => n109, B1 => B(26), B2 => n107, 
                           ZN => n39);
   U62 : INV_X1 port map( A => n38, ZN => Y(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n110, B1 => B(27), B2 => n107, 
                           ZN => n38);
   U64 : INV_X1 port map( A => n37, ZN => Y(28));
   U65 : AOI22_X1 port map( A1 => A(28), A2 => n109, B1 => B(28), B2 => n107, 
                           ZN => n37);
   U66 : INV_X1 port map( A => n36, ZN => Y(29));
   U67 : AOI22_X1 port map( A1 => A(29), A2 => n110, B1 => B(29), B2 => n107, 
                           ZN => n36);
   U68 : INV_X1 port map( A => n35, ZN => Y(30));
   U69 : AOI22_X1 port map( A1 => A(30), A2 => n109, B1 => B(30), B2 => n107, 
                           ZN => n35);
   U70 : INV_X1 port map( A => n34, ZN => Y(31));
   U71 : AOI22_X1 port map( A1 => A(31), A2 => n110, B1 => n107, B2 => B(31), 
                           ZN => n34);
   U72 : BUF_X1 port map( A => SEL, Z => n108);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_1 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_1;

architecture SYN_Behavioral of MUX3to1_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n131, D => n134, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n132, D => n135, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n132, D => n136, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n132, D => n137, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n132, D => n138, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n132, D => n139, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n132, D => n140, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n132, D => n141, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n132, D => n142, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n132, D => n143, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n132, D => n144, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n133, D => n145, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n132, D => n146, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n133, D => n147, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n133, D => n148, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n133, D => n149, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n133, D => n150, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n133, D => n151, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n133, D => n152, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n133, D => n153, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n133, D => n154, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n133, D => n155, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n131, D => n156, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n131, D => n157, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n131, D => n158, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n131, D => n159, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n131, D => n160, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n131, D => n161, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n131, D => n162, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n131, D => n163, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n131, D => n164, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n131, D => n165, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n119, A2 => n128, A3 => n125, ZN => N12);
   U4 : BUF_X1 port map( A => n37, Z => n122);
   U5 : BUF_X1 port map( A => n36, Z => n126);
   U6 : BUF_X1 port map( A => n35, Z => n127);
   U7 : BUF_X1 port map( A => N12, Z => n132);
   U8 : BUF_X1 port map( A => N12, Z => n131);
   U9 : BUF_X1 port map( A => N12, Z => n133);
   U10 : BUF_X1 port map( A => n126, Z => n124);
   U11 : BUF_X1 port map( A => n126, Z => n123);
   U12 : BUF_X1 port map( A => n122, Z => n119);
   U13 : BUF_X1 port map( A => n122, Z => n120);
   U14 : BUF_X1 port map( A => n127, Z => n128);
   U15 : BUF_X1 port map( A => n127, Z => n129);
   U16 : BUF_X1 port map( A => n126, Z => n125);
   U17 : BUF_X1 port map( A => n122, Z => n121);
   U18 : BUF_X1 port map( A => n127, Z => n130);
   U19 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n37);
   U20 : NOR2_X1 port map( A1 => n166, A2 => SEL(0), ZN => n36);
   U21 : AND2_X1 port map( A1 => SEL(0), A2 => n166, ZN => n35);
   U22 : INV_X1 port map( A => SEL(1), ZN => n166);
   U23 : INV_X1 port map( A => n68, ZN => n165);
   U24 : AOI222_X1 port map( A1 => B(0), A2 => n128, B1 => C(0), B2 => n125, C1
                           => A(0), C2 => n119, ZN => n68);
   U25 : INV_X1 port map( A => n67, ZN => n164);
   U26 : AOI222_X1 port map( A1 => B(1), A2 => n128, B1 => C(1), B2 => n125, C1
                           => A(1), C2 => n119, ZN => n67);
   U27 : INV_X1 port map( A => n66, ZN => n163);
   U28 : AOI222_X1 port map( A1 => B(2), A2 => n128, B1 => C(2), B2 => n125, C1
                           => A(2), C2 => n119, ZN => n66);
   U29 : INV_X1 port map( A => n65, ZN => n162);
   U30 : AOI222_X1 port map( A1 => B(3), A2 => n128, B1 => C(3), B2 => n125, C1
                           => A(3), C2 => n119, ZN => n65);
   U31 : INV_X1 port map( A => n64, ZN => n161);
   U32 : AOI222_X1 port map( A1 => B(4), A2 => n128, B1 => C(4), B2 => n125, C1
                           => A(4), C2 => n119, ZN => n64);
   U33 : INV_X1 port map( A => n63, ZN => n160);
   U34 : AOI222_X1 port map( A1 => B(5), A2 => n128, B1 => C(5), B2 => n125, C1
                           => A(5), C2 => n119, ZN => n63);
   U35 : INV_X1 port map( A => n62, ZN => n159);
   U36 : AOI222_X1 port map( A1 => B(6), A2 => n128, B1 => C(6), B2 => n125, C1
                           => A(6), C2 => n119, ZN => n62);
   U37 : INV_X1 port map( A => n61, ZN => n158);
   U38 : AOI222_X1 port map( A1 => B(7), A2 => n128, B1 => C(7), B2 => n125, C1
                           => A(7), C2 => n119, ZN => n61);
   U39 : INV_X1 port map( A => n60, ZN => n157);
   U40 : AOI222_X1 port map( A1 => B(8), A2 => n128, B1 => C(8), B2 => n124, C1
                           => A(8), C2 => n119, ZN => n60);
   U41 : INV_X1 port map( A => n59, ZN => n156);
   U42 : AOI222_X1 port map( A1 => B(9), A2 => n128, B1 => C(9), B2 => n124, C1
                           => A(9), C2 => n119, ZN => n59);
   U43 : INV_X1 port map( A => n58, ZN => n155);
   U44 : AOI222_X1 port map( A1 => B(10), A2 => n128, B1 => C(10), B2 => n124, 
                           C1 => A(10), C2 => n119, ZN => n58);
   U45 : INV_X1 port map( A => n57, ZN => n154);
   U46 : AOI222_X1 port map( A1 => B(11), A2 => n129, B1 => C(11), B2 => n124, 
                           C1 => A(11), C2 => n120, ZN => n57);
   U47 : INV_X1 port map( A => n56, ZN => n153);
   U48 : AOI222_X1 port map( A1 => B(12), A2 => n129, B1 => C(12), B2 => n124, 
                           C1 => A(12), C2 => n120, ZN => n56);
   U49 : INV_X1 port map( A => n55, ZN => n152);
   U50 : AOI222_X1 port map( A1 => B(13), A2 => n129, B1 => C(13), B2 => n124, 
                           C1 => A(13), C2 => n120, ZN => n55);
   U51 : INV_X1 port map( A => n54, ZN => n151);
   U52 : AOI222_X1 port map( A1 => B(14), A2 => n129, B1 => C(14), B2 => n124, 
                           C1 => A(14), C2 => n120, ZN => n54);
   U53 : INV_X1 port map( A => n53, ZN => n150);
   U54 : AOI222_X1 port map( A1 => B(15), A2 => n129, B1 => C(15), B2 => n124, 
                           C1 => A(15), C2 => n120, ZN => n53);
   U55 : INV_X1 port map( A => n52, ZN => n149);
   U56 : AOI222_X1 port map( A1 => B(16), A2 => n129, B1 => C(16), B2 => n124, 
                           C1 => A(16), C2 => n120, ZN => n52);
   U57 : INV_X1 port map( A => n51, ZN => n148);
   U58 : AOI222_X1 port map( A1 => B(17), A2 => n129, B1 => C(17), B2 => n124, 
                           C1 => A(17), C2 => n120, ZN => n51);
   U59 : INV_X1 port map( A => n50, ZN => n147);
   U60 : AOI222_X1 port map( A1 => B(18), A2 => n129, B1 => C(18), B2 => n124, 
                           C1 => A(18), C2 => n120, ZN => n50);
   U61 : INV_X1 port map( A => n49, ZN => n146);
   U62 : AOI222_X1 port map( A1 => B(19), A2 => n129, B1 => C(19), B2 => n124, 
                           C1 => A(19), C2 => n120, ZN => n49);
   U63 : INV_X1 port map( A => n48, ZN => n145);
   U64 : AOI222_X1 port map( A1 => B(20), A2 => n129, B1 => C(20), B2 => n123, 
                           C1 => A(20), C2 => n120, ZN => n48);
   U65 : INV_X1 port map( A => n47, ZN => n144);
   U66 : AOI222_X1 port map( A1 => B(21), A2 => n129, B1 => C(21), B2 => n123, 
                           C1 => A(21), C2 => n120, ZN => n47);
   U67 : INV_X1 port map( A => n46, ZN => n143);
   U68 : AOI222_X1 port map( A1 => B(22), A2 => n129, B1 => C(22), B2 => n123, 
                           C1 => A(22), C2 => n120, ZN => n46);
   U69 : INV_X1 port map( A => n45, ZN => n142);
   U70 : AOI222_X1 port map( A1 => B(23), A2 => n130, B1 => C(23), B2 => n123, 
                           C1 => A(23), C2 => n121, ZN => n45);
   U71 : INV_X1 port map( A => n44, ZN => n141);
   U72 : AOI222_X1 port map( A1 => B(24), A2 => n130, B1 => C(24), B2 => n123, 
                           C1 => A(24), C2 => n121, ZN => n44);
   U73 : INV_X1 port map( A => n43, ZN => n140);
   U74 : AOI222_X1 port map( A1 => B(25), A2 => n130, B1 => C(25), B2 => n123, 
                           C1 => A(25), C2 => n121, ZN => n43);
   U75 : INV_X1 port map( A => n42, ZN => n139);
   U76 : AOI222_X1 port map( A1 => B(26), A2 => n130, B1 => C(26), B2 => n123, 
                           C1 => A(26), C2 => n121, ZN => n42);
   U77 : INV_X1 port map( A => n41, ZN => n138);
   U78 : AOI222_X1 port map( A1 => B(27), A2 => n130, B1 => C(27), B2 => n123, 
                           C1 => A(27), C2 => n121, ZN => n41);
   U79 : INV_X1 port map( A => n40, ZN => n137);
   U80 : AOI222_X1 port map( A1 => B(28), A2 => n130, B1 => C(28), B2 => n123, 
                           C1 => A(28), C2 => n121, ZN => n40);
   U81 : INV_X1 port map( A => n39, ZN => n136);
   U82 : AOI222_X1 port map( A1 => B(29), A2 => n130, B1 => C(29), B2 => n123, 
                           C1 => A(29), C2 => n121, ZN => n39);
   U83 : INV_X1 port map( A => n38, ZN => n135);
   U84 : AOI222_X1 port map( A1 => B(30), A2 => n130, B1 => C(30), B2 => n123, 
                           C1 => A(30), C2 => n121, ZN => n38);
   U85 : INV_X1 port map( A => n34, ZN => n134);
   U86 : AOI222_X1 port map( A1 => B(31), A2 => n130, B1 => C(31), B2 => n123, 
                           C1 => A(31), C2 => n121, ZN => n34);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_2 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_2;

architecture SYN_Behavioral of MUX3to1_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n132, D => n134, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n132, D => n135, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n132, D => n136, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n131, D => n137, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n132, D => n138, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n132, D => n139, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n132, D => n140, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n132, D => n141, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n132, D => n142, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n132, D => n143, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n132, D => n144, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n133, D => n145, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n133, D => n146, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n132, D => n147, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n133, D => n148, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n133, D => n149, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n133, D => n150, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n133, D => n151, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n133, D => n152, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n133, D => n153, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n133, D => n154, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n133, D => n155, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n131, D => n156, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n131, D => n157, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n131, D => n158, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n131, D => n159, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n131, D => n160, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n131, D => n161, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n131, D => n162, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n131, D => n163, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n131, D => n164, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n131, D => n165, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n119, A2 => n128, A3 => n125, ZN => N12);
   U4 : BUF_X1 port map( A => n37, Z => n122);
   U5 : BUF_X1 port map( A => n36, Z => n126);
   U6 : BUF_X1 port map( A => n35, Z => n127);
   U7 : BUF_X1 port map( A => N12, Z => n131);
   U8 : BUF_X1 port map( A => N12, Z => n132);
   U9 : BUF_X1 port map( A => N12, Z => n133);
   U10 : BUF_X1 port map( A => n126, Z => n124);
   U11 : BUF_X1 port map( A => n126, Z => n123);
   U12 : BUF_X1 port map( A => n122, Z => n119);
   U13 : BUF_X1 port map( A => n122, Z => n120);
   U14 : BUF_X1 port map( A => n127, Z => n128);
   U15 : BUF_X1 port map( A => n127, Z => n129);
   U16 : BUF_X1 port map( A => n126, Z => n125);
   U17 : BUF_X1 port map( A => n122, Z => n121);
   U18 : BUF_X1 port map( A => n127, Z => n130);
   U19 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n37);
   U20 : NOR2_X1 port map( A1 => n166, A2 => SEL(0), ZN => n36);
   U21 : AND2_X1 port map( A1 => SEL(0), A2 => n166, ZN => n35);
   U22 : INV_X1 port map( A => SEL(1), ZN => n166);
   U23 : INV_X1 port map( A => n68, ZN => n165);
   U24 : AOI222_X1 port map( A1 => B(0), A2 => n128, B1 => C(0), B2 => n125, C1
                           => A(0), C2 => n119, ZN => n68);
   U25 : INV_X1 port map( A => n67, ZN => n164);
   U26 : AOI222_X1 port map( A1 => B(1), A2 => n128, B1 => C(1), B2 => n125, C1
                           => A(1), C2 => n119, ZN => n67);
   U27 : INV_X1 port map( A => n66, ZN => n163);
   U28 : AOI222_X1 port map( A1 => B(2), A2 => n128, B1 => C(2), B2 => n125, C1
                           => A(2), C2 => n119, ZN => n66);
   U29 : INV_X1 port map( A => n65, ZN => n162);
   U30 : AOI222_X1 port map( A1 => B(3), A2 => n128, B1 => C(3), B2 => n125, C1
                           => A(3), C2 => n119, ZN => n65);
   U31 : INV_X1 port map( A => n64, ZN => n161);
   U32 : AOI222_X1 port map( A1 => B(4), A2 => n128, B1 => C(4), B2 => n125, C1
                           => A(4), C2 => n119, ZN => n64);
   U33 : INV_X1 port map( A => n63, ZN => n160);
   U34 : AOI222_X1 port map( A1 => B(5), A2 => n128, B1 => C(5), B2 => n125, C1
                           => A(5), C2 => n119, ZN => n63);
   U35 : INV_X1 port map( A => n62, ZN => n159);
   U36 : AOI222_X1 port map( A1 => B(6), A2 => n128, B1 => C(6), B2 => n125, C1
                           => A(6), C2 => n119, ZN => n62);
   U37 : INV_X1 port map( A => n61, ZN => n158);
   U38 : AOI222_X1 port map( A1 => B(7), A2 => n128, B1 => C(7), B2 => n125, C1
                           => A(7), C2 => n119, ZN => n61);
   U39 : INV_X1 port map( A => n60, ZN => n157);
   U40 : AOI222_X1 port map( A1 => B(8), A2 => n128, B1 => C(8), B2 => n124, C1
                           => A(8), C2 => n119, ZN => n60);
   U41 : INV_X1 port map( A => n59, ZN => n156);
   U42 : AOI222_X1 port map( A1 => B(9), A2 => n128, B1 => C(9), B2 => n124, C1
                           => A(9), C2 => n119, ZN => n59);
   U43 : INV_X1 port map( A => n58, ZN => n155);
   U44 : AOI222_X1 port map( A1 => B(10), A2 => n128, B1 => C(10), B2 => n124, 
                           C1 => A(10), C2 => n119, ZN => n58);
   U45 : INV_X1 port map( A => n57, ZN => n154);
   U46 : AOI222_X1 port map( A1 => B(11), A2 => n129, B1 => C(11), B2 => n124, 
                           C1 => A(11), C2 => n120, ZN => n57);
   U47 : INV_X1 port map( A => n56, ZN => n153);
   U48 : AOI222_X1 port map( A1 => B(12), A2 => n129, B1 => C(12), B2 => n124, 
                           C1 => A(12), C2 => n120, ZN => n56);
   U49 : INV_X1 port map( A => n55, ZN => n152);
   U50 : AOI222_X1 port map( A1 => B(13), A2 => n129, B1 => C(13), B2 => n124, 
                           C1 => A(13), C2 => n120, ZN => n55);
   U51 : INV_X1 port map( A => n54, ZN => n151);
   U52 : AOI222_X1 port map( A1 => B(14), A2 => n129, B1 => C(14), B2 => n124, 
                           C1 => A(14), C2 => n120, ZN => n54);
   U53 : INV_X1 port map( A => n53, ZN => n150);
   U54 : AOI222_X1 port map( A1 => B(15), A2 => n129, B1 => C(15), B2 => n124, 
                           C1 => A(15), C2 => n120, ZN => n53);
   U55 : INV_X1 port map( A => n52, ZN => n149);
   U56 : AOI222_X1 port map( A1 => B(16), A2 => n129, B1 => C(16), B2 => n124, 
                           C1 => A(16), C2 => n120, ZN => n52);
   U57 : INV_X1 port map( A => n51, ZN => n148);
   U58 : AOI222_X1 port map( A1 => B(17), A2 => n129, B1 => C(17), B2 => n124, 
                           C1 => A(17), C2 => n120, ZN => n51);
   U59 : INV_X1 port map( A => n50, ZN => n147);
   U60 : AOI222_X1 port map( A1 => B(18), A2 => n129, B1 => C(18), B2 => n124, 
                           C1 => A(18), C2 => n120, ZN => n50);
   U61 : INV_X1 port map( A => n49, ZN => n146);
   U62 : AOI222_X1 port map( A1 => B(19), A2 => n129, B1 => C(19), B2 => n124, 
                           C1 => A(19), C2 => n120, ZN => n49);
   U63 : INV_X1 port map( A => n48, ZN => n145);
   U64 : AOI222_X1 port map( A1 => B(20), A2 => n129, B1 => C(20), B2 => n123, 
                           C1 => A(20), C2 => n120, ZN => n48);
   U65 : INV_X1 port map( A => n47, ZN => n144);
   U66 : AOI222_X1 port map( A1 => B(21), A2 => n129, B1 => C(21), B2 => n123, 
                           C1 => A(21), C2 => n120, ZN => n47);
   U67 : INV_X1 port map( A => n46, ZN => n143);
   U68 : AOI222_X1 port map( A1 => B(22), A2 => n129, B1 => C(22), B2 => n123, 
                           C1 => A(22), C2 => n120, ZN => n46);
   U69 : INV_X1 port map( A => n45, ZN => n142);
   U70 : AOI222_X1 port map( A1 => B(23), A2 => n130, B1 => C(23), B2 => n123, 
                           C1 => A(23), C2 => n121, ZN => n45);
   U71 : INV_X1 port map( A => n44, ZN => n141);
   U72 : AOI222_X1 port map( A1 => B(24), A2 => n130, B1 => C(24), B2 => n123, 
                           C1 => A(24), C2 => n121, ZN => n44);
   U73 : INV_X1 port map( A => n43, ZN => n140);
   U74 : AOI222_X1 port map( A1 => B(25), A2 => n130, B1 => C(25), B2 => n123, 
                           C1 => A(25), C2 => n121, ZN => n43);
   U75 : INV_X1 port map( A => n42, ZN => n139);
   U76 : AOI222_X1 port map( A1 => B(26), A2 => n130, B1 => C(26), B2 => n123, 
                           C1 => A(26), C2 => n121, ZN => n42);
   U77 : INV_X1 port map( A => n41, ZN => n138);
   U78 : AOI222_X1 port map( A1 => B(27), A2 => n130, B1 => C(27), B2 => n123, 
                           C1 => A(27), C2 => n121, ZN => n41);
   U79 : INV_X1 port map( A => n40, ZN => n137);
   U80 : AOI222_X1 port map( A1 => B(28), A2 => n130, B1 => C(28), B2 => n123, 
                           C1 => A(28), C2 => n121, ZN => n40);
   U81 : INV_X1 port map( A => n39, ZN => n136);
   U82 : AOI222_X1 port map( A1 => B(29), A2 => n130, B1 => C(29), B2 => n123, 
                           C1 => A(29), C2 => n121, ZN => n39);
   U83 : INV_X1 port map( A => n38, ZN => n135);
   U84 : AOI222_X1 port map( A1 => B(30), A2 => n130, B1 => C(30), B2 => n123, 
                           C1 => A(30), C2 => n121, ZN => n38);
   U85 : INV_X1 port map( A => n34, ZN => n134);
   U86 : AOI222_X1 port map( A1 => B(31), A2 => n130, B1 => C(31), B2 => n123, 
                           C1 => A(31), C2 => n121, ZN => n34);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_3 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_3;

architecture SYN_Behavioral of MUX3to1_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n132, D => n134, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n132, D => n135, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n132, D => n136, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n132, D => n137, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n132, D => n138, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n132, D => n139, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n132, D => n140, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n131, D => n141, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n132, D => n142, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n132, D => n143, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n132, D => n144, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n133, D => n145, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n133, D => n146, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n133, D => n147, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n133, D => n148, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n133, D => n149, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n133, D => n150, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n133, D => n151, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n133, D => n152, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n133, D => n153, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n133, D => n154, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n132, D => n155, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n131, D => n156, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n131, D => n157, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n131, D => n158, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n131, D => n159, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n131, D => n160, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n131, D => n161, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n131, D => n162, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n131, D => n163, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n131, D => n164, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n131, D => n165, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n119, A2 => n128, A3 => n125, ZN => N12);
   U4 : BUF_X1 port map( A => n37, Z => n122);
   U5 : BUF_X1 port map( A => n36, Z => n126);
   U6 : BUF_X1 port map( A => n35, Z => n127);
   U7 : BUF_X1 port map( A => N12, Z => n131);
   U8 : BUF_X1 port map( A => N12, Z => n132);
   U9 : BUF_X1 port map( A => N12, Z => n133);
   U10 : BUF_X1 port map( A => n126, Z => n124);
   U11 : BUF_X1 port map( A => n126, Z => n123);
   U12 : BUF_X1 port map( A => n122, Z => n119);
   U13 : BUF_X1 port map( A => n122, Z => n120);
   U14 : BUF_X1 port map( A => n127, Z => n128);
   U15 : BUF_X1 port map( A => n127, Z => n129);
   U16 : BUF_X1 port map( A => n126, Z => n125);
   U17 : BUF_X1 port map( A => n122, Z => n121);
   U18 : BUF_X1 port map( A => n127, Z => n130);
   U19 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n37);
   U20 : NOR2_X1 port map( A1 => n166, A2 => SEL(0), ZN => n36);
   U21 : AND2_X1 port map( A1 => SEL(0), A2 => n166, ZN => n35);
   U22 : INV_X1 port map( A => SEL(1), ZN => n166);
   U23 : INV_X1 port map( A => n68, ZN => n165);
   U24 : AOI222_X1 port map( A1 => B(0), A2 => n128, B1 => C(0), B2 => n125, C1
                           => A(0), C2 => n119, ZN => n68);
   U25 : INV_X1 port map( A => n67, ZN => n164);
   U26 : AOI222_X1 port map( A1 => B(1), A2 => n128, B1 => C(1), B2 => n125, C1
                           => A(1), C2 => n119, ZN => n67);
   U27 : INV_X1 port map( A => n66, ZN => n163);
   U28 : AOI222_X1 port map( A1 => B(2), A2 => n128, B1 => C(2), B2 => n125, C1
                           => A(2), C2 => n119, ZN => n66);
   U29 : INV_X1 port map( A => n65, ZN => n162);
   U30 : AOI222_X1 port map( A1 => B(3), A2 => n128, B1 => C(3), B2 => n125, C1
                           => A(3), C2 => n119, ZN => n65);
   U31 : INV_X1 port map( A => n64, ZN => n161);
   U32 : AOI222_X1 port map( A1 => B(4), A2 => n128, B1 => C(4), B2 => n125, C1
                           => A(4), C2 => n119, ZN => n64);
   U33 : INV_X1 port map( A => n63, ZN => n160);
   U34 : AOI222_X1 port map( A1 => B(5), A2 => n128, B1 => C(5), B2 => n125, C1
                           => A(5), C2 => n119, ZN => n63);
   U35 : INV_X1 port map( A => n62, ZN => n159);
   U36 : AOI222_X1 port map( A1 => B(6), A2 => n128, B1 => C(6), B2 => n125, C1
                           => A(6), C2 => n119, ZN => n62);
   U37 : INV_X1 port map( A => n61, ZN => n158);
   U38 : AOI222_X1 port map( A1 => B(7), A2 => n128, B1 => C(7), B2 => n125, C1
                           => A(7), C2 => n119, ZN => n61);
   U39 : INV_X1 port map( A => n60, ZN => n157);
   U40 : AOI222_X1 port map( A1 => B(8), A2 => n128, B1 => C(8), B2 => n124, C1
                           => A(8), C2 => n119, ZN => n60);
   U41 : INV_X1 port map( A => n59, ZN => n156);
   U42 : AOI222_X1 port map( A1 => B(9), A2 => n128, B1 => C(9), B2 => n124, C1
                           => A(9), C2 => n119, ZN => n59);
   U43 : INV_X1 port map( A => n58, ZN => n155);
   U44 : AOI222_X1 port map( A1 => B(10), A2 => n128, B1 => C(10), B2 => n124, 
                           C1 => A(10), C2 => n119, ZN => n58);
   U45 : INV_X1 port map( A => n57, ZN => n154);
   U46 : AOI222_X1 port map( A1 => B(11), A2 => n129, B1 => C(11), B2 => n124, 
                           C1 => A(11), C2 => n120, ZN => n57);
   U47 : INV_X1 port map( A => n56, ZN => n153);
   U48 : AOI222_X1 port map( A1 => B(12), A2 => n129, B1 => C(12), B2 => n124, 
                           C1 => A(12), C2 => n120, ZN => n56);
   U49 : INV_X1 port map( A => n55, ZN => n152);
   U50 : AOI222_X1 port map( A1 => B(13), A2 => n129, B1 => C(13), B2 => n124, 
                           C1 => A(13), C2 => n120, ZN => n55);
   U51 : INV_X1 port map( A => n54, ZN => n151);
   U52 : AOI222_X1 port map( A1 => B(14), A2 => n129, B1 => C(14), B2 => n124, 
                           C1 => A(14), C2 => n120, ZN => n54);
   U53 : INV_X1 port map( A => n53, ZN => n150);
   U54 : AOI222_X1 port map( A1 => B(15), A2 => n129, B1 => C(15), B2 => n124, 
                           C1 => A(15), C2 => n120, ZN => n53);
   U55 : INV_X1 port map( A => n52, ZN => n149);
   U56 : AOI222_X1 port map( A1 => B(16), A2 => n129, B1 => C(16), B2 => n124, 
                           C1 => A(16), C2 => n120, ZN => n52);
   U57 : INV_X1 port map( A => n51, ZN => n148);
   U58 : AOI222_X1 port map( A1 => B(17), A2 => n129, B1 => C(17), B2 => n124, 
                           C1 => A(17), C2 => n120, ZN => n51);
   U59 : INV_X1 port map( A => n50, ZN => n147);
   U60 : AOI222_X1 port map( A1 => B(18), A2 => n129, B1 => C(18), B2 => n124, 
                           C1 => A(18), C2 => n120, ZN => n50);
   U61 : INV_X1 port map( A => n49, ZN => n146);
   U62 : AOI222_X1 port map( A1 => B(19), A2 => n129, B1 => C(19), B2 => n124, 
                           C1 => A(19), C2 => n120, ZN => n49);
   U63 : INV_X1 port map( A => n48, ZN => n145);
   U64 : AOI222_X1 port map( A1 => B(20), A2 => n129, B1 => C(20), B2 => n123, 
                           C1 => A(20), C2 => n120, ZN => n48);
   U65 : INV_X1 port map( A => n47, ZN => n144);
   U66 : AOI222_X1 port map( A1 => B(21), A2 => n129, B1 => C(21), B2 => n123, 
                           C1 => A(21), C2 => n120, ZN => n47);
   U67 : INV_X1 port map( A => n46, ZN => n143);
   U68 : AOI222_X1 port map( A1 => B(22), A2 => n129, B1 => C(22), B2 => n123, 
                           C1 => A(22), C2 => n120, ZN => n46);
   U69 : INV_X1 port map( A => n45, ZN => n142);
   U70 : AOI222_X1 port map( A1 => B(23), A2 => n130, B1 => C(23), B2 => n123, 
                           C1 => A(23), C2 => n121, ZN => n45);
   U71 : INV_X1 port map( A => n44, ZN => n141);
   U72 : AOI222_X1 port map( A1 => B(24), A2 => n130, B1 => C(24), B2 => n123, 
                           C1 => A(24), C2 => n121, ZN => n44);
   U73 : INV_X1 port map( A => n43, ZN => n140);
   U74 : AOI222_X1 port map( A1 => B(25), A2 => n130, B1 => C(25), B2 => n123, 
                           C1 => A(25), C2 => n121, ZN => n43);
   U75 : INV_X1 port map( A => n42, ZN => n139);
   U76 : AOI222_X1 port map( A1 => B(26), A2 => n130, B1 => C(26), B2 => n123, 
                           C1 => A(26), C2 => n121, ZN => n42);
   U77 : INV_X1 port map( A => n41, ZN => n138);
   U78 : AOI222_X1 port map( A1 => B(27), A2 => n130, B1 => C(27), B2 => n123, 
                           C1 => A(27), C2 => n121, ZN => n41);
   U79 : INV_X1 port map( A => n40, ZN => n137);
   U80 : AOI222_X1 port map( A1 => B(28), A2 => n130, B1 => C(28), B2 => n123, 
                           C1 => A(28), C2 => n121, ZN => n40);
   U81 : INV_X1 port map( A => n39, ZN => n136);
   U82 : AOI222_X1 port map( A1 => B(29), A2 => n130, B1 => C(29), B2 => n123, 
                           C1 => A(29), C2 => n121, ZN => n39);
   U83 : INV_X1 port map( A => n38, ZN => n135);
   U84 : AOI222_X1 port map( A1 => B(30), A2 => n130, B1 => C(30), B2 => n123, 
                           C1 => A(30), C2 => n121, ZN => n38);
   U85 : INV_X1 port map( A => n34, ZN => n134);
   U86 : AOI222_X1 port map( A1 => B(31), A2 => n130, B1 => C(31), B2 => n123, 
                           C1 => A(31), C2 => n121, ZN => n34);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_5;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n105, n106, n107, n140 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n140, Z => n106);
   U2 : BUF_X1 port map( A => n140, Z => n105);
   U3 : BUF_X1 port map( A => n140, Z => n107);
   U4 : INV_X1 port map( A => n61, ZN => Y(4));
   U5 : AOI22_X1 port map( A1 => A(4), A2 => n105, B1 => B(4), B2 => SEL, ZN =>
                           n61);
   U6 : INV_X1 port map( A => n64, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n105, B1 => B(1), B2 => SEL, ZN =>
                           n64);
   U8 : INV_X1 port map( A => n65, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n105, B1 => B(0), B2 => SEL, ZN =>
                           n65);
   U10 : INV_X1 port map( A => n63, ZN => Y(2));
   U11 : AOI22_X1 port map( A1 => A(2), A2 => n105, B1 => B(2), B2 => SEL, ZN 
                           => n63);
   U12 : INV_X1 port map( A => n62, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n105, B1 => B(3), B2 => SEL, ZN 
                           => n62);
   U14 : INV_X1 port map( A => n53, ZN => Y(12));
   U15 : AOI22_X1 port map( A1 => A(12), A2 => n106, B1 => B(12), B2 => SEL, ZN
                           => n53);
   U16 : INV_X1 port map( A => n57, ZN => Y(8));
   U17 : AOI22_X1 port map( A1 => A(8), A2 => n105, B1 => B(8), B2 => SEL, ZN 
                           => n57);
   U18 : INV_X1 port map( A => n59, ZN => Y(6));
   U19 : AOI22_X1 port map( A1 => A(6), A2 => n105, B1 => B(6), B2 => SEL, ZN 
                           => n59);
   U20 : INV_X1 port map( A => n55, ZN => Y(10));
   U21 : AOI22_X1 port map( A1 => A(10), A2 => n105, B1 => B(10), B2 => SEL, ZN
                           => n55);
   U22 : INV_X1 port map( A => n51, ZN => Y(14));
   U23 : AOI22_X1 port map( A1 => A(14), A2 => n106, B1 => B(14), B2 => SEL, ZN
                           => n51);
   U24 : INV_X1 port map( A => n50, ZN => Y(15));
   U25 : AOI22_X1 port map( A1 => A(15), A2 => n106, B1 => B(15), B2 => SEL, ZN
                           => n50);
   U26 : INV_X1 port map( A => n52, ZN => Y(13));
   U27 : AOI22_X1 port map( A1 => A(13), A2 => n106, B1 => B(13), B2 => SEL, ZN
                           => n52);
   U28 : INV_X1 port map( A => n54, ZN => Y(11));
   U29 : AOI22_X1 port map( A1 => A(11), A2 => n105, B1 => B(11), B2 => SEL, ZN
                           => n54);
   U30 : INV_X1 port map( A => n56, ZN => Y(9));
   U31 : AOI22_X1 port map( A1 => A(9), A2 => n105, B1 => B(9), B2 => SEL, ZN 
                           => n56);
   U32 : INV_X1 port map( A => n58, ZN => Y(7));
   U33 : AOI22_X1 port map( A1 => A(7), A2 => n105, B1 => B(7), B2 => SEL, ZN 
                           => n58);
   U34 : INV_X1 port map( A => n60, ZN => Y(5));
   U35 : AOI22_X1 port map( A1 => A(5), A2 => n105, B1 => B(5), B2 => SEL, ZN 
                           => n60);
   U36 : INV_X1 port map( A => n49, ZN => Y(16));
   U37 : AOI22_X1 port map( A1 => A(16), A2 => n106, B1 => B(16), B2 => SEL, ZN
                           => n49);
   U38 : INV_X1 port map( A => n45, ZN => Y(20));
   U39 : AOI22_X1 port map( A1 => A(20), A2 => n106, B1 => B(20), B2 => SEL, ZN
                           => n45);
   U40 : INV_X1 port map( A => n41, ZN => Y(24));
   U41 : AOI22_X1 port map( A1 => A(24), A2 => n107, B1 => B(24), B2 => SEL, ZN
                           => n41);
   U42 : INV_X1 port map( A => n48, ZN => Y(17));
   U43 : AOI22_X1 port map( A1 => A(17), A2 => n106, B1 => B(17), B2 => SEL, ZN
                           => n48);
   U44 : INV_X1 port map( A => n44, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n106, B1 => B(21), B2 => SEL, ZN
                           => n44);
   U46 : INV_X1 port map( A => n40, ZN => Y(25));
   U47 : AOI22_X1 port map( A1 => A(25), A2 => n107, B1 => B(25), B2 => SEL, ZN
                           => n40);
   U48 : INV_X1 port map( A => n37, ZN => Y(28));
   U49 : AOI22_X1 port map( A1 => A(28), A2 => n107, B1 => B(28), B2 => SEL, ZN
                           => n37);
   U50 : INV_X1 port map( A => n47, ZN => Y(18));
   U51 : AOI22_X1 port map( A1 => A(18), A2 => n106, B1 => B(18), B2 => SEL, ZN
                           => n47);
   U52 : INV_X1 port map( A => n46, ZN => Y(19));
   U53 : AOI22_X1 port map( A1 => A(19), A2 => n106, B1 => B(19), B2 => SEL, ZN
                           => n46);
   U54 : INV_X1 port map( A => n43, ZN => Y(22));
   U55 : AOI22_X1 port map( A1 => A(22), A2 => n106, B1 => B(22), B2 => SEL, ZN
                           => n43);
   U56 : INV_X1 port map( A => n42, ZN => Y(23));
   U57 : AOI22_X1 port map( A1 => A(23), A2 => n106, B1 => B(23), B2 => SEL, ZN
                           => n42);
   U58 : INV_X1 port map( A => n39, ZN => Y(26));
   U59 : AOI22_X1 port map( A1 => A(26), A2 => n107, B1 => B(26), B2 => SEL, ZN
                           => n39);
   U60 : INV_X1 port map( A => n38, ZN => Y(27));
   U61 : AOI22_X1 port map( A1 => A(27), A2 => n107, B1 => B(27), B2 => SEL, ZN
                           => n38);
   U62 : INV_X1 port map( A => n36, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n107, B1 => B(29), B2 => SEL, ZN
                           => n36);
   U64 : INV_X1 port map( A => n35, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n107, B1 => B(30), B2 => SEL, ZN
                           => n35);
   U66 : INV_X1 port map( A => n34, ZN => Y(31));
   U67 : AOI22_X1 port map( A1 => A(31), A2 => n107, B1 => SEL, B2 => B(31), ZN
                           => n34);
   U68 : INV_X1 port map( A => SEL, ZN => n140);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_6;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n105, n106, n107, n140 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n140, Z => n106);
   U2 : BUF_X1 port map( A => n140, Z => n105);
   U3 : BUF_X1 port map( A => n140, Z => n107);
   U4 : INV_X1 port map( A => n65, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n105, B1 => B(0), B2 => SEL, ZN =>
                           n65);
   U6 : INV_X1 port map( A => n64, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n105, B1 => B(1), B2 => SEL, ZN =>
                           n64);
   U8 : INV_X1 port map( A => n63, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n105, B1 => B(2), B2 => SEL, ZN =>
                           n63);
   U10 : INV_X1 port map( A => n62, ZN => Y(3));
   U11 : AOI22_X1 port map( A1 => A(3), A2 => n105, B1 => B(3), B2 => SEL, ZN 
                           => n62);
   U12 : INV_X1 port map( A => n61, ZN => Y(4));
   U13 : AOI22_X1 port map( A1 => A(4), A2 => n105, B1 => B(4), B2 => SEL, ZN 
                           => n61);
   U14 : INV_X1 port map( A => n60, ZN => Y(5));
   U15 : AOI22_X1 port map( A1 => A(5), A2 => n105, B1 => B(5), B2 => SEL, ZN 
                           => n60);
   U16 : INV_X1 port map( A => n59, ZN => Y(6));
   U17 : AOI22_X1 port map( A1 => A(6), A2 => n105, B1 => B(6), B2 => SEL, ZN 
                           => n59);
   U18 : INV_X1 port map( A => n58, ZN => Y(7));
   U19 : AOI22_X1 port map( A1 => A(7), A2 => n105, B1 => B(7), B2 => SEL, ZN 
                           => n58);
   U20 : INV_X1 port map( A => n57, ZN => Y(8));
   U21 : AOI22_X1 port map( A1 => A(8), A2 => n105, B1 => B(8), B2 => SEL, ZN 
                           => n57);
   U22 : INV_X1 port map( A => n56, ZN => Y(9));
   U23 : AOI22_X1 port map( A1 => A(9), A2 => n105, B1 => B(9), B2 => SEL, ZN 
                           => n56);
   U24 : INV_X1 port map( A => n55, ZN => Y(10));
   U25 : AOI22_X1 port map( A1 => A(10), A2 => n105, B1 => B(10), B2 => SEL, ZN
                           => n55);
   U26 : INV_X1 port map( A => n54, ZN => Y(11));
   U27 : AOI22_X1 port map( A1 => A(11), A2 => n105, B1 => B(11), B2 => SEL, ZN
                           => n54);
   U28 : INV_X1 port map( A => n53, ZN => Y(12));
   U29 : AOI22_X1 port map( A1 => A(12), A2 => n106, B1 => B(12), B2 => SEL, ZN
                           => n53);
   U30 : INV_X1 port map( A => n52, ZN => Y(13));
   U31 : AOI22_X1 port map( A1 => A(13), A2 => n106, B1 => B(13), B2 => SEL, ZN
                           => n52);
   U32 : INV_X1 port map( A => n51, ZN => Y(14));
   U33 : AOI22_X1 port map( A1 => A(14), A2 => n106, B1 => B(14), B2 => SEL, ZN
                           => n51);
   U34 : INV_X1 port map( A => n50, ZN => Y(15));
   U35 : AOI22_X1 port map( A1 => A(15), A2 => n106, B1 => B(15), B2 => SEL, ZN
                           => n50);
   U36 : INV_X1 port map( A => n49, ZN => Y(16));
   U37 : AOI22_X1 port map( A1 => A(16), A2 => n106, B1 => B(16), B2 => SEL, ZN
                           => n49);
   U38 : INV_X1 port map( A => n48, ZN => Y(17));
   U39 : AOI22_X1 port map( A1 => A(17), A2 => n106, B1 => B(17), B2 => SEL, ZN
                           => n48);
   U40 : INV_X1 port map( A => n47, ZN => Y(18));
   U41 : AOI22_X1 port map( A1 => A(18), A2 => n106, B1 => B(18), B2 => SEL, ZN
                           => n47);
   U42 : INV_X1 port map( A => n46, ZN => Y(19));
   U43 : AOI22_X1 port map( A1 => A(19), A2 => n106, B1 => B(19), B2 => SEL, ZN
                           => n46);
   U44 : INV_X1 port map( A => n45, ZN => Y(20));
   U45 : AOI22_X1 port map( A1 => A(20), A2 => n106, B1 => B(20), B2 => SEL, ZN
                           => n45);
   U46 : INV_X1 port map( A => n44, ZN => Y(21));
   U47 : AOI22_X1 port map( A1 => A(21), A2 => n106, B1 => B(21), B2 => SEL, ZN
                           => n44);
   U48 : INV_X1 port map( A => n43, ZN => Y(22));
   U49 : AOI22_X1 port map( A1 => A(22), A2 => n106, B1 => B(22), B2 => SEL, ZN
                           => n43);
   U50 : INV_X1 port map( A => n42, ZN => Y(23));
   U51 : AOI22_X1 port map( A1 => A(23), A2 => n106, B1 => B(23), B2 => SEL, ZN
                           => n42);
   U52 : INV_X1 port map( A => n41, ZN => Y(24));
   U53 : AOI22_X1 port map( A1 => A(24), A2 => n107, B1 => B(24), B2 => SEL, ZN
                           => n41);
   U54 : INV_X1 port map( A => n40, ZN => Y(25));
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n107, B1 => B(25), B2 => SEL, ZN
                           => n40);
   U56 : INV_X1 port map( A => n39, ZN => Y(26));
   U57 : AOI22_X1 port map( A1 => A(26), A2 => n107, B1 => B(26), B2 => SEL, ZN
                           => n39);
   U58 : INV_X1 port map( A => n38, ZN => Y(27));
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n107, B1 => B(27), B2 => SEL, ZN
                           => n38);
   U60 : INV_X1 port map( A => n37, ZN => Y(28));
   U61 : AOI22_X1 port map( A1 => A(28), A2 => n107, B1 => B(28), B2 => SEL, ZN
                           => n37);
   U62 : INV_X1 port map( A => n36, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n107, B1 => B(29), B2 => SEL, ZN
                           => n36);
   U64 : INV_X1 port map( A => n34, ZN => Y(31));
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n107, B1 => SEL, B2 => B(31), ZN
                           => n34);
   U66 : INV_X1 port map( A => n35, ZN => Y(30));
   U67 : AOI22_X1 port map( A1 => A(30), A2 => n107, B1 => B(30), B2 => SEL, ZN
                           => n35);
   U68 : INV_X1 port map( A => SEL, ZN => n140);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_7;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n96, n97, n98, n99, n100, n101, n102 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n101, ZN => n99);
   U2 : INV_X1 port map( A => n42, ZN => Y(23));
   U3 : INV_X1 port map( A => n43, ZN => Y(22));
   U4 : INV_X1 port map( A => n44, ZN => Y(21));
   U5 : INV_X1 port map( A => n45, ZN => Y(20));
   U6 : INV_X1 port map( A => n46, ZN => Y(19));
   U7 : INV_X1 port map( A => n47, ZN => Y(18));
   U8 : INV_X1 port map( A => n48, ZN => Y(17));
   U9 : INV_X1 port map( A => n49, ZN => Y(16));
   U10 : INV_X1 port map( A => n50, ZN => Y(15));
   U11 : INV_X1 port map( A => n51, ZN => Y(14));
   U12 : INV_X1 port map( A => n52, ZN => Y(13));
   U13 : INV_X1 port map( A => n53, ZN => Y(12));
   U14 : INV_X1 port map( A => n35, ZN => Y(30));
   U15 : INV_X1 port map( A => n36, ZN => Y(29));
   U16 : INV_X1 port map( A => n37, ZN => Y(28));
   U17 : INV_X1 port map( A => n38, ZN => Y(27));
   U18 : INV_X1 port map( A => n39, ZN => Y(26));
   U19 : INV_X1 port map( A => n40, ZN => Y(25));
   U20 : INV_X1 port map( A => n41, ZN => Y(24));
   U21 : INV_X1 port map( A => n34, ZN => Y(31));
   U22 : INV_X1 port map( A => n54, ZN => Y(11));
   U23 : INV_X1 port map( A => n55, ZN => Y(10));
   U24 : INV_X1 port map( A => n56, ZN => Y(9));
   U25 : INV_X1 port map( A => n57, ZN => Y(8));
   U26 : INV_X1 port map( A => n58, ZN => Y(7));
   U27 : INV_X1 port map( A => n59, ZN => Y(6));
   U28 : INV_X1 port map( A => n60, ZN => Y(5));
   U29 : INV_X1 port map( A => n61, ZN => Y(4));
   U30 : INV_X1 port map( A => n62, ZN => Y(3));
   U31 : BUF_X1 port map( A => SEL, Z => n101);
   U32 : INV_X1 port map( A => n64, ZN => Y(1));
   U33 : INV_X1 port map( A => n63, ZN => Y(2));
   U34 : BUF_X2 port map( A => n102, Z => n96);
   U35 : CLKBUF_X1 port map( A => n102, Z => n97);
   U36 : CLKBUF_X1 port map( A => n102, Z => n98);
   U37 : BUF_X1 port map( A => SEL, Z => n102);
   U38 : AOI22_X1 port map( A1 => A(12), A2 => n100, B1 => B(12), B2 => n97, ZN
                           => n53);
   U39 : AOI22_X1 port map( A1 => A(13), A2 => n100, B1 => B(13), B2 => n97, ZN
                           => n52);
   U40 : AOI22_X1 port map( A1 => A(14), A2 => n100, B1 => B(14), B2 => n97, ZN
                           => n51);
   U41 : AOI22_X1 port map( A1 => A(15), A2 => n100, B1 => B(15), B2 => n97, ZN
                           => n50);
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n100, B1 => B(16), B2 => n97, ZN
                           => n49);
   U43 : AOI22_X1 port map( A1 => A(17), A2 => n100, B1 => B(17), B2 => n97, ZN
                           => n48);
   U44 : AOI22_X1 port map( A1 => A(18), A2 => n100, B1 => B(18), B2 => n97, ZN
                           => n47);
   U45 : AOI22_X1 port map( A1 => A(19), A2 => n100, B1 => B(19), B2 => n97, ZN
                           => n46);
   U46 : AOI22_X1 port map( A1 => A(20), A2 => n100, B1 => B(20), B2 => n97, ZN
                           => n45);
   U47 : AOI22_X1 port map( A1 => A(21), A2 => n100, B1 => B(21), B2 => n97, ZN
                           => n44);
   U48 : AOI22_X1 port map( A1 => A(22), A2 => n100, B1 => B(22), B2 => n97, ZN
                           => n43);
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n100, B1 => B(23), B2 => n97, ZN
                           => n42);
   U50 : AOI22_X1 port map( A1 => A(24), A2 => n100, B1 => B(24), B2 => n98, ZN
                           => n41);
   U51 : AOI22_X1 port map( A1 => A(25), A2 => n100, B1 => B(25), B2 => n98, ZN
                           => n40);
   U52 : AOI22_X1 port map( A1 => A(26), A2 => n100, B1 => B(26), B2 => n98, ZN
                           => n39);
   U53 : AOI22_X1 port map( A1 => A(27), A2 => n100, B1 => B(27), B2 => n98, ZN
                           => n38);
   U54 : AOI22_X1 port map( A1 => A(28), A2 => n100, B1 => B(28), B2 => n98, ZN
                           => n37);
   U55 : AOI22_X1 port map( A1 => A(29), A2 => n100, B1 => B(29), B2 => n98, ZN
                           => n36);
   U56 : AOI22_X1 port map( A1 => A(30), A2 => n100, B1 => B(30), B2 => n98, ZN
                           => n35);
   U57 : AOI22_X1 port map( A1 => A(31), A2 => n100, B1 => n98, B2 => B(31), ZN
                           => n34);
   U58 : INV_X1 port map( A => n101, ZN => n100);
   U59 : INV_X1 port map( A => n65, ZN => Y(0));
   U60 : AOI22_X1 port map( A1 => A(3), A2 => n99, B1 => B(3), B2 => n96, ZN =>
                           n62);
   U61 : AOI22_X1 port map( A1 => A(4), A2 => n99, B1 => B(4), B2 => n96, ZN =>
                           n61);
   U62 : AOI22_X1 port map( A1 => A(5), A2 => n99, B1 => B(5), B2 => n96, ZN =>
                           n60);
   U63 : AOI22_X1 port map( A1 => A(6), A2 => n99, B1 => B(6), B2 => n96, ZN =>
                           n59);
   U64 : AOI22_X1 port map( A1 => A(7), A2 => n99, B1 => B(7), B2 => n96, ZN =>
                           n58);
   U65 : AOI22_X1 port map( A1 => A(8), A2 => n99, B1 => B(8), B2 => n96, ZN =>
                           n57);
   U66 : AOI22_X1 port map( A1 => A(9), A2 => n99, B1 => B(9), B2 => n96, ZN =>
                           n56);
   U67 : AOI22_X1 port map( A1 => A(10), A2 => n99, B1 => B(10), B2 => n96, ZN 
                           => n55);
   U68 : AOI22_X1 port map( A1 => A(11), A2 => n99, B1 => B(11), B2 => n96, ZN 
                           => n54);
   U69 : AOI22_X1 port map( A1 => A(2), A2 => n99, B1 => B(2), B2 => n96, ZN =>
                           n63);
   U70 : AOI22_X1 port map( A1 => A(1), A2 => n99, B1 => B(1), B2 => n96, ZN =>
                           n64);
   U71 : AOI22_X1 port map( A1 => A(0), A2 => n99, B1 => B(0), B2 => n96, ZN =>
                           n65);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_8 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_8;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n101, n102, n103, n136 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n136, Z => n101);
   U2 : BUF_X1 port map( A => n136, Z => n102);
   U3 : BUF_X1 port map( A => n136, Z => n103);
   U4 : INV_X1 port map( A => n64, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n101, B1 => B(1), B2 => SEL, ZN =>
                           n64);
   U6 : INV_X1 port map( A => n63, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n101, B1 => B(2), B2 => SEL, ZN =>
                           n63);
   U8 : INV_X1 port map( A => n62, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n101, B1 => B(3), B2 => SEL, ZN =>
                           n62);
   U10 : INV_X1 port map( A => n61, ZN => Y(4));
   U11 : AOI22_X1 port map( A1 => A(4), A2 => n101, B1 => B(4), B2 => SEL, ZN 
                           => n61);
   U12 : INV_X1 port map( A => n60, ZN => Y(5));
   U13 : AOI22_X1 port map( A1 => A(5), A2 => n101, B1 => B(5), B2 => SEL, ZN 
                           => n60);
   U14 : INV_X1 port map( A => n59, ZN => Y(6));
   U15 : AOI22_X1 port map( A1 => A(6), A2 => n101, B1 => B(6), B2 => SEL, ZN 
                           => n59);
   U16 : INV_X1 port map( A => n58, ZN => Y(7));
   U17 : AOI22_X1 port map( A1 => A(7), A2 => n101, B1 => B(7), B2 => SEL, ZN 
                           => n58);
   U18 : INV_X1 port map( A => n57, ZN => Y(8));
   U19 : AOI22_X1 port map( A1 => A(8), A2 => n101, B1 => B(8), B2 => SEL, ZN 
                           => n57);
   U20 : INV_X1 port map( A => n56, ZN => Y(9));
   U21 : AOI22_X1 port map( A1 => A(9), A2 => n101, B1 => B(9), B2 => SEL, ZN 
                           => n56);
   U22 : INV_X1 port map( A => n55, ZN => Y(10));
   U23 : AOI22_X1 port map( A1 => A(10), A2 => n101, B1 => B(10), B2 => SEL, ZN
                           => n55);
   U24 : INV_X1 port map( A => n54, ZN => Y(11));
   U25 : AOI22_X1 port map( A1 => A(11), A2 => n101, B1 => B(11), B2 => SEL, ZN
                           => n54);
   U26 : INV_X1 port map( A => n53, ZN => Y(12));
   U27 : AOI22_X1 port map( A1 => A(12), A2 => n102, B1 => B(12), B2 => SEL, ZN
                           => n53);
   U28 : INV_X1 port map( A => n52, ZN => Y(13));
   U29 : AOI22_X1 port map( A1 => A(13), A2 => n102, B1 => B(13), B2 => SEL, ZN
                           => n52);
   U30 : INV_X1 port map( A => n51, ZN => Y(14));
   U31 : AOI22_X1 port map( A1 => A(14), A2 => n102, B1 => B(14), B2 => SEL, ZN
                           => n51);
   U32 : INV_X1 port map( A => n50, ZN => Y(15));
   U33 : AOI22_X1 port map( A1 => A(15), A2 => n102, B1 => B(15), B2 => SEL, ZN
                           => n50);
   U34 : INV_X1 port map( A => n49, ZN => Y(16));
   U35 : AOI22_X1 port map( A1 => A(16), A2 => n102, B1 => B(16), B2 => SEL, ZN
                           => n49);
   U36 : INV_X1 port map( A => n48, ZN => Y(17));
   U37 : INV_X1 port map( A => n47, ZN => Y(18));
   U38 : INV_X1 port map( A => n46, ZN => Y(19));
   U39 : INV_X1 port map( A => n45, ZN => Y(20));
   U40 : INV_X1 port map( A => n44, ZN => Y(21));
   U41 : INV_X1 port map( A => n43, ZN => Y(22));
   U42 : INV_X1 port map( A => n42, ZN => Y(23));
   U43 : AOI22_X1 port map( A1 => A(23), A2 => n102, B1 => B(23), B2 => SEL, ZN
                           => n42);
   U44 : INV_X1 port map( A => n41, ZN => Y(24));
   U45 : AOI22_X1 port map( A1 => A(24), A2 => n103, B1 => B(24), B2 => SEL, ZN
                           => n41);
   U46 : INV_X1 port map( A => n40, ZN => Y(25));
   U47 : INV_X1 port map( A => n39, ZN => Y(26));
   U48 : INV_X1 port map( A => n38, ZN => Y(27));
   U49 : INV_X1 port map( A => n37, ZN => Y(28));
   U50 : INV_X1 port map( A => n36, ZN => Y(29));
   U51 : INV_X1 port map( A => n35, ZN => Y(30));
   U52 : INV_X1 port map( A => n65, ZN => Y(0));
   U53 : AOI22_X1 port map( A1 => A(0), A2 => n101, B1 => B(0), B2 => SEL, ZN 
                           => n65);
   U54 : INV_X1 port map( A => SEL, ZN => n136);
   U55 : INV_X1 port map( A => n34, ZN => Y(31));
   U56 : AOI22_X1 port map( A1 => A(19), A2 => n102, B1 => B(19), B2 => SEL, ZN
                           => n46);
   U57 : AOI22_X1 port map( A1 => A(17), A2 => n102, B1 => B(17), B2 => SEL, ZN
                           => n48);
   U58 : AOI22_X1 port map( A1 => A(22), A2 => n102, B1 => B(22), B2 => SEL, ZN
                           => n43);
   U59 : AOI22_X1 port map( A1 => A(30), A2 => n103, B1 => B(30), B2 => SEL, ZN
                           => n35);
   U60 : AOI22_X1 port map( A1 => A(29), A2 => n103, B1 => B(29), B2 => SEL, ZN
                           => n36);
   U61 : AOI22_X1 port map( A1 => A(28), A2 => n103, B1 => B(28), B2 => SEL, ZN
                           => n37);
   U62 : AOI22_X1 port map( A1 => A(27), A2 => n103, B1 => B(27), B2 => SEL, ZN
                           => n38);
   U63 : AOI22_X1 port map( A1 => A(26), A2 => n103, B1 => B(26), B2 => SEL, ZN
                           => n39);
   U64 : AOI22_X1 port map( A1 => A(25), A2 => n103, B1 => B(25), B2 => SEL, ZN
                           => n40);
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n103, B1 => SEL, B2 => B(31), ZN
                           => n34);
   U66 : AOI22_X1 port map( A1 => A(20), A2 => n102, B1 => B(20), B2 => SEL, ZN
                           => n45);
   U67 : AOI22_X1 port map( A1 => A(21), A2 => n102, B1 => B(21), B2 => SEL, ZN
                           => n44);
   U68 : AOI22_X1 port map( A1 => A(18), A2 => n102, B1 => B(18), B2 => SEL, ZN
                           => n47);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_0;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n69, Z => n72);
   U2 : BUF_X1 port map( A => n69, Z => n73);
   U3 : BUF_X1 port map( A => n73, Z => n68);
   U4 : BUF_X1 port map( A => n73, Z => n66);
   U5 : BUF_X1 port map( A => n73, Z => n67);
   U6 : INV_X1 port map( A => n72, ZN => n70);
   U7 : INV_X1 port map( A => n54, ZN => Y(1));
   U8 : BUF_X1 port map( A => SEL, Z => n69);
   U9 : INV_X1 port map( A => n65, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n70, B1 => B(0), B2 => n66, ZN =>
                           n65);
   U11 : INV_X1 port map( A => n36, ZN => Y(7));
   U12 : AOI22_X1 port map( A1 => A(7), A2 => n71, B1 => B(7), B2 => n68, ZN =>
                           n36);
   U13 : INV_X1 port map( A => n38, ZN => Y(5));
   U14 : AOI22_X1 port map( A1 => A(5), A2 => n71, B1 => B(5), B2 => n68, ZN =>
                           n38);
   U15 : INV_X1 port map( A => n37, ZN => Y(6));
   U16 : INV_X1 port map( A => n40, ZN => Y(3));
   U17 : AOI22_X1 port map( A1 => A(3), A2 => n71, B1 => B(3), B2 => n67, ZN =>
                           n40);
   U18 : INV_X1 port map( A => n39, ZN => Y(4));
   U19 : AOI22_X1 port map( A1 => A(4), A2 => n71, B1 => B(4), B2 => n68, ZN =>
                           n39);
   U20 : INV_X1 port map( A => n64, ZN => Y(10));
   U21 : AOI22_X1 port map( A1 => A(10), A2 => n70, B1 => B(10), B2 => n66, ZN 
                           => n64);
   U22 : INV_X1 port map( A => n35, ZN => Y(8));
   U23 : AOI22_X1 port map( A1 => A(8), A2 => n71, B1 => B(8), B2 => n68, ZN =>
                           n35);
   U24 : INV_X1 port map( A => n34, ZN => Y(9));
   U25 : AOI22_X1 port map( A1 => A(9), A2 => n71, B1 => n68, B2 => B(9), ZN =>
                           n34);
   U26 : INV_X1 port map( A => n63, ZN => Y(11));
   U27 : AOI22_X1 port map( A1 => A(11), A2 => n70, B1 => B(11), B2 => n66, ZN 
                           => n63);
   U28 : INV_X1 port map( A => n60, ZN => Y(14));
   U29 : AOI22_X1 port map( A1 => A(14), A2 => n70, B1 => B(14), B2 => n66, ZN 
                           => n60);
   U30 : INV_X1 port map( A => n59, ZN => Y(15));
   U31 : AOI22_X1 port map( A1 => A(15), A2 => n70, B1 => B(15), B2 => n66, ZN 
                           => n59);
   U32 : INV_X1 port map( A => n61, ZN => Y(13));
   U33 : AOI22_X1 port map( A1 => A(13), A2 => n70, B1 => B(13), B2 => n66, ZN 
                           => n61);
   U34 : INV_X1 port map( A => n62, ZN => Y(12));
   U35 : AOI22_X1 port map( A1 => A(12), A2 => n70, B1 => B(12), B2 => n66, ZN 
                           => n62);
   U36 : INV_X1 port map( A => n57, ZN => Y(17));
   U37 : AOI22_X1 port map( A1 => A(17), A2 => n70, B1 => B(17), B2 => n66, ZN 
                           => n57);
   U38 : INV_X1 port map( A => n56, ZN => Y(18));
   U39 : AOI22_X1 port map( A1 => A(18), A2 => n70, B1 => B(18), B2 => n66, ZN 
                           => n56);
   U40 : INV_X1 port map( A => n55, ZN => Y(19));
   U41 : AOI22_X1 port map( A1 => A(19), A2 => n70, B1 => B(19), B2 => n66, ZN 
                           => n55);
   U42 : INV_X1 port map( A => n58, ZN => Y(16));
   U43 : AOI22_X1 port map( A1 => A(16), A2 => n70, B1 => B(16), B2 => n66, ZN 
                           => n58);
   U44 : INV_X1 port map( A => n52, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n71, B1 => B(21), B2 => n67, ZN 
                           => n52);
   U46 : INV_X1 port map( A => n51, ZN => Y(22));
   U47 : AOI22_X1 port map( A1 => A(22), A2 => n71, B1 => B(22), B2 => n67, ZN 
                           => n51);
   U48 : INV_X1 port map( A => n50, ZN => Y(23));
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n71, B1 => B(23), B2 => n67, ZN 
                           => n50);
   U50 : INV_X1 port map( A => n53, ZN => Y(20));
   U51 : AOI22_X1 port map( A1 => A(20), A2 => n71, B1 => B(20), B2 => n66, ZN 
                           => n53);
   U52 : INV_X1 port map( A => n48, ZN => Y(25));
   U53 : AOI22_X1 port map( A1 => A(25), A2 => n71, B1 => B(25), B2 => n67, ZN 
                           => n48);
   U54 : INV_X1 port map( A => n47, ZN => Y(26));
   U55 : AOI22_X1 port map( A1 => A(26), A2 => n71, B1 => B(26), B2 => n67, ZN 
                           => n47);
   U56 : INV_X1 port map( A => n49, ZN => Y(24));
   U57 : AOI22_X1 port map( A1 => A(24), A2 => n71, B1 => B(24), B2 => n67, ZN 
                           => n49);
   U58 : INV_X1 port map( A => n46, ZN => Y(27));
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n71, B1 => B(27), B2 => n67, ZN 
                           => n46);
   U60 : INV_X1 port map( A => n45, ZN => Y(28));
   U61 : AOI22_X1 port map( A1 => A(28), A2 => n71, B1 => B(28), B2 => n67, ZN 
                           => n45);
   U62 : INV_X1 port map( A => n44, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n71, B1 => B(29), B2 => n67, ZN 
                           => n44);
   U64 : INV_X1 port map( A => n42, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n71, B1 => B(30), B2 => n67, ZN 
                           => n42);
   U66 : INV_X1 port map( A => n41, ZN => Y(31));
   U67 : AOI22_X1 port map( A1 => A(31), A2 => n71, B1 => B(31), B2 => n67, ZN 
                           => n41);
   U68 : INV_X1 port map( A => n72, ZN => n71);
   U69 : AOI22_X1 port map( A1 => A(2), A2 => n71, B1 => B(2), B2 => n68, ZN =>
                           n43);
   U70 : AOI22_X1 port map( A1 => A(6), A2 => n71, B1 => B(6), B2 => n68, ZN =>
                           n37);
   U71 : INV_X1 port map( A => n43, ZN => Y(2));
   U72 : AOI22_X1 port map( A1 => A(1), A2 => n70, B1 => B(1), B2 => n68, ZN =>
                           n54);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_0 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_0;

architecture SYN_Behavioral of MUX3to1_NBIT32_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n84, D => n117, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n84, D => n116, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n84, D => n115, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n84, D => n114, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n84, D => n113, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n84, D => n112, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n84, D => n111, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n84, D => n110, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n84, D => n109, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n84, D => n108, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n83, D => n107, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n85, D => n106, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n85, D => n105, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n85, D => n104, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n85, D => n103, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n85, D => n102, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n85, D => n101, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n85, D => n100, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n85, D => n99, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n85, D => n98, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n85, D => n97, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n84, D => n96, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n83, D => n95, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n83, D => n94, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n83, D => n93, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n83, D => n92, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n83, D => n91, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n83, D => n90, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n83, D => n89, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n83, D => n88, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n83, D => n87, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n83, D => n86, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n71, A2 => n80, A3 => n77, ZN => N12);
   U4 : BUF_X1 port map( A => n37, Z => n74);
   U5 : BUF_X1 port map( A => n36, Z => n78);
   U6 : BUF_X1 port map( A => n35, Z => n79);
   U7 : BUF_X1 port map( A => N12, Z => n83);
   U8 : BUF_X1 port map( A => N12, Z => n84);
   U9 : BUF_X1 port map( A => N12, Z => n85);
   U10 : BUF_X1 port map( A => n78, Z => n76);
   U11 : BUF_X1 port map( A => n78, Z => n75);
   U12 : BUF_X1 port map( A => n74, Z => n71);
   U13 : BUF_X1 port map( A => n74, Z => n72);
   U14 : BUF_X1 port map( A => n79, Z => n80);
   U15 : BUF_X1 port map( A => n79, Z => n81);
   U16 : BUF_X1 port map( A => n78, Z => n77);
   U17 : BUF_X1 port map( A => n74, Z => n73);
   U18 : BUF_X1 port map( A => n79, Z => n82);
   U19 : INV_X1 port map( A => SEL(1), ZN => n118);
   U20 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n37);
   U21 : NOR2_X1 port map( A1 => n118, A2 => SEL(0), ZN => n36);
   U22 : AND2_X1 port map( A1 => SEL(0), A2 => n118, ZN => n35);
   U23 : INV_X1 port map( A => n68, ZN => n86);
   U24 : AOI222_X1 port map( A1 => B(0), A2 => n80, B1 => C(0), B2 => n77, C1 
                           => A(0), C2 => n71, ZN => n68);
   U25 : INV_X1 port map( A => n67, ZN => n87);
   U26 : AOI222_X1 port map( A1 => B(1), A2 => n80, B1 => C(1), B2 => n77, C1 
                           => A(1), C2 => n71, ZN => n67);
   U27 : INV_X1 port map( A => n66, ZN => n88);
   U28 : AOI222_X1 port map( A1 => B(2), A2 => n80, B1 => C(2), B2 => n77, C1 
                           => A(2), C2 => n71, ZN => n66);
   U29 : INV_X1 port map( A => n65, ZN => n89);
   U30 : AOI222_X1 port map( A1 => B(3), A2 => n80, B1 => C(3), B2 => n77, C1 
                           => A(3), C2 => n71, ZN => n65);
   U31 : INV_X1 port map( A => n64, ZN => n90);
   U32 : AOI222_X1 port map( A1 => B(4), A2 => n80, B1 => C(4), B2 => n77, C1 
                           => A(4), C2 => n71, ZN => n64);
   U33 : INV_X1 port map( A => n63, ZN => n91);
   U34 : AOI222_X1 port map( A1 => B(5), A2 => n80, B1 => C(5), B2 => n77, C1 
                           => A(5), C2 => n71, ZN => n63);
   U35 : INV_X1 port map( A => n62, ZN => n92);
   U36 : AOI222_X1 port map( A1 => B(6), A2 => n80, B1 => C(6), B2 => n77, C1 
                           => A(6), C2 => n71, ZN => n62);
   U37 : INV_X1 port map( A => n61, ZN => n93);
   U38 : AOI222_X1 port map( A1 => B(7), A2 => n80, B1 => C(7), B2 => n77, C1 
                           => A(7), C2 => n71, ZN => n61);
   U39 : INV_X1 port map( A => n60, ZN => n94);
   U40 : AOI222_X1 port map( A1 => B(8), A2 => n80, B1 => C(8), B2 => n76, C1 
                           => A(8), C2 => n71, ZN => n60);
   U41 : INV_X1 port map( A => n59, ZN => n95);
   U42 : AOI222_X1 port map( A1 => B(9), A2 => n80, B1 => C(9), B2 => n76, C1 
                           => A(9), C2 => n71, ZN => n59);
   U43 : INV_X1 port map( A => n58, ZN => n96);
   U44 : AOI222_X1 port map( A1 => B(10), A2 => n80, B1 => C(10), B2 => n76, C1
                           => A(10), C2 => n71, ZN => n58);
   U45 : INV_X1 port map( A => n57, ZN => n97);
   U46 : AOI222_X1 port map( A1 => B(11), A2 => n81, B1 => C(11), B2 => n76, C1
                           => A(11), C2 => n72, ZN => n57);
   U47 : INV_X1 port map( A => n56, ZN => n98);
   U48 : AOI222_X1 port map( A1 => B(12), A2 => n81, B1 => C(12), B2 => n76, C1
                           => A(12), C2 => n72, ZN => n56);
   U49 : INV_X1 port map( A => n55, ZN => n99);
   U50 : AOI222_X1 port map( A1 => B(13), A2 => n81, B1 => C(13), B2 => n76, C1
                           => A(13), C2 => n72, ZN => n55);
   U51 : INV_X1 port map( A => n54, ZN => n100);
   U52 : AOI222_X1 port map( A1 => B(14), A2 => n81, B1 => C(14), B2 => n76, C1
                           => A(14), C2 => n72, ZN => n54);
   U53 : INV_X1 port map( A => n53, ZN => n101);
   U54 : AOI222_X1 port map( A1 => B(15), A2 => n81, B1 => C(15), B2 => n76, C1
                           => A(15), C2 => n72, ZN => n53);
   U55 : INV_X1 port map( A => n52, ZN => n102);
   U56 : AOI222_X1 port map( A1 => B(16), A2 => n81, B1 => C(16), B2 => n76, C1
                           => A(16), C2 => n72, ZN => n52);
   U57 : INV_X1 port map( A => n51, ZN => n103);
   U58 : AOI222_X1 port map( A1 => B(17), A2 => n81, B1 => C(17), B2 => n76, C1
                           => A(17), C2 => n72, ZN => n51);
   U59 : INV_X1 port map( A => n50, ZN => n104);
   U60 : AOI222_X1 port map( A1 => B(18), A2 => n81, B1 => C(18), B2 => n76, C1
                           => A(18), C2 => n72, ZN => n50);
   U61 : INV_X1 port map( A => n49, ZN => n105);
   U62 : AOI222_X1 port map( A1 => B(19), A2 => n81, B1 => C(19), B2 => n76, C1
                           => A(19), C2 => n72, ZN => n49);
   U63 : INV_X1 port map( A => n48, ZN => n106);
   U64 : AOI222_X1 port map( A1 => B(20), A2 => n81, B1 => C(20), B2 => n75, C1
                           => A(20), C2 => n72, ZN => n48);
   U65 : INV_X1 port map( A => n47, ZN => n107);
   U66 : AOI222_X1 port map( A1 => B(21), A2 => n81, B1 => C(21), B2 => n75, C1
                           => A(21), C2 => n72, ZN => n47);
   U67 : INV_X1 port map( A => n46, ZN => n108);
   U68 : AOI222_X1 port map( A1 => B(22), A2 => n81, B1 => C(22), B2 => n75, C1
                           => A(22), C2 => n72, ZN => n46);
   U69 : INV_X1 port map( A => n45, ZN => n109);
   U70 : AOI222_X1 port map( A1 => B(23), A2 => n82, B1 => C(23), B2 => n75, C1
                           => A(23), C2 => n73, ZN => n45);
   U71 : INV_X1 port map( A => n44, ZN => n110);
   U72 : AOI222_X1 port map( A1 => B(24), A2 => n82, B1 => C(24), B2 => n75, C1
                           => A(24), C2 => n73, ZN => n44);
   U73 : INV_X1 port map( A => n43, ZN => n111);
   U74 : AOI222_X1 port map( A1 => B(25), A2 => n82, B1 => C(25), B2 => n75, C1
                           => A(25), C2 => n73, ZN => n43);
   U75 : INV_X1 port map( A => n42, ZN => n112);
   U76 : AOI222_X1 port map( A1 => B(26), A2 => n82, B1 => C(26), B2 => n75, C1
                           => A(26), C2 => n73, ZN => n42);
   U77 : INV_X1 port map( A => n41, ZN => n113);
   U78 : AOI222_X1 port map( A1 => B(27), A2 => n82, B1 => C(27), B2 => n75, C1
                           => A(27), C2 => n73, ZN => n41);
   U79 : INV_X1 port map( A => n40, ZN => n114);
   U80 : AOI222_X1 port map( A1 => B(28), A2 => n82, B1 => C(28), B2 => n75, C1
                           => A(28), C2 => n73, ZN => n40);
   U81 : INV_X1 port map( A => n39, ZN => n115);
   U82 : AOI222_X1 port map( A1 => B(29), A2 => n82, B1 => C(29), B2 => n75, C1
                           => A(29), C2 => n73, ZN => n39);
   U83 : INV_X1 port map( A => n38, ZN => n116);
   U84 : AOI222_X1 port map( A1 => B(30), A2 => n82, B1 => C(30), B2 => n75, C1
                           => A(30), C2 => n73, ZN => n38);
   U85 : INV_X1 port map( A => n34, ZN => n117);
   U86 : AOI222_X1 port map( A1 => B(31), A2 => n82, B1 => C(31), B2 => n75, C1
                           => A(31), C2 => n73, ZN => n34);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Sum : out std_logic_vector 
         (31 downto 0));

end PC_adder_1;

architecture SYN_Behavioral of PC_adder_1 is

   component PC_adder_1_DW01_add_0_DW01_add_128
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1583 : std_logic;

begin
   
   n1 <= '0';
   add_16 : PC_adder_1_DW01_add_0_DW01_add_128 port map( A(31) => A(31), A(30) 
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => n1, SUM(31) => Sum(31),
                           SUM(30) => Sum(30), SUM(29) => Sum(29), SUM(28) => 
                           Sum(28), SUM(27) => Sum(27), SUM(26) => Sum(26), 
                           SUM(25) => Sum(25), SUM(24) => Sum(24), SUM(23) => 
                           Sum(23), SUM(22) => Sum(22), SUM(21) => Sum(21), 
                           SUM(20) => Sum(20), SUM(19) => Sum(19), SUM(18) => 
                           Sum(18), SUM(17) => Sum(17), SUM(16) => Sum(16), 
                           SUM(15) => Sum(15), SUM(14) => Sum(14), SUM(13) => 
                           Sum(13), SUM(12) => Sum(12), SUM(11) => Sum(11), 
                           SUM(10) => Sum(10), SUM(9) => Sum(9), SUM(8) => 
                           Sum(8), SUM(7) => Sum(7), SUM(6) => Sum(6), SUM(5) 
                           => Sum(5), SUM(4) => Sum(4), SUM(3) => Sum(3), 
                           SUM(2) => Sum(2), SUM(1) => Sum(1), SUM(0) => Sum(0)
                           , CO => n_1583);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Sum : out std_logic_vector 
         (31 downto 0));

end PC_adder_0;

architecture SYN_Behavioral of PC_adder_0 is

   component PC_adder_0_DW01_add_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1584 : std_logic;

begin
   
   n2 <= '0';
   add_16 : PC_adder_0_DW01_add_2 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(31) => Sum(31), 
                           SUM(30) => Sum(30), SUM(29) => Sum(29), SUM(28) => 
                           Sum(28), SUM(27) => Sum(27), SUM(26) => Sum(26), 
                           SUM(25) => Sum(25), SUM(24) => Sum(24), SUM(23) => 
                           Sum(23), SUM(22) => Sum(22), SUM(21) => Sum(21), 
                           SUM(20) => Sum(20), SUM(19) => Sum(19), SUM(18) => 
                           Sum(18), SUM(17) => Sum(17), SUM(16) => Sum(16), 
                           SUM(15) => Sum(15), SUM(14) => Sum(14), SUM(13) => 
                           Sum(13), SUM(12) => Sum(12), SUM(11) => Sum(11), 
                           SUM(10) => Sum(10), SUM(9) => Sum(9), SUM(8) => 
                           Sum(8), SUM(7) => Sum(7), SUM(6) => Sum(6), SUM(5) 
                           => Sum(5), SUM(4) => Sum(4), SUM(3) => Sum(3), 
                           SUM(2) => Sum(2), SUM(1) => Sum(1), SUM(0) => Sum(0)
                           , CO => n_1584);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_4 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_4;

architecture SYN_Behavioral of REG_NBIT32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n215, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n215, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n215, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n215, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n215, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n215, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n215, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n215, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n215, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n216, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n215, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n216, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n215, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n216, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n216, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n215, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n217, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n217, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n217, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n217, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n216, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n216, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n216, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n216, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n206, Z => n214);
   U3 : BUF_X1 port map( A => n206, Z => n213);
   U4 : BUF_X1 port map( A => n214, Z => n208);
   U5 : BUF_X1 port map( A => n214, Z => n207);
   U6 : BUF_X1 port map( A => n214, Z => n209);
   U7 : BUF_X1 port map( A => n213, Z => n211);
   U8 : BUF_X1 port map( A => n213, Z => n210);
   U9 : BUF_X1 port map( A => n218, Z => n216);
   U10 : BUF_X1 port map( A => n218, Z => n215);
   U11 : BUF_X1 port map( A => n218, Z => n217);
   U12 : BUF_X1 port map( A => n213, Z => n212);
   U13 : INV_X1 port map( A => reset, ZN => n218);
   U14 : BUF_X1 port map( A => enable, Z => n206);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n2, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n212, A2 => data_in(0), ZN => n2);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n209, A => n3, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n207, ZN => n3);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n209, A => n4, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n207, ZN => n4);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n5, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n207, ZN => n5);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n209, A => n6, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n207, ZN => n6);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n209, A => n7, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n208, ZN => n7);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n8, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n208, ZN => n8);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n209, A => n9, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n208, ZN => n9);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n210, A => n10, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n208, ZN => n10);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n210, A => n11, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n209, ZN => n11);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n12, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n208, ZN => n12);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n210, A => n13, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n209, ZN => n13);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n210, A => n14, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n209, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n210, A => n15, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n209, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n210, A => n16, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n209, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n210, A => n17, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n209, ZN => n17);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n211, A => n18, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n209, ZN => n18);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n211, A => n19, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n208, ZN => n19);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n211, A => n20, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n208, ZN => n20);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n211, A => n21, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n208, ZN => n21);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n211, A => n22, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n208, ZN => n22);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n211, A => n23, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n208, ZN => n23);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n24, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n208, ZN => n24);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n211, A => n25, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n208, ZN => n25);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n211, A => n26, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n207, ZN => n26);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n211, A => n27, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n207, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n211, A => n28, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n207, ZN => n28);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n211, A => n29, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n207, ZN => n29);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n212, A => n30, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n207, ZN => n30);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n212, A => n31, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n207, ZN => n31);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n212, A => n32, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n207, ZN => n32);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n210, A => n33, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n207, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_5 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_5;

architecture SYN_Behavioral of REG_NBIT32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n215, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n215, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n215, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n215, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n215, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n215, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n215, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n215, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n216, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n216, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n215, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n215, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n215, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n216, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n215, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n217, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n216, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n216, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n216, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n216, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n206, Z => n214);
   U3 : BUF_X1 port map( A => n206, Z => n213);
   U4 : BUF_X1 port map( A => n214, Z => n208);
   U5 : BUF_X1 port map( A => n214, Z => n207);
   U6 : BUF_X1 port map( A => n214, Z => n209);
   U7 : BUF_X1 port map( A => n213, Z => n211);
   U8 : BUF_X1 port map( A => n213, Z => n210);
   U9 : BUF_X1 port map( A => n218, Z => n216);
   U10 : BUF_X1 port map( A => n218, Z => n215);
   U11 : BUF_X1 port map( A => n218, Z => n217);
   U12 : BUF_X1 port map( A => n213, Z => n212);
   U13 : INV_X1 port map( A => reset, ZN => n218);
   U14 : BUF_X1 port map( A => enable, Z => n206);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n2, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n212, A2 => data_in(0), ZN => n2);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n209, A => n3, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n207, ZN => n3);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n209, A => n4, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n207, ZN => n4);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n5, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n207, ZN => n5);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n209, A => n6, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n207, ZN => n6);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n209, A => n7, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n208, ZN => n7);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n8, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n208, ZN => n8);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n209, A => n9, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n208, ZN => n9);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n210, A => n10, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n208, ZN => n10);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n210, A => n11, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n209, ZN => n11);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n12, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n208, ZN => n12);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n210, A => n13, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n209, ZN => n13);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n210, A => n14, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n209, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n210, A => n15, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n209, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n210, A => n16, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n209, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n210, A => n17, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n209, ZN => n17);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n211, A => n18, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n209, ZN => n18);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n211, A => n19, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n208, ZN => n19);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n211, A => n20, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n208, ZN => n20);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n211, A => n21, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n208, ZN => n21);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n211, A => n22, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n208, ZN => n22);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n211, A => n23, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n208, ZN => n23);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n24, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n208, ZN => n24);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n211, A => n25, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n208, ZN => n25);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n211, A => n26, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n207, ZN => n26);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n211, A => n27, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n207, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n211, A => n28, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n207, ZN => n28);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n211, A => n29, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n207, ZN => n29);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n212, A => n30, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n207, ZN => n30);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n212, A => n31, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n207, ZN => n31);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n212, A => n32, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n207, ZN => n32);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n210, A => n33, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n207, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT7 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (6 
         downto 0);  data_out : out std_logic_vector (6 downto 0));

end REG_NBIT7;

architecture SYN_Behavioral of REG_NBIT7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n22, 
      n2, n3, n4, n5, n6, n7, n21, n26, n27, n28, n29 : std_logic;

begin
   
   reg_reg_6_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n29, Q => 
                           data_out(6), QN => n14);
   reg_reg_5_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n29, Q => 
                           data_out(5), QN => n13);
   reg_reg_4_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n29, Q => 
                           data_out(4), QN => n12);
   reg_reg_3_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n29, Q => 
                           data_out(3), QN => n11);
   reg_reg_2_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n29, Q => 
                           data_out(2), QN => n10);
   reg_reg_1_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n29, Q => 
                           data_out(1), QN => n9);
   reg_reg_0_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n29, Q => 
                           data_out(0), QN => n8);
   U2 : INV_X1 port map( A => reset, ZN => n29);
   U3 : BUF_X1 port map( A => n28, Z => n26);
   U4 : BUF_X1 port map( A => enable, Z => n28);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n26, A => n21, ZN => n15);
   U6 : NAND2_X1 port map( A1 => data_in(0), A2 => n26, ZN => n21);
   U7 : OAI21_X1 port map( B1 => n9, B2 => n26, A => n7, ZN => n16);
   U8 : NAND2_X1 port map( A1 => data_in(1), A2 => n26, ZN => n7);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n26, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => data_in(2), A2 => n26, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n11, B2 => n26, A => n5, ZN => n18);
   U12 : NAND2_X1 port map( A1 => data_in(3), A2 => n26, ZN => n5);
   U13 : OAI21_X1 port map( B1 => n12, B2 => n26, A => n4, ZN => n19);
   U14 : NAND2_X1 port map( A1 => data_in(4), A2 => n26, ZN => n4);
   U15 : OAI21_X1 port map( B1 => n13, B2 => n26, A => n3, ZN => n20);
   U16 : NAND2_X1 port map( A1 => data_in(5), A2 => n26, ZN => n3);
   U17 : OAI21_X1 port map( B1 => n14, B2 => n27, A => n2, ZN => n22);
   U18 : NAND2_X1 port map( A1 => n27, A2 => data_in(6), ZN => n2);
   U19 : BUF_X1 port map( A => n28, Z => n27);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_7 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_7;

architecture SYN_Behavioral of REG_NBIT32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n216, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n216, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n216, Q => 
                           data_out(29), QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n216, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n216, Q => 
                           data_out(27), QN => n147);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n216, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n216, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n216, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n218, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n218, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n218, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n217, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n218, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n218, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n218, Q => 
                           data_out(17), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n218, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n217, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n218, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n217, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n217, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n216, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n216, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n216, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n217, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n216, Q => 
                           data_out(0), QN => n174);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n217, Q => 
                           data_out(16), QN => n158);
   U2 : BUF_X1 port map( A => n207, Z => n215);
   U3 : BUF_X1 port map( A => n207, Z => n214);
   U4 : BUF_X1 port map( A => n215, Z => n209);
   U5 : BUF_X1 port map( A => n215, Z => n208);
   U6 : BUF_X1 port map( A => n215, Z => n210);
   U7 : BUF_X1 port map( A => n214, Z => n212);
   U8 : BUF_X1 port map( A => n214, Z => n211);
   U9 : BUF_X1 port map( A => n219, Z => n217);
   U10 : BUF_X1 port map( A => n219, Z => n216);
   U11 : BUF_X1 port map( A => n219, Z => n218);
   U12 : BUF_X1 port map( A => n214, Z => n213);
   U13 : INV_X1 port map( A => reset, ZN => n219);
   U14 : BUF_X1 port map( A => enable, Z => n207);
   U15 : OAI21_X1 port map( B1 => n158, B2 => n212, A => n18, ZN => n126);
   U16 : NAND2_X1 port map( A1 => data_in(16), A2 => n210, ZN => n18);
   U17 : OAI21_X1 port map( B1 => n174, B2 => n211, A => n2, ZN => n142);
   U18 : NAND2_X1 port map( A1 => n213, A2 => data_in(0), ZN => n2);
   U19 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n3, ZN => n141);
   U20 : NAND2_X1 port map( A1 => data_in(1), A2 => n208, ZN => n3);
   U21 : OAI21_X1 port map( B1 => n172, B2 => n210, A => n4, ZN => n140);
   U22 : NAND2_X1 port map( A1 => data_in(2), A2 => n208, ZN => n4);
   U23 : OAI21_X1 port map( B1 => n171, B2 => n211, A => n5, ZN => n139);
   U24 : NAND2_X1 port map( A1 => data_in(3), A2 => n208, ZN => n5);
   U25 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n6, ZN => n138);
   U26 : NAND2_X1 port map( A1 => data_in(4), A2 => n208, ZN => n6);
   U27 : OAI21_X1 port map( B1 => n169, B2 => n210, A => n7, ZN => n137);
   U28 : NAND2_X1 port map( A1 => data_in(5), A2 => n209, ZN => n7);
   U29 : OAI21_X1 port map( B1 => n168, B2 => n211, A => n8, ZN => n136);
   U30 : NAND2_X1 port map( A1 => data_in(6), A2 => n209, ZN => n8);
   U31 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n9, ZN => n135);
   U32 : NAND2_X1 port map( A1 => data_in(7), A2 => n209, ZN => n9);
   U33 : OAI21_X1 port map( B1 => n166, B2 => n211, A => n10, ZN => n134);
   U34 : NAND2_X1 port map( A1 => data_in(8), A2 => n209, ZN => n10);
   U35 : OAI21_X1 port map( B1 => n165, B2 => n211, A => n11, ZN => n133);
   U36 : NAND2_X1 port map( A1 => data_in(9), A2 => n210, ZN => n11);
   U37 : OAI21_X1 port map( B1 => n164, B2 => n211, A => n12, ZN => n132);
   U38 : NAND2_X1 port map( A1 => data_in(10), A2 => n209, ZN => n12);
   U39 : OAI21_X1 port map( B1 => n163, B2 => n211, A => n13, ZN => n131);
   U40 : NAND2_X1 port map( A1 => data_in(11), A2 => n210, ZN => n13);
   U41 : OAI21_X1 port map( B1 => n162, B2 => n211, A => n14, ZN => n130);
   U42 : NAND2_X1 port map( A1 => data_in(12), A2 => n210, ZN => n14);
   U43 : OAI21_X1 port map( B1 => n161, B2 => n211, A => n15, ZN => n129);
   U44 : NAND2_X1 port map( A1 => data_in(13), A2 => n210, ZN => n15);
   U45 : OAI21_X1 port map( B1 => n160, B2 => n211, A => n16, ZN => n128);
   U46 : NAND2_X1 port map( A1 => data_in(14), A2 => n210, ZN => n16);
   U47 : OAI21_X1 port map( B1 => n159, B2 => n211, A => n17, ZN => n127);
   U48 : NAND2_X1 port map( A1 => data_in(15), A2 => n210, ZN => n17);
   U49 : OAI21_X1 port map( B1 => n157, B2 => n212, A => n19, ZN => n125);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n209, ZN => n19);
   U51 : OAI21_X1 port map( B1 => n156, B2 => n212, A => n20, ZN => n124);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n209, ZN => n20);
   U53 : OAI21_X1 port map( B1 => n155, B2 => n212, A => n21, ZN => n123);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n209, ZN => n21);
   U55 : OAI21_X1 port map( B1 => n154, B2 => n212, A => n22, ZN => n122);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n209, ZN => n22);
   U57 : OAI21_X1 port map( B1 => n153, B2 => n212, A => n23, ZN => n121);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n209, ZN => n23);
   U59 : OAI21_X1 port map( B1 => n152, B2 => n212, A => n24, ZN => n120);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n209, ZN => n24);
   U61 : OAI21_X1 port map( B1 => n151, B2 => n212, A => n25, ZN => n119);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n209, ZN => n25);
   U63 : OAI21_X1 port map( B1 => n150, B2 => n212, A => n26, ZN => n118);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n208, ZN => n26);
   U65 : OAI21_X1 port map( B1 => n149, B2 => n212, A => n27, ZN => n117);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n208, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n148, B2 => n212, A => n28, ZN => n116);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n208, ZN => n28);
   U69 : OAI21_X1 port map( B1 => n147, B2 => n212, A => n29, ZN => n115);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n208, ZN => n29);
   U71 : OAI21_X1 port map( B1 => n146, B2 => n213, A => n30, ZN => n114);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n208, ZN => n30);
   U73 : OAI21_X1 port map( B1 => n145, B2 => n213, A => n31, ZN => n113);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n208, ZN => n31);
   U75 : OAI21_X1 port map( B1 => n144, B2 => n213, A => n32, ZN => n112);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n208, ZN => n32);
   U77 : OAI21_X1 port map( B1 => n143, B2 => n211, A => n33, ZN => n111);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n208, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_8 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_8;

architecture SYN_Behavioral of REG_NBIT32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n216, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n216, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n216, Q => 
                           data_out(29), QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n216, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n216, Q => 
                           data_out(27), QN => n147);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n216, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n216, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n216, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n216, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n217, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n217, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n217, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n217, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n217, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n217, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n217, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n217, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n217, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n218, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n218, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n218, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n218, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n218, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n218, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n218, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n218, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n174);
   U2 : BUF_X1 port map( A => n207, Z => n215);
   U3 : BUF_X1 port map( A => n207, Z => n214);
   U4 : BUF_X1 port map( A => n215, Z => n209);
   U5 : BUF_X1 port map( A => n215, Z => n208);
   U6 : BUF_X1 port map( A => n215, Z => n210);
   U7 : BUF_X1 port map( A => n214, Z => n212);
   U8 : BUF_X1 port map( A => n214, Z => n211);
   U9 : BUF_X1 port map( A => n219, Z => n217);
   U10 : BUF_X1 port map( A => n219, Z => n216);
   U11 : BUF_X1 port map( A => n219, Z => n218);
   U12 : BUF_X1 port map( A => n214, Z => n213);
   U13 : INV_X1 port map( A => reset, ZN => n219);
   U14 : BUF_X1 port map( A => enable, Z => n207);
   U15 : OAI21_X1 port map( B1 => n174, B2 => n211, A => n2, ZN => n142);
   U16 : NAND2_X1 port map( A1 => n213, A2 => data_in(0), ZN => n2);
   U17 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n3, ZN => n141);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n208, ZN => n3);
   U19 : OAI21_X1 port map( B1 => n172, B2 => n210, A => n4, ZN => n140);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n208, ZN => n4);
   U21 : OAI21_X1 port map( B1 => n171, B2 => n211, A => n5, ZN => n139);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n208, ZN => n5);
   U23 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n6, ZN => n138);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n208, ZN => n6);
   U25 : OAI21_X1 port map( B1 => n169, B2 => n210, A => n7, ZN => n137);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n209, ZN => n7);
   U27 : OAI21_X1 port map( B1 => n168, B2 => n211, A => n8, ZN => n136);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n209, ZN => n8);
   U29 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n9, ZN => n135);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n209, ZN => n9);
   U31 : OAI21_X1 port map( B1 => n166, B2 => n211, A => n10, ZN => n134);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n209, ZN => n10);
   U33 : OAI21_X1 port map( B1 => n165, B2 => n211, A => n11, ZN => n133);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n210, ZN => n11);
   U35 : OAI21_X1 port map( B1 => n164, B2 => n211, A => n12, ZN => n132);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n209, ZN => n12);
   U37 : OAI21_X1 port map( B1 => n163, B2 => n211, A => n13, ZN => n131);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n210, ZN => n13);
   U39 : OAI21_X1 port map( B1 => n162, B2 => n211, A => n14, ZN => n130);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n210, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n161, B2 => n211, A => n15, ZN => n129);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n210, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n160, B2 => n211, A => n16, ZN => n128);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n210, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n159, B2 => n211, A => n17, ZN => n127);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n210, ZN => n17);
   U47 : OAI21_X1 port map( B1 => n158, B2 => n212, A => n18, ZN => n126);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n210, ZN => n18);
   U49 : OAI21_X1 port map( B1 => n157, B2 => n212, A => n19, ZN => n125);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n209, ZN => n19);
   U51 : OAI21_X1 port map( B1 => n156, B2 => n212, A => n20, ZN => n124);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n209, ZN => n20);
   U53 : OAI21_X1 port map( B1 => n155, B2 => n212, A => n21, ZN => n123);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n209, ZN => n21);
   U55 : OAI21_X1 port map( B1 => n154, B2 => n212, A => n22, ZN => n122);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n209, ZN => n22);
   U57 : OAI21_X1 port map( B1 => n153, B2 => n212, A => n23, ZN => n121);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n209, ZN => n23);
   U59 : OAI21_X1 port map( B1 => n152, B2 => n212, A => n24, ZN => n120);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n209, ZN => n24);
   U61 : OAI21_X1 port map( B1 => n151, B2 => n212, A => n25, ZN => n119);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n209, ZN => n25);
   U63 : OAI21_X1 port map( B1 => n150, B2 => n212, A => n26, ZN => n118);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n208, ZN => n26);
   U65 : OAI21_X1 port map( B1 => n149, B2 => n212, A => n27, ZN => n117);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n208, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n148, B2 => n212, A => n28, ZN => n116);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n208, ZN => n28);
   U69 : OAI21_X1 port map( B1 => n147, B2 => n212, A => n29, ZN => n115);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n208, ZN => n29);
   U71 : OAI21_X1 port map( B1 => n146, B2 => n213, A => n30, ZN => n114);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n208, ZN => n30);
   U73 : OAI21_X1 port map( B1 => n145, B2 => n213, A => n31, ZN => n113);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n208, ZN => n31);
   U75 : OAI21_X1 port map( B1 => n144, B2 => n213, A => n32, ZN => n112);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n208, ZN => n32);
   U77 : OAI21_X1 port map( B1 => n143, B2 => n211, A => n33, ZN => n111);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n208, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_9 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_9;

architecture SYN_Behavioral of REG_NBIT32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n216, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n216, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n216, Q => 
                           data_out(29), QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n216, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n216, Q => 
                           data_out(27), QN => n147);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n216, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n216, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n216, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n216, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n217, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n216, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n217, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n217, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n217, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n217, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n217, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n217, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n217, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n216, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n218, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n218, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n218, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n218, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n218, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n218, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n218, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n218, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n174);
   U2 : BUF_X1 port map( A => n207, Z => n215);
   U3 : BUF_X1 port map( A => n207, Z => n214);
   U4 : BUF_X1 port map( A => n215, Z => n209);
   U5 : BUF_X1 port map( A => n215, Z => n210);
   U6 : BUF_X1 port map( A => n214, Z => n212);
   U7 : BUF_X1 port map( A => n214, Z => n211);
   U8 : BUF_X1 port map( A => n215, Z => n208);
   U9 : BUF_X1 port map( A => n219, Z => n217);
   U10 : BUF_X1 port map( A => n219, Z => n216);
   U11 : BUF_X1 port map( A => n219, Z => n218);
   U12 : BUF_X1 port map( A => n214, Z => n213);
   U13 : INV_X1 port map( A => reset, ZN => n219);
   U14 : BUF_X1 port map( A => enable, Z => n207);
   U15 : OAI21_X1 port map( B1 => n174, B2 => n211, A => n2, ZN => n142);
   U16 : NAND2_X1 port map( A1 => n213, A2 => data_in(0), ZN => n2);
   U17 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n3, ZN => n141);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n208, ZN => n3);
   U19 : OAI21_X1 port map( B1 => n172, B2 => n210, A => n4, ZN => n140);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n208, ZN => n4);
   U21 : OAI21_X1 port map( B1 => n171, B2 => n211, A => n5, ZN => n139);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n208, ZN => n5);
   U23 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n6, ZN => n138);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n208, ZN => n6);
   U25 : OAI21_X1 port map( B1 => n169, B2 => n210, A => n7, ZN => n137);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n209, ZN => n7);
   U27 : OAI21_X1 port map( B1 => n168, B2 => n211, A => n8, ZN => n136);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n209, ZN => n8);
   U29 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n9, ZN => n135);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n209, ZN => n9);
   U31 : OAI21_X1 port map( B1 => n166, B2 => n211, A => n10, ZN => n134);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n209, ZN => n10);
   U33 : OAI21_X1 port map( B1 => n165, B2 => n211, A => n11, ZN => n133);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n210, ZN => n11);
   U35 : OAI21_X1 port map( B1 => n164, B2 => n211, A => n12, ZN => n132);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n209, ZN => n12);
   U37 : OAI21_X1 port map( B1 => n163, B2 => n211, A => n13, ZN => n131);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n210, ZN => n13);
   U39 : OAI21_X1 port map( B1 => n162, B2 => n211, A => n14, ZN => n130);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n210, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n161, B2 => n211, A => n15, ZN => n129);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n210, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n160, B2 => n211, A => n16, ZN => n128);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n210, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n159, B2 => n211, A => n17, ZN => n127);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n210, ZN => n17);
   U47 : OAI21_X1 port map( B1 => n158, B2 => n212, A => n18, ZN => n126);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n210, ZN => n18);
   U49 : OAI21_X1 port map( B1 => n157, B2 => n212, A => n19, ZN => n125);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n209, ZN => n19);
   U51 : OAI21_X1 port map( B1 => n156, B2 => n212, A => n20, ZN => n124);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n209, ZN => n20);
   U53 : OAI21_X1 port map( B1 => n155, B2 => n212, A => n21, ZN => n123);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n209, ZN => n21);
   U55 : OAI21_X1 port map( B1 => n154, B2 => n212, A => n22, ZN => n122);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n209, ZN => n22);
   U57 : OAI21_X1 port map( B1 => n153, B2 => n212, A => n23, ZN => n121);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n209, ZN => n23);
   U59 : OAI21_X1 port map( B1 => n152, B2 => n212, A => n24, ZN => n120);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n209, ZN => n24);
   U61 : OAI21_X1 port map( B1 => n151, B2 => n212, A => n25, ZN => n119);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n209, ZN => n25);
   U63 : OAI21_X1 port map( B1 => n150, B2 => n212, A => n26, ZN => n118);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n208, ZN => n26);
   U65 : OAI21_X1 port map( B1 => n149, B2 => n212, A => n27, ZN => n117);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n208, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n148, B2 => n212, A => n28, ZN => n116);
   U68 : OAI21_X1 port map( B1 => n147, B2 => n212, A => n29, ZN => n115);
   U69 : NAND2_X1 port map( A1 => data_in(27), A2 => n208, ZN => n29);
   U70 : OAI21_X1 port map( B1 => n146, B2 => n213, A => n30, ZN => n114);
   U71 : NAND2_X1 port map( A1 => data_in(28), A2 => n208, ZN => n30);
   U72 : OAI21_X1 port map( B1 => n145, B2 => n213, A => n31, ZN => n113);
   U73 : NAND2_X1 port map( A1 => data_in(29), A2 => n208, ZN => n31);
   U74 : OAI21_X1 port map( B1 => n144, B2 => n213, A => n32, ZN => n112);
   U75 : NAND2_X1 port map( A1 => data_in(30), A2 => n208, ZN => n32);
   U76 : OAI21_X1 port map( B1 => n143, B2 => n211, A => n33, ZN => n111);
   U77 : NAND2_X1 port map( A1 => data_in(31), A2 => n208, ZN => n33);
   U78 : NAND2_X1 port map( A1 => data_in(26), A2 => n208, ZN => n28);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_10 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_10;

architecture SYN_Behavioral of REG_NBIT32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n216, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n216, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n216, Q => 
                           data_out(29), QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n216, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n216, Q => 
                           data_out(27), QN => n147);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n216, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n216, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n216, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n216, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n216, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n216, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n217, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n217, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n217, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n217, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n217, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n217, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n217, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n217, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n217, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n217, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n217, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n218, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n218, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n218, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n218, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n218, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n218, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n218, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n218, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n216, Q => 
                           data_out(0), QN => n174);
   U2 : BUF_X1 port map( A => n207, Z => n215);
   U3 : BUF_X1 port map( A => n207, Z => n214);
   U4 : BUF_X1 port map( A => n220, Z => n219);
   U5 : BUF_X1 port map( A => n215, Z => n209);
   U6 : BUF_X1 port map( A => n215, Z => n208);
   U7 : BUF_X1 port map( A => n215, Z => n210);
   U8 : BUF_X1 port map( A => n214, Z => n212);
   U9 : BUF_X1 port map( A => n214, Z => n211);
   U10 : BUF_X1 port map( A => n219, Z => n217);
   U11 : BUF_X1 port map( A => n219, Z => n216);
   U12 : BUF_X1 port map( A => n219, Z => n218);
   U13 : BUF_X1 port map( A => n214, Z => n213);
   U14 : INV_X1 port map( A => reset, ZN => n220);
   U15 : BUF_X1 port map( A => enable, Z => n207);
   U16 : OAI21_X1 port map( B1 => n174, B2 => n211, A => n2, ZN => n142);
   U17 : NAND2_X1 port map( A1 => n213, A2 => data_in(0), ZN => n2);
   U18 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n3, ZN => n141);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n208, ZN => n3);
   U20 : OAI21_X1 port map( B1 => n172, B2 => n210, A => n4, ZN => n140);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n208, ZN => n4);
   U22 : OAI21_X1 port map( B1 => n171, B2 => n211, A => n5, ZN => n139);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n208, ZN => n5);
   U24 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n6, ZN => n138);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n208, ZN => n6);
   U26 : OAI21_X1 port map( B1 => n169, B2 => n210, A => n7, ZN => n137);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n209, ZN => n7);
   U28 : OAI21_X1 port map( B1 => n168, B2 => n211, A => n8, ZN => n136);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n209, ZN => n8);
   U30 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n9, ZN => n135);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n209, ZN => n9);
   U32 : OAI21_X1 port map( B1 => n166, B2 => n211, A => n10, ZN => n134);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n209, ZN => n10);
   U34 : OAI21_X1 port map( B1 => n165, B2 => n211, A => n11, ZN => n133);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n210, ZN => n11);
   U36 : OAI21_X1 port map( B1 => n164, B2 => n211, A => n12, ZN => n132);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n209, ZN => n12);
   U38 : OAI21_X1 port map( B1 => n163, B2 => n211, A => n13, ZN => n131);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n210, ZN => n13);
   U40 : OAI21_X1 port map( B1 => n162, B2 => n211, A => n14, ZN => n130);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n210, ZN => n14);
   U42 : OAI21_X1 port map( B1 => n161, B2 => n211, A => n15, ZN => n129);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n210, ZN => n15);
   U44 : OAI21_X1 port map( B1 => n160, B2 => n211, A => n16, ZN => n128);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n210, ZN => n16);
   U46 : OAI21_X1 port map( B1 => n159, B2 => n211, A => n17, ZN => n127);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n210, ZN => n17);
   U48 : OAI21_X1 port map( B1 => n158, B2 => n212, A => n18, ZN => n126);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n210, ZN => n18);
   U50 : OAI21_X1 port map( B1 => n157, B2 => n212, A => n19, ZN => n125);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n209, ZN => n19);
   U52 : OAI21_X1 port map( B1 => n156, B2 => n212, A => n20, ZN => n124);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n209, ZN => n20);
   U54 : OAI21_X1 port map( B1 => n155, B2 => n212, A => n21, ZN => n123);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n209, ZN => n21);
   U56 : OAI21_X1 port map( B1 => n154, B2 => n212, A => n22, ZN => n122);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n209, ZN => n22);
   U58 : OAI21_X1 port map( B1 => n153, B2 => n212, A => n23, ZN => n121);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n209, ZN => n23);
   U60 : OAI21_X1 port map( B1 => n152, B2 => n212, A => n24, ZN => n120);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n209, ZN => n24);
   U62 : OAI21_X1 port map( B1 => n151, B2 => n212, A => n25, ZN => n119);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n209, ZN => n25);
   U64 : OAI21_X1 port map( B1 => n150, B2 => n212, A => n26, ZN => n118);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n208, ZN => n26);
   U66 : OAI21_X1 port map( B1 => n149, B2 => n212, A => n27, ZN => n117);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n208, ZN => n27);
   U68 : OAI21_X1 port map( B1 => n148, B2 => n212, A => n28, ZN => n116);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n208, ZN => n28);
   U70 : OAI21_X1 port map( B1 => n147, B2 => n212, A => n29, ZN => n115);
   U71 : NAND2_X1 port map( A1 => data_in(27), A2 => n208, ZN => n29);
   U72 : OAI21_X1 port map( B1 => n146, B2 => n213, A => n30, ZN => n114);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n208, ZN => n30);
   U74 : OAI21_X1 port map( B1 => n145, B2 => n213, A => n31, ZN => n113);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n208, ZN => n31);
   U76 : OAI21_X1 port map( B1 => n144, B2 => n213, A => n32, ZN => n112);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n208, ZN => n32);
   U78 : OAI21_X1 port map( B1 => n143, B2 => n211, A => n33, ZN => n111);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n208, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FFD_1;

architecture SYN_BEHAVIORAL of FFD_1 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n10, n11, n12, n13, n_1585 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n10, CK => CK, RN => n13, Q => Q_port, QN => 
                           n_1585);
   U2 : INV_X1 port map( A => n3, ZN => n10);
   U3 : INV_X1 port map( A => RESET, ZN => n13);
   U4 : INV_X1 port map( A => n11, ZN => n12);
   U5 : BUF_X1 port map( A => ENABLE, Z => n11);
   U6 : OAI22_X1 port map( A1 => n11, A2 => Q_port, B1 => D, B2 => n12, ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_11 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_11;

architecture SYN_Behavioral of REG_NBIT32_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n215, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n215, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n215, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n215, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n215, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n215, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n215, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n215, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n215, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n215, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n215, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n215, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n216, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n216, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n216, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n216, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n216, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n216, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n217, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n216, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n206, Z => n214);
   U3 : BUF_X1 port map( A => n206, Z => n213);
   U4 : BUF_X1 port map( A => n219, Z => n218);
   U5 : BUF_X1 port map( A => n214, Z => n208);
   U6 : BUF_X1 port map( A => n214, Z => n207);
   U7 : BUF_X1 port map( A => n214, Z => n209);
   U8 : BUF_X1 port map( A => n213, Z => n211);
   U9 : BUF_X1 port map( A => n213, Z => n210);
   U10 : BUF_X1 port map( A => n218, Z => n216);
   U11 : BUF_X1 port map( A => n218, Z => n215);
   U12 : BUF_X1 port map( A => n218, Z => n217);
   U13 : BUF_X1 port map( A => n213, Z => n212);
   U14 : INV_X1 port map( A => reset, ZN => n219);
   U15 : BUF_X1 port map( A => enable, Z => n206);
   U16 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n2, ZN => n141);
   U17 : NAND2_X1 port map( A1 => n212, A2 => data_in(0), ZN => n2);
   U18 : OAI21_X1 port map( B1 => n172, B2 => n209, A => n3, ZN => n140);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n207, ZN => n3);
   U20 : OAI21_X1 port map( B1 => n171, B2 => n209, A => n4, ZN => n139);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n207, ZN => n4);
   U22 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n5, ZN => n138);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n207, ZN => n5);
   U24 : OAI21_X1 port map( B1 => n169, B2 => n209, A => n6, ZN => n137);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n207, ZN => n6);
   U26 : OAI21_X1 port map( B1 => n168, B2 => n209, A => n7, ZN => n136);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n208, ZN => n7);
   U28 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n8, ZN => n135);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n208, ZN => n8);
   U30 : OAI21_X1 port map( B1 => n166, B2 => n209, A => n9, ZN => n134);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n208, ZN => n9);
   U32 : OAI21_X1 port map( B1 => n165, B2 => n210, A => n10, ZN => n133);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n208, ZN => n10);
   U34 : OAI21_X1 port map( B1 => n164, B2 => n210, A => n11, ZN => n132);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n209, ZN => n11);
   U36 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n12, ZN => n131);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n208, ZN => n12);
   U38 : OAI21_X1 port map( B1 => n162, B2 => n210, A => n13, ZN => n130);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n209, ZN => n13);
   U40 : OAI21_X1 port map( B1 => n161, B2 => n210, A => n14, ZN => n129);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n209, ZN => n14);
   U42 : OAI21_X1 port map( B1 => n160, B2 => n210, A => n15, ZN => n128);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n209, ZN => n15);
   U44 : OAI21_X1 port map( B1 => n159, B2 => n210, A => n16, ZN => n127);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n209, ZN => n16);
   U46 : OAI21_X1 port map( B1 => n158, B2 => n210, A => n17, ZN => n126);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n209, ZN => n17);
   U48 : OAI21_X1 port map( B1 => n157, B2 => n211, A => n18, ZN => n125);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n209, ZN => n18);
   U50 : OAI21_X1 port map( B1 => n156, B2 => n211, A => n19, ZN => n124);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n208, ZN => n19);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n211, A => n20, ZN => n123);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n208, ZN => n20);
   U54 : OAI21_X1 port map( B1 => n154, B2 => n211, A => n21, ZN => n122);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n208, ZN => n21);
   U56 : OAI21_X1 port map( B1 => n153, B2 => n211, A => n22, ZN => n121);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n208, ZN => n22);
   U58 : OAI21_X1 port map( B1 => n152, B2 => n211, A => n23, ZN => n120);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n208, ZN => n23);
   U60 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n24, ZN => n119);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n208, ZN => n24);
   U62 : OAI21_X1 port map( B1 => n150, B2 => n211, A => n25, ZN => n118);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n208, ZN => n25);
   U64 : OAI21_X1 port map( B1 => n149, B2 => n211, A => n26, ZN => n117);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n207, ZN => n26);
   U66 : OAI21_X1 port map( B1 => n148, B2 => n211, A => n27, ZN => n116);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n207, ZN => n27);
   U68 : OAI21_X1 port map( B1 => n147, B2 => n211, A => n28, ZN => n115);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n207, ZN => n28);
   U70 : OAI21_X1 port map( B1 => n146, B2 => n211, A => n29, ZN => n114);
   U71 : NAND2_X1 port map( A1 => data_in(27), A2 => n207, ZN => n29);
   U72 : OAI21_X1 port map( B1 => n145, B2 => n212, A => n30, ZN => n113);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n207, ZN => n30);
   U74 : OAI21_X1 port map( B1 => n144, B2 => n212, A => n31, ZN => n112);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n207, ZN => n31);
   U76 : OAI21_X1 port map( B1 => n143, B2 => n212, A => n32, ZN => n111);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n207, ZN => n32);
   U78 : OAI21_X1 port map( B1 => n142, B2 => n210, A => n33, ZN => n110);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n207, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_12 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_12;

architecture SYN_Behavioral of REG_NBIT32_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n44, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n45, n46, n167, n168, n169, n170, n171, n172, n173, n174, n175,
      n176, n177, n178, n179, n180 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n176, Q => 
                           data_out(31), QN => n127);
   reg_reg_30_inst : DFFR_X1 port map( D => n96, CK => clk, RN => n176, Q => 
                           data_out(30), QN => n128);
   reg_reg_29_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n176, Q => 
                           data_out(29), QN => n129);
   reg_reg_28_inst : DFFR_X1 port map( D => n98, CK => clk, RN => n176, Q => 
                           data_out(28), QN => n130);
   reg_reg_27_inst : DFFR_X1 port map( D => n99, CK => clk, RN => n177, Q => 
                           data_out(27), QN => n131);
   reg_reg_26_inst : DFFR_X1 port map( D => n100, CK => clk, RN => n177, Q => 
                           data_out(26), QN => n132);
   reg_reg_25_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n177, Q => 
                           data_out(25), QN => n133);
   reg_reg_24_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n177, Q => 
                           data_out(24), QN => n134);
   reg_reg_23_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n177, Q => 
                           data_out(23), QN => n135);
   reg_reg_22_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n177, Q => 
                           data_out(22), QN => n136);
   reg_reg_21_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n177, Q => 
                           data_out(21), QN => n137);
   reg_reg_20_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n177, Q => 
                           data_out(20), QN => n138);
   reg_reg_19_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n177, Q => 
                           data_out(19), QN => n139);
   reg_reg_18_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n177, Q => 
                           data_out(18), QN => n140);
   reg_reg_17_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n177, Q => 
                           data_out(17), QN => n141);
   reg_reg_16_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n177, Q => 
                           data_out(16), QN => n142);
   reg_reg_15_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n178, Q => 
                           data_out(15), QN => n143);
   reg_reg_14_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n178, Q => 
                           data_out(14), QN => n144);
   reg_reg_13_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n178, Q => 
                           data_out(13), QN => n145);
   reg_reg_12_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n178, Q => 
                           data_out(12), QN => n146);
   reg_reg_11_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n178, Q => 
                           data_out(11), QN => n46);
   reg_reg_10_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n178, Q => 
                           data_out(10), QN => n45);
   reg_reg_9_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n178, Q => 
                           data_out(9), QN => n43);
   reg_reg_8_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n178, Q => 
                           data_out(8), QN => n42);
   reg_reg_7_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n176, Q => 
                           data_out(7), QN => n41);
   reg_reg_6_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n176, Q => 
                           data_out(6), QN => n40);
   reg_reg_5_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n176, Q => 
                           data_out(5), QN => n39);
   reg_reg_4_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n176, Q => 
                           data_out(4), QN => n38);
   reg_reg_3_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n176, Q => 
                           data_out(3), QN => n37);
   reg_reg_2_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n176, Q => 
                           data_out(2), QN => n36);
   reg_reg_1_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n176, Q => 
                           data_out(1), QN => n35);
   reg_reg_0_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n176, Q => 
                           data_out(0), QN => n34);
   U2 : BUF_X1 port map( A => n167, Z => n175);
   U3 : BUF_X1 port map( A => n167, Z => n174);
   U4 : BUF_X1 port map( A => n180, Z => n179);
   U5 : BUF_X1 port map( A => n175, Z => n169);
   U6 : BUF_X1 port map( A => n175, Z => n168);
   U7 : BUF_X1 port map( A => n175, Z => n170);
   U8 : BUF_X1 port map( A => n174, Z => n172);
   U9 : BUF_X1 port map( A => n174, Z => n171);
   U10 : BUF_X1 port map( A => n179, Z => n177);
   U11 : BUF_X1 port map( A => n179, Z => n176);
   U12 : BUF_X1 port map( A => n179, Z => n178);
   U13 : BUF_X1 port map( A => n174, Z => n173);
   U14 : INV_X1 port map( A => reset, ZN => n180);
   U15 : BUF_X1 port map( A => enable, Z => n167);
   U16 : OAI21_X1 port map( B1 => n34, B2 => n170, A => n7, ZN => n126);
   U17 : NAND2_X1 port map( A1 => data_in(0), A2 => n169, ZN => n7);
   U18 : OAI21_X1 port map( B1 => n35, B2 => n171, A => n8, ZN => n125);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n169, ZN => n8);
   U20 : OAI21_X1 port map( B1 => n36, B2 => n170, A => n9, ZN => n124);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n169, ZN => n9);
   U22 : OAI21_X1 port map( B1 => n37, B2 => n171, A => n10, ZN => n123);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n169, ZN => n10);
   U24 : OAI21_X1 port map( B1 => n38, B2 => n171, A => n11, ZN => n122);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n170, ZN => n11);
   U26 : OAI21_X1 port map( B1 => n39, B2 => n171, A => n12, ZN => n121);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n169, ZN => n12);
   U28 : OAI21_X1 port map( B1 => n40, B2 => n171, A => n13, ZN => n120);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n170, ZN => n13);
   U30 : OAI21_X1 port map( B1 => n41, B2 => n171, A => n14, ZN => n119);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n170, ZN => n14);
   U32 : OAI21_X1 port map( B1 => n42, B2 => n171, A => n15, ZN => n118);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n170, ZN => n15);
   U34 : OAI21_X1 port map( B1 => n43, B2 => n171, A => n16, ZN => n117);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n170, ZN => n16);
   U36 : OAI21_X1 port map( B1 => n45, B2 => n171, A => n17, ZN => n116);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n170, ZN => n17);
   U38 : OAI21_X1 port map( B1 => n46, B2 => n172, A => n18, ZN => n115);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n170, ZN => n18);
   U40 : OAI21_X1 port map( B1 => n146, B2 => n172, A => n19, ZN => n114);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n169, ZN => n19);
   U42 : OAI21_X1 port map( B1 => n145, B2 => n172, A => n20, ZN => n113);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n169, ZN => n20);
   U44 : OAI21_X1 port map( B1 => n144, B2 => n172, A => n21, ZN => n112);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n169, ZN => n21);
   U46 : OAI21_X1 port map( B1 => n143, B2 => n172, A => n22, ZN => n111);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n169, ZN => n22);
   U48 : OAI21_X1 port map( B1 => n142, B2 => n172, A => n23, ZN => n110);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n169, ZN => n23);
   U50 : OAI21_X1 port map( B1 => n141, B2 => n172, A => n24, ZN => n109);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n169, ZN => n24);
   U52 : OAI21_X1 port map( B1 => n140, B2 => n172, A => n25, ZN => n108);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n169, ZN => n25);
   U54 : OAI21_X1 port map( B1 => n139, B2 => n172, A => n26, ZN => n107);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n168, ZN => n26);
   U56 : OAI21_X1 port map( B1 => n138, B2 => n172, A => n27, ZN => n106);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n168, ZN => n27);
   U58 : OAI21_X1 port map( B1 => n137, B2 => n172, A => n28, ZN => n105);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n168, ZN => n28);
   U60 : OAI21_X1 port map( B1 => n136, B2 => n172, A => n29, ZN => n104);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n168, ZN => n29);
   U62 : OAI21_X1 port map( B1 => n135, B2 => n173, A => n30, ZN => n103);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n168, ZN => n30);
   U64 : OAI21_X1 port map( B1 => n134, B2 => n173, A => n31, ZN => n102);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n168, ZN => n31);
   U66 : OAI21_X1 port map( B1 => n133, B2 => n173, A => n32, ZN => n101);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n168, ZN => n32);
   U68 : OAI21_X1 port map( B1 => n132, B2 => n171, A => n33, ZN => n100);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n168, ZN => n33);
   U70 : OAI21_X1 port map( B1 => n131, B2 => n171, A => n2, ZN => n99);
   U71 : NAND2_X1 port map( A1 => n173, A2 => data_in(27), ZN => n2);
   U72 : OAI21_X1 port map( B1 => n130, B2 => n170, A => n3, ZN => n98);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n168, ZN => n3);
   U74 : OAI21_X1 port map( B1 => n129, B2 => n170, A => n4, ZN => n97);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n168, ZN => n4);
   U76 : OAI21_X1 port map( B1 => n128, B2 => n171, A => n5, ZN => n96);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n168, ZN => n5);
   U78 : OAI21_X1 port map( B1 => n127, B2 => n170, A => n6, ZN => n44);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n168, ZN => n6);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FFD_0;

architecture SYN_BEHAVIORAL of FFD_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n2, n3, n5 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n5, Q => Q, QN => n3);
   U2 : INV_X1 port map( A => RESET, ZN => n5);
   U3 : OAI21_X1 port map( B1 => n3, B2 => ENABLE, A => n2, ZN => n4);
   U4 : NAND2_X1 port map( A1 => ENABLE, A2 => D, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_13 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_13;

architecture SYN_Behavioral of REG_NBIT32_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n211, Q => 
                           data_out(31), QN => n140);
   reg_reg_30_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n211, Q => 
                           data_out(30), QN => n141);
   reg_reg_29_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n212, Q => 
                           data_out(29), QN => n142);
   reg_reg_28_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n212, Q => 
                           data_out(28), QN => n143);
   reg_reg_27_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n212, Q => 
                           data_out(27), QN => n144);
   reg_reg_26_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n211, Q => 
                           data_out(26), QN => n34);
   reg_reg_25_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n212, Q => 
                           data_out(25), QN => n145);
   reg_reg_24_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n212, Q => 
                           data_out(24), QN => n146);
   reg_reg_23_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n211, Q => 
                           data_out(23), QN => n147);
   reg_reg_22_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n212, Q => 
                           data_out(22), QN => n148);
   reg_reg_21_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n211, Q => 
                           data_out(21), QN => n149);
   reg_reg_20_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n212, Q => 
                           data_out(20), QN => n150);
   reg_reg_19_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n212, Q => 
                           data_out(19), QN => n151);
   reg_reg_18_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n213, Q => 
                           data_out(18), QN => n152);
   reg_reg_17_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n212, Q => 
                           data_out(17), QN => n153);
   reg_reg_16_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n212, Q => 
                           data_out(16), QN => n154);
   reg_reg_15_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n213, Q => 
                           data_out(15), QN => n155);
   reg_reg_14_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n213, Q => 
                           data_out(14), QN => n156);
   reg_reg_13_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n213, Q => 
                           data_out(13), QN => n157);
   reg_reg_12_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n212, Q => 
                           data_out(12), QN => n158);
   reg_reg_11_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n213, Q => 
                           data_out(11), QN => n159);
   reg_reg_10_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n213, Q => 
                           data_out(10), QN => n160);
   reg_reg_9_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n213, Q => 
                           data_out(9), QN => n161);
   reg_reg_8_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n213, Q => 
                           data_out(8), QN => n162);
   reg_reg_7_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n212, Q => 
                           data_out(7), QN => n163);
   reg_reg_6_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n211, Q => 
                           data_out(6), QN => n164);
   reg_reg_5_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n211, Q => 
                           data_out(5), QN => n165);
   reg_reg_4_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n211, Q => 
                           data_out(4), QN => n166);
   reg_reg_3_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n211, Q => 
                           data_out(3), QN => n167);
   reg_reg_2_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n211, Q => 
                           data_out(2), QN => n168);
   reg_reg_1_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n211, Q => 
                           data_out(1), QN => n169);
   reg_reg_0_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n211, Q => 
                           data_out(0), QN => n170);
   U2 : BUF_X1 port map( A => n202, Z => n210);
   U3 : BUF_X1 port map( A => n202, Z => n209);
   U4 : BUF_X1 port map( A => n215, Z => n214);
   U5 : BUF_X1 port map( A => n210, Z => n205);
   U6 : BUF_X1 port map( A => n209, Z => n207);
   U7 : BUF_X1 port map( A => n209, Z => n206);
   U8 : BUF_X1 port map( A => n210, Z => n203);
   U9 : BUF_X1 port map( A => n210, Z => n204);
   U10 : BUF_X1 port map( A => n214, Z => n212);
   U11 : BUF_X1 port map( A => n214, Z => n211);
   U12 : BUF_X1 port map( A => n214, Z => n213);
   U13 : BUF_X1 port map( A => n209, Z => n208);
   U14 : INV_X1 port map( A => reset, ZN => n215);
   U15 : BUF_X1 port map( A => enable, Z => n202);
   U16 : OAI21_X1 port map( B1 => n170, B2 => n206, A => n2, ZN => n139);
   U17 : NAND2_X1 port map( A1 => n208, A2 => data_in(0), ZN => n2);
   U18 : OAI21_X1 port map( B1 => n169, B2 => n205, A => n3, ZN => n138);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n203, ZN => n3);
   U20 : OAI21_X1 port map( B1 => n168, B2 => n205, A => n4, ZN => n137);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n203, ZN => n4);
   U22 : OAI21_X1 port map( B1 => n167, B2 => n206, A => n5, ZN => n136);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n203, ZN => n5);
   U24 : OAI21_X1 port map( B1 => n166, B2 => n205, A => n6, ZN => n135);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n203, ZN => n6);
   U26 : OAI21_X1 port map( B1 => n165, B2 => n205, A => n7, ZN => n134);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n204, ZN => n7);
   U28 : OAI21_X1 port map( B1 => n164, B2 => n206, A => n8, ZN => n133);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n204, ZN => n8);
   U30 : OAI21_X1 port map( B1 => n163, B2 => n205, A => n9, ZN => n132);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n204, ZN => n9);
   U32 : OAI21_X1 port map( B1 => n162, B2 => n206, A => n10, ZN => n131);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n204, ZN => n10);
   U34 : OAI21_X1 port map( B1 => n161, B2 => n206, A => n11, ZN => n130);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n205, ZN => n11);
   U36 : OAI21_X1 port map( B1 => n160, B2 => n206, A => n12, ZN => n129);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n204, ZN => n12);
   U38 : OAI21_X1 port map( B1 => n159, B2 => n206, A => n13, ZN => n128);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n205, ZN => n13);
   U40 : OAI21_X1 port map( B1 => n158, B2 => n206, A => n14, ZN => n127);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n205, ZN => n14);
   U42 : OAI21_X1 port map( B1 => n157, B2 => n206, A => n15, ZN => n126);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n205, ZN => n15);
   U44 : OAI21_X1 port map( B1 => n156, B2 => n206, A => n16, ZN => n125);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n205, ZN => n16);
   U46 : OAI21_X1 port map( B1 => n155, B2 => n206, A => n17, ZN => n124);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n205, ZN => n17);
   U48 : OAI21_X1 port map( B1 => n154, B2 => n207, A => n18, ZN => n123);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n205, ZN => n18);
   U50 : OAI21_X1 port map( B1 => n153, B2 => n207, A => n19, ZN => n122);
   U51 : OAI21_X1 port map( B1 => n152, B2 => n207, A => n20, ZN => n121);
   U52 : OAI21_X1 port map( B1 => n151, B2 => n207, A => n21, ZN => n120);
   U53 : OAI21_X1 port map( B1 => n150, B2 => n207, A => n22, ZN => n119);
   U54 : OAI21_X1 port map( B1 => n149, B2 => n207, A => n23, ZN => n118);
   U55 : OAI21_X1 port map( B1 => n148, B2 => n207, A => n24, ZN => n117);
   U56 : OAI21_X1 port map( B1 => n147, B2 => n207, A => n25, ZN => n116);
   U57 : NAND2_X1 port map( A1 => data_in(23), A2 => n204, ZN => n25);
   U58 : OAI21_X1 port map( B1 => n146, B2 => n207, A => n26, ZN => n115);
   U59 : NAND2_X1 port map( A1 => data_in(24), A2 => n203, ZN => n26);
   U60 : OAI21_X1 port map( B1 => n145, B2 => n207, A => n27, ZN => n114);
   U61 : OAI21_X1 port map( B1 => n34, B2 => n207, A => n28, ZN => n113);
   U62 : OAI21_X1 port map( B1 => n144, B2 => n207, A => n29, ZN => n112);
   U63 : OAI21_X1 port map( B1 => n143, B2 => n208, A => n30, ZN => n111);
   U64 : OAI21_X1 port map( B1 => n142, B2 => n208, A => n31, ZN => n110);
   U65 : NAND2_X1 port map( A1 => data_in(29), A2 => n203, ZN => n31);
   U66 : OAI21_X1 port map( B1 => n141, B2 => n208, A => n32, ZN => n109);
   U67 : NAND2_X1 port map( A1 => data_in(30), A2 => n203, ZN => n32);
   U68 : OAI21_X1 port map( B1 => n140, B2 => n206, A => n33, ZN => n108);
   U69 : NAND2_X1 port map( A1 => data_in(31), A2 => n203, ZN => n33);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n203, ZN => n29);
   U71 : NAND2_X1 port map( A1 => data_in(19), A2 => n204, ZN => n21);
   U72 : NAND2_X1 port map( A1 => data_in(17), A2 => n204, ZN => n19);
   U73 : NAND2_X1 port map( A1 => data_in(22), A2 => n204, ZN => n24);
   U74 : NAND2_X1 port map( A1 => data_in(25), A2 => n203, ZN => n27);
   U75 : NAND2_X1 port map( A1 => data_in(20), A2 => n204, ZN => n22);
   U76 : NAND2_X1 port map( A1 => data_in(21), A2 => n204, ZN => n23);
   U77 : NAND2_X1 port map( A1 => data_in(18), A2 => n204, ZN => n20);
   U78 : NAND2_X1 port map( A1 => data_in(26), A2 => n203, ZN => n28);
   U79 : NAND2_X1 port map( A1 => data_in(28), A2 => n203, ZN => n30);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_14 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_14;

architecture SYN_Behavioral of REG_NBIT32_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n215, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n215, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n215, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n215, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n215, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n215, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n215, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n215, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n215, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n215, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n215, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n216, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n216, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n216, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n215, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n217, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n217, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n217, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n217, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n216, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n216, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n216, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n216, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n206, Z => n214);
   U3 : BUF_X1 port map( A => n206, Z => n213);
   U4 : BUF_X1 port map( A => n219, Z => n218);
   U5 : BUF_X1 port map( A => n214, Z => n208);
   U6 : BUF_X1 port map( A => n214, Z => n207);
   U7 : BUF_X1 port map( A => n214, Z => n209);
   U8 : BUF_X1 port map( A => n213, Z => n211);
   U9 : BUF_X1 port map( A => n213, Z => n210);
   U10 : BUF_X1 port map( A => n218, Z => n216);
   U11 : BUF_X1 port map( A => n218, Z => n215);
   U12 : BUF_X1 port map( A => n218, Z => n217);
   U13 : BUF_X1 port map( A => n213, Z => n212);
   U14 : INV_X1 port map( A => reset, ZN => n219);
   U15 : BUF_X1 port map( A => enable, Z => n206);
   U16 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n2, ZN => n141);
   U17 : NAND2_X1 port map( A1 => n212, A2 => data_in(0), ZN => n2);
   U18 : OAI21_X1 port map( B1 => n172, B2 => n209, A => n3, ZN => n140);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n207, ZN => n3);
   U20 : OAI21_X1 port map( B1 => n171, B2 => n209, A => n4, ZN => n139);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n207, ZN => n4);
   U22 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n5, ZN => n138);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n207, ZN => n5);
   U24 : OAI21_X1 port map( B1 => n169, B2 => n209, A => n6, ZN => n137);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n207, ZN => n6);
   U26 : OAI21_X1 port map( B1 => n168, B2 => n209, A => n7, ZN => n136);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n208, ZN => n7);
   U28 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n8, ZN => n135);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n208, ZN => n8);
   U30 : OAI21_X1 port map( B1 => n166, B2 => n209, A => n9, ZN => n134);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n208, ZN => n9);
   U32 : OAI21_X1 port map( B1 => n165, B2 => n210, A => n10, ZN => n133);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n208, ZN => n10);
   U34 : OAI21_X1 port map( B1 => n164, B2 => n210, A => n11, ZN => n132);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n209, ZN => n11);
   U36 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n12, ZN => n131);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n208, ZN => n12);
   U38 : OAI21_X1 port map( B1 => n162, B2 => n210, A => n13, ZN => n130);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n209, ZN => n13);
   U40 : OAI21_X1 port map( B1 => n161, B2 => n210, A => n14, ZN => n129);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n209, ZN => n14);
   U42 : OAI21_X1 port map( B1 => n160, B2 => n210, A => n15, ZN => n128);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n209, ZN => n15);
   U44 : OAI21_X1 port map( B1 => n159, B2 => n210, A => n16, ZN => n127);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n209, ZN => n16);
   U46 : OAI21_X1 port map( B1 => n158, B2 => n210, A => n17, ZN => n126);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n209, ZN => n17);
   U48 : OAI21_X1 port map( B1 => n157, B2 => n211, A => n18, ZN => n125);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n209, ZN => n18);
   U50 : OAI21_X1 port map( B1 => n156, B2 => n211, A => n19, ZN => n124);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n208, ZN => n19);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n211, A => n20, ZN => n123);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n208, ZN => n20);
   U54 : OAI21_X1 port map( B1 => n154, B2 => n211, A => n21, ZN => n122);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n208, ZN => n21);
   U56 : OAI21_X1 port map( B1 => n153, B2 => n211, A => n22, ZN => n121);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n208, ZN => n22);
   U58 : OAI21_X1 port map( B1 => n152, B2 => n211, A => n23, ZN => n120);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n208, ZN => n23);
   U60 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n24, ZN => n119);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n208, ZN => n24);
   U62 : OAI21_X1 port map( B1 => n150, B2 => n211, A => n25, ZN => n118);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n208, ZN => n25);
   U64 : OAI21_X1 port map( B1 => n149, B2 => n211, A => n26, ZN => n117);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n207, ZN => n26);
   U66 : OAI21_X1 port map( B1 => n148, B2 => n211, A => n27, ZN => n116);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n207, ZN => n27);
   U68 : OAI21_X1 port map( B1 => n147, B2 => n211, A => n28, ZN => n115);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n207, ZN => n28);
   U70 : OAI21_X1 port map( B1 => n146, B2 => n211, A => n29, ZN => n114);
   U71 : NAND2_X1 port map( A1 => data_in(27), A2 => n207, ZN => n29);
   U72 : OAI21_X1 port map( B1 => n145, B2 => n212, A => n30, ZN => n113);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n207, ZN => n30);
   U74 : OAI21_X1 port map( B1 => n144, B2 => n212, A => n31, ZN => n112);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n207, ZN => n31);
   U76 : OAI21_X1 port map( B1 => n143, B2 => n212, A => n32, ZN => n111);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n207, ZN => n32);
   U78 : OAI21_X1 port map( B1 => n142, B2 => n210, A => n33, ZN => n110);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n207, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_15 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_15;

architecture SYN_Behavioral of REG_NBIT32_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n215, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n215, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n215, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n215, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n215, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n215, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n215, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n215, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n215, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n215, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n215, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n215, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n216, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n216, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n216, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n216, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n216, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n216, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n216, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n216, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n216, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n216, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n217, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n217, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n217, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n206, Z => n214);
   U3 : BUF_X1 port map( A => n206, Z => n213);
   U4 : BUF_X1 port map( A => n214, Z => n208);
   U5 : BUF_X1 port map( A => n214, Z => n207);
   U6 : BUF_X1 port map( A => n214, Z => n209);
   U7 : BUF_X1 port map( A => n213, Z => n211);
   U8 : BUF_X1 port map( A => n213, Z => n210);
   U9 : BUF_X1 port map( A => n218, Z => n216);
   U10 : BUF_X1 port map( A => n218, Z => n215);
   U11 : BUF_X1 port map( A => n218, Z => n217);
   U12 : BUF_X1 port map( A => n213, Z => n212);
   U13 : INV_X1 port map( A => reset, ZN => n218);
   U14 : BUF_X1 port map( A => enable, Z => n206);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n2, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n212, A2 => data_in(0), ZN => n2);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n209, A => n3, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n207, ZN => n3);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n209, A => n4, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n207, ZN => n4);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n5, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n207, ZN => n5);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n209, A => n6, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n207, ZN => n6);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n209, A => n7, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n208, ZN => n7);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n8, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n208, ZN => n8);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n209, A => n9, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n208, ZN => n9);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n210, A => n10, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n208, ZN => n10);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n210, A => n11, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n209, ZN => n11);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n12, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n208, ZN => n12);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n210, A => n13, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n209, ZN => n13);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n210, A => n14, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n209, ZN => n14);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n210, A => n15, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n209, ZN => n15);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n210, A => n16, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n209, ZN => n16);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n210, A => n17, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n209, ZN => n17);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n211, A => n18, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n209, ZN => n18);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n211, A => n19, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n208, ZN => n19);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n211, A => n20, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n208, ZN => n20);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n211, A => n21, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n208, ZN => n21);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n211, A => n22, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n208, ZN => n22);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n211, A => n23, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n208, ZN => n23);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n24, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n208, ZN => n24);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n211, A => n25, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n208, ZN => n25);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n211, A => n26, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n207, ZN => n26);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n211, A => n27, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n207, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n211, A => n28, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n207, ZN => n28);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n211, A => n29, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n207, ZN => n29);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n212, A => n30, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n207, ZN => n30);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n212, A => n31, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n207, ZN => n31);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n212, A => n32, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n207, ZN => n32);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n210, A => n33, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n207, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_16 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_16;

architecture SYN_Behavioral of REG_NBIT32_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n60, n61, n62, n63, n64, n92, n93, n94, n95, n96, n97, n98, n99, n100
      , n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
      n163 : std_logic;

begin
   
   reg_reg_30_inst : DFFR_X1 port map( D => n61, CK => clk, RN => n160, Q => 
                           data_out(30), QN => n48);
   reg_reg_29_inst : DFFR_X1 port map( D => n62, CK => clk, RN => n160, Q => 
                           data_out(29), QN => n47);
   reg_reg_28_inst : DFFR_X1 port map( D => n63, CK => clk, RN => n160, Q => 
                           data_out(28), QN => n46);
   reg_reg_27_inst : DFFR_X1 port map( D => n64, CK => clk, RN => n161, Q => 
                           data_out(27), QN => n45);
   reg_reg_26_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n161, Q => 
                           data_out(26), QN => n44);
   reg_reg_25_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n161, Q => 
                           data_out(25), QN => n43);
   reg_reg_24_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n161, Q => 
                           data_out(24), QN => n42);
   reg_reg_23_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n160, Q => 
                           data_out(23), QN => n41);
   reg_reg_22_inst : DFFR_X1 port map( D => n96, CK => clk, RN => n160, Q => 
                           data_out(22), QN => n40);
   reg_reg_21_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n160, Q => 
                           data_out(21), QN => n39);
   reg_reg_20_inst : DFFR_X1 port map( D => n98, CK => clk, RN => n160, Q => 
                           data_out(20), QN => n38);
   reg_reg_19_inst : DFFR_X1 port map( D => n99, CK => clk, RN => n160, Q => 
                           data_out(19), QN => n37);
   reg_reg_18_inst : DFFR_X1 port map( D => n100, CK => clk, RN => n160, Q => 
                           data_out(18), QN => n36);
   reg_reg_17_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n160, Q => 
                           data_out(17), QN => n35);
   reg_reg_16_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n160, Q => 
                           data_out(16), QN => n34);
   reg_reg_15_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n161, Q => 
                           data_out(15), QN => n119);
   reg_reg_14_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n161, Q => 
                           data_out(14), QN => n120);
   reg_reg_13_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n161, Q => 
                           data_out(13), QN => n121);
   reg_reg_12_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n161, Q => 
                           data_out(12), QN => n122);
   reg_reg_11_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n162, Q => 
                           data_out(11), QN => n123);
   reg_reg_10_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n162, Q => 
                           data_out(10), QN => n124);
   reg_reg_9_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n162, Q => 
                           data_out(9), QN => n125);
   reg_reg_8_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n162, Q => 
                           data_out(8), QN => n126);
   reg_reg_7_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n162, Q => 
                           data_out(7), QN => n127);
   reg_reg_6_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n162, Q => 
                           data_out(6), QN => n128);
   reg_reg_5_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n162, Q => 
                           data_out(5), QN => n129);
   reg_reg_4_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n162, Q => 
                           data_out(4), QN => n130);
   reg_reg_3_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n161, Q => 
                           data_out(3), QN => n131);
   reg_reg_2_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n161, Q => 
                           data_out(2), QN => n132);
   reg_reg_1_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n161, Q => 
                           data_out(1), QN => n133);
   reg_reg_0_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n161, Q => 
                           data_out(0), QN => n134);
   reg_reg_31_inst : DFFR_X1 port map( D => n60, CK => clk, RN => n160, Q => 
                           data_out(31), QN => n49);
   U2 : BUF_X1 port map( A => n151, Z => n159);
   U3 : BUF_X1 port map( A => n151, Z => n158);
   U4 : BUF_X1 port map( A => n159, Z => n153);
   U5 : BUF_X1 port map( A => n159, Z => n152);
   U6 : BUF_X1 port map( A => n159, Z => n154);
   U7 : BUF_X1 port map( A => n158, Z => n157);
   U8 : BUF_X1 port map( A => n158, Z => n156);
   U9 : BUF_X1 port map( A => n158, Z => n155);
   U10 : BUF_X1 port map( A => n163, Z => n161);
   U11 : BUF_X1 port map( A => n163, Z => n160);
   U12 : BUF_X1 port map( A => n163, Z => n162);
   U13 : INV_X1 port map( A => reset, ZN => n163);
   U14 : BUF_X1 port map( A => enable, Z => n151);
   U15 : OAI21_X1 port map( B1 => n48, B2 => n155, A => n13, ZN => n61);
   U16 : NAND2_X1 port map( A1 => data_in(30), A2 => n154, ZN => n13);
   U17 : OAI21_X1 port map( B1 => n45, B2 => n155, A => n10, ZN => n64);
   U18 : OAI21_X1 port map( B1 => n47, B2 => n155, A => n12, ZN => n62);
   U19 : NAND2_X1 port map( A1 => data_in(29), A2 => n153, ZN => n12);
   U20 : OAI21_X1 port map( B1 => n44, B2 => n154, A => n9, ZN => n92);
   U21 : NAND2_X1 port map( A1 => data_in(26), A2 => n153, ZN => n9);
   U22 : OAI21_X1 port map( B1 => n119, B2 => n157, A => n30, ZN => n103);
   U23 : NAND2_X1 port map( A1 => data_in(15), A2 => n152, ZN => n30);
   U24 : OAI21_X1 port map( B1 => n41, B2 => n154, A => n6, ZN => n95);
   U25 : NAND2_X1 port map( A1 => data_in(23), A2 => n152, ZN => n6);
   U26 : OAI21_X1 port map( B1 => n46, B2 => n155, A => n11, ZN => n63);
   U27 : NAND2_X1 port map( A1 => data_in(28), A2 => n154, ZN => n11);
   U28 : OAI21_X1 port map( B1 => n43, B2 => n155, A => n8, ZN => n93);
   U29 : NAND2_X1 port map( A1 => data_in(25), A2 => n153, ZN => n8);
   U30 : OAI21_X1 port map( B1 => n120, B2 => n156, A => n29, ZN => n104);
   U31 : NAND2_X1 port map( A1 => data_in(14), A2 => n152, ZN => n29);
   U32 : OAI21_X1 port map( B1 => n40, B2 => n155, A => n5, ZN => n96);
   U33 : NAND2_X1 port map( A1 => data_in(22), A2 => n152, ZN => n5);
   U34 : OAI21_X1 port map( B1 => n37, B2 => n155, A => n2, ZN => n99);
   U35 : NAND2_X1 port map( A1 => n157, A2 => data_in(19), ZN => n2);
   U36 : OAI21_X1 port map( B1 => n123, B2 => n156, A => n26, ZN => n107);
   U37 : NAND2_X1 port map( A1 => data_in(11), A2 => n152, ZN => n26);
   U38 : OAI21_X1 port map( B1 => n42, B2 => n154, A => n7, ZN => n94);
   U39 : NAND2_X1 port map( A1 => data_in(24), A2 => n153, ZN => n7);
   U40 : OAI21_X1 port map( B1 => n39, B2 => n154, A => n4, ZN => n97);
   U41 : NAND2_X1 port map( A1 => data_in(21), A2 => n152, ZN => n4);
   U42 : OAI21_X1 port map( B1 => n121, B2 => n156, A => n28, ZN => n105);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n152, ZN => n28);
   U44 : OAI21_X1 port map( B1 => n124, B2 => n156, A => n25, ZN => n108);
   U45 : NAND2_X1 port map( A1 => data_in(10), A2 => n153, ZN => n25);
   U46 : OAI21_X1 port map( B1 => n36, B2 => n155, A => n33, ZN => n100);
   U47 : NAND2_X1 port map( A1 => data_in(18), A2 => n152, ZN => n33);
   U48 : OAI21_X1 port map( B1 => n127, B2 => n156, A => n22, ZN => n111);
   U49 : NAND2_X1 port map( A1 => data_in(7), A2 => n153, ZN => n22);
   U50 : OAI21_X1 port map( B1 => n38, B2 => n154, A => n3, ZN => n98);
   U51 : NAND2_X1 port map( A1 => data_in(20), A2 => n152, ZN => n3);
   U52 : OAI21_X1 port map( B1 => n35, B2 => n157, A => n32, ZN => n101);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n152, ZN => n32);
   U54 : OAI21_X1 port map( B1 => n128, B2 => n156, A => n21, ZN => n112);
   U55 : NAND2_X1 port map( A1 => data_in(6), A2 => n153, ZN => n21);
   U56 : OAI21_X1 port map( B1 => n122, B2 => n156, A => n27, ZN => n106);
   U57 : NAND2_X1 port map( A1 => data_in(12), A2 => n152, ZN => n27);
   U58 : OAI21_X1 port map( B1 => n125, B2 => n156, A => n24, ZN => n109);
   U59 : NAND2_X1 port map( A1 => data_in(9), A2 => n153, ZN => n24);
   U60 : OAI21_X1 port map( B1 => n34, B2 => n157, A => n31, ZN => n102);
   U61 : NAND2_X1 port map( A1 => data_in(16), A2 => n152, ZN => n31);
   U62 : OAI21_X1 port map( B1 => n126, B2 => n156, A => n23, ZN => n110);
   U63 : NAND2_X1 port map( A1 => data_in(8), A2 => n153, ZN => n23);
   U64 : OAI21_X1 port map( B1 => n129, B2 => n156, A => n20, ZN => n113);
   U65 : NAND2_X1 port map( A1 => data_in(5), A2 => n153, ZN => n20);
   U66 : OAI21_X1 port map( B1 => n131, B2 => n156, A => n18, ZN => n115);
   U67 : NAND2_X1 port map( A1 => data_in(3), A2 => n154, ZN => n18);
   U68 : OAI21_X1 port map( B1 => n130, B2 => n156, A => n19, ZN => n114);
   U69 : NAND2_X1 port map( A1 => data_in(4), A2 => n153, ZN => n19);
   U70 : OAI21_X1 port map( B1 => n133, B2 => n155, A => n16, ZN => n117);
   U71 : NAND2_X1 port map( A1 => data_in(1), A2 => n154, ZN => n16);
   U72 : OAI21_X1 port map( B1 => n132, B2 => n155, A => n17, ZN => n116);
   U73 : NAND2_X1 port map( A1 => data_in(2), A2 => n154, ZN => n17);
   U74 : OAI21_X1 port map( B1 => n134, B2 => n155, A => n15, ZN => n118);
   U75 : NAND2_X1 port map( A1 => data_in(0), A2 => n154, ZN => n15);
   U76 : OAI21_X1 port map( B1 => n49, B2 => n155, A => n14, ZN => n60);
   U77 : NAND2_X1 port map( A1 => data_in(27), A2 => n153, ZN => n10);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n154, ZN => n14);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_17 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_17;

architecture SYN_Behavioral of REG_NBIT32_17 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n216, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n216, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n216, Q => 
                           data_out(29), QN => n145);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n216, Q => 
                           data_out(26), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n216, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n216, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n217, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n216, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n217, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n217, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n217, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n217, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n216, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n217, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n217, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n217, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n216, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n218, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n218, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n218, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n218, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n218, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n218, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n218, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n217, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n217, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n217, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n218, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n217, Q => 
                           data_out(0), QN => n174);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n216, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n216, Q => 
                           data_out(27), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n216, Q => 
                           data_out(25), QN => n149);
   U2 : BUF_X1 port map( A => n207, Z => n215);
   U3 : BUF_X1 port map( A => n207, Z => n214);
   U4 : BUF_X1 port map( A => n215, Z => n209);
   U5 : BUF_X1 port map( A => n215, Z => n208);
   U6 : BUF_X1 port map( A => n215, Z => n210);
   U7 : BUF_X1 port map( A => n214, Z => n213);
   U8 : BUF_X1 port map( A => n214, Z => n212);
   U9 : BUF_X1 port map( A => n214, Z => n211);
   U10 : BUF_X1 port map( A => n219, Z => n216);
   U11 : BUF_X1 port map( A => n219, Z => n217);
   U12 : BUF_X1 port map( A => n219, Z => n218);
   U13 : INV_X1 port map( A => reset, ZN => n219);
   U14 : BUF_X1 port map( A => enable, Z => n207);
   U15 : OAI21_X1 port map( B1 => n147, B2 => n212, A => n29, ZN => n115);
   U16 : NAND2_X1 port map( A1 => data_in(27), A2 => n208, ZN => n29);
   U17 : OAI21_X1 port map( B1 => n173, B2 => n210, A => n3, ZN => n141);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n208, ZN => n3);
   U19 : OAI21_X1 port map( B1 => n172, B2 => n210, A => n4, ZN => n140);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n208, ZN => n4);
   U21 : OAI21_X1 port map( B1 => n171, B2 => n211, A => n5, ZN => n139);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n208, ZN => n5);
   U23 : OAI21_X1 port map( B1 => n170, B2 => n210, A => n6, ZN => n138);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n208, ZN => n6);
   U25 : OAI21_X1 port map( B1 => n169, B2 => n210, A => n7, ZN => n137);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n209, ZN => n7);
   U27 : OAI21_X1 port map( B1 => n168, B2 => n211, A => n8, ZN => n136);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n209, ZN => n8);
   U29 : OAI21_X1 port map( B1 => n167, B2 => n210, A => n9, ZN => n135);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n209, ZN => n9);
   U31 : OAI21_X1 port map( B1 => n166, B2 => n211, A => n10, ZN => n134);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n209, ZN => n10);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n211, A => n12, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(10), A2 => n209, ZN => n12);
   U35 : OAI21_X1 port map( B1 => n157, B2 => n212, A => n19, ZN => n125);
   U36 : NAND2_X1 port map( A1 => data_in(17), A2 => n209, ZN => n19);
   U37 : OAI21_X1 port map( B1 => n156, B2 => n212, A => n20, ZN => n124);
   U38 : NAND2_X1 port map( A1 => data_in(18), A2 => n209, ZN => n20);
   U39 : OAI21_X1 port map( B1 => n155, B2 => n212, A => n21, ZN => n123);
   U40 : NAND2_X1 port map( A1 => data_in(19), A2 => n209, ZN => n21);
   U41 : OAI21_X1 port map( B1 => n154, B2 => n212, A => n22, ZN => n122);
   U42 : NAND2_X1 port map( A1 => data_in(20), A2 => n209, ZN => n22);
   U43 : OAI21_X1 port map( B1 => n153, B2 => n212, A => n23, ZN => n121);
   U44 : NAND2_X1 port map( A1 => data_in(21), A2 => n209, ZN => n23);
   U45 : OAI21_X1 port map( B1 => n152, B2 => n212, A => n24, ZN => n120);
   U46 : NAND2_X1 port map( A1 => data_in(22), A2 => n209, ZN => n24);
   U47 : OAI21_X1 port map( B1 => n151, B2 => n212, A => n25, ZN => n119);
   U48 : NAND2_X1 port map( A1 => data_in(23), A2 => n209, ZN => n25);
   U49 : OAI21_X1 port map( B1 => n150, B2 => n212, A => n26, ZN => n118);
   U50 : NAND2_X1 port map( A1 => data_in(24), A2 => n208, ZN => n26);
   U51 : OAI21_X1 port map( B1 => n148, B2 => n212, A => n28, ZN => n116);
   U52 : NAND2_X1 port map( A1 => data_in(26), A2 => n208, ZN => n28);
   U53 : OAI21_X1 port map( B1 => n145, B2 => n213, A => n31, ZN => n113);
   U54 : NAND2_X1 port map( A1 => data_in(29), A2 => n208, ZN => n31);
   U55 : OAI21_X1 port map( B1 => n144, B2 => n213, A => n32, ZN => n112);
   U56 : NAND2_X1 port map( A1 => data_in(30), A2 => n208, ZN => n32);
   U57 : OAI21_X1 port map( B1 => n143, B2 => n211, A => n33, ZN => n111);
   U58 : NAND2_X1 port map( A1 => data_in(31), A2 => n208, ZN => n33);
   U59 : OAI21_X1 port map( B1 => n165, B2 => n211, A => n11, ZN => n133);
   U60 : NAND2_X1 port map( A1 => data_in(9), A2 => n210, ZN => n11);
   U61 : OAI21_X1 port map( B1 => n163, B2 => n211, A => n13, ZN => n131);
   U62 : NAND2_X1 port map( A1 => data_in(11), A2 => n210, ZN => n13);
   U63 : OAI21_X1 port map( B1 => n162, B2 => n211, A => n14, ZN => n130);
   U64 : NAND2_X1 port map( A1 => data_in(12), A2 => n210, ZN => n14);
   U65 : OAI21_X1 port map( B1 => n161, B2 => n211, A => n15, ZN => n129);
   U66 : NAND2_X1 port map( A1 => data_in(13), A2 => n210, ZN => n15);
   U67 : OAI21_X1 port map( B1 => n160, B2 => n211, A => n16, ZN => n128);
   U68 : NAND2_X1 port map( A1 => data_in(14), A2 => n210, ZN => n16);
   U69 : OAI21_X1 port map( B1 => n159, B2 => n211, A => n17, ZN => n127);
   U70 : NAND2_X1 port map( A1 => data_in(15), A2 => n210, ZN => n17);
   U71 : OAI21_X1 port map( B1 => n158, B2 => n212, A => n18, ZN => n126);
   U72 : NAND2_X1 port map( A1 => data_in(16), A2 => n210, ZN => n18);
   U73 : OAI21_X1 port map( B1 => n149, B2 => n212, A => n27, ZN => n117);
   U74 : NAND2_X1 port map( A1 => data_in(25), A2 => n208, ZN => n27);
   U75 : NAND2_X1 port map( A1 => data_in(28), A2 => n208, ZN => n30);
   U76 : OAI21_X1 port map( B1 => n174, B2 => n211, A => n2, ZN => n142);
   U77 : NAND2_X1 port map( A1 => n213, A2 => data_in(0), ZN => n2);
   U78 : OAI21_X1 port map( B1 => n146, B2 => n213, A => n30, ZN => n114);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_0 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_0;

architecture SYN_Behavioral of REG_NBIT32_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77
      , n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
      n92, n93, n94, n95, n97, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n96, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110 : std_logic;

begin
   
   reg_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n107, Q => 
                           data_out(30), QN => n64);
   reg_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n107, Q => 
                           data_out(29), QN => n63);
   reg_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n107, Q => 
                           data_out(28), QN => n62);
   reg_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n61);
   reg_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n60);
   reg_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n59);
   reg_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n58);
   reg_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n107, Q => 
                           data_out(23), QN => n57);
   reg_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n107, Q => 
                           data_out(22), QN => n56);
   reg_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n55);
   reg_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n54);
   reg_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n53);
   reg_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n52);
   reg_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n51);
   reg_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n50);
   reg_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n108, Q => 
                           data_out(15), QN => n48);
   reg_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n108, Q => 
                           data_out(14), QN => n47);
   reg_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n108, Q => 
                           data_out(13), QN => n46);
   reg_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n108, Q => 
                           data_out(12), QN => n45);
   reg_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n109, Q => 
                           data_out(11), QN => n44);
   reg_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n109, Q => 
                           data_out(10), QN => n43);
   reg_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n109, Q => 
                           data_out(9), QN => n42);
   reg_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n109, Q => 
                           data_out(8), QN => n41);
   reg_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n109, Q => 
                           data_out(7), QN => n40);
   reg_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n109, Q => 
                           data_out(6), QN => n39);
   reg_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n109, Q => 
                           data_out(5), QN => n38);
   reg_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n109, Q => 
                           data_out(4), QN => n37);
   reg_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n108, Q => 
                           data_out(3), QN => n36);
   reg_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n108, Q => 
                           data_out(2), QN => n35);
   reg_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n108, Q => 
                           data_out(1), QN => n34);
   reg_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n108, Q => 
                           data_out(0), QN => n33);
   reg_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n107, Q => 
                           data_out(31), QN => n96);
   U2 : BUF_X1 port map( A => n98, Z => n106);
   U3 : BUF_X1 port map( A => n98, Z => n105);
   U4 : BUF_X1 port map( A => n106, Z => n99);
   U5 : BUF_X1 port map( A => n106, Z => n100);
   U6 : BUF_X1 port map( A => n106, Z => n101);
   U7 : BUF_X1 port map( A => n105, Z => n104);
   U8 : BUF_X1 port map( A => n105, Z => n103);
   U9 : BUF_X1 port map( A => n105, Z => n102);
   U10 : BUF_X1 port map( A => n110, Z => n108);
   U11 : BUF_X1 port map( A => n110, Z => n107);
   U12 : BUF_X1 port map( A => n110, Z => n109);
   U13 : INV_X1 port map( A => reset, ZN => n110);
   U14 : BUF_X1 port map( A => enable, Z => n98);
   U15 : OAI21_X1 port map( B1 => n64, B2 => n101, A => n3, ZN => n95);
   U16 : NAND2_X1 port map( A1 => data_in(30), A2 => n99, ZN => n3);
   U17 : OAI21_X1 port map( B1 => n61, B2 => n101, A => n6, ZN => n92);
   U18 : OAI21_X1 port map( B1 => n63, B2 => n101, A => n4, ZN => n94);
   U19 : NAND2_X1 port map( A1 => data_in(29), A2 => n99, ZN => n4);
   U20 : OAI21_X1 port map( B1 => n60, B2 => n101, A => n7, ZN => n91);
   U21 : NAND2_X1 port map( A1 => data_in(26), A2 => n100, ZN => n7);
   U22 : OAI21_X1 port map( B1 => n48, B2 => n103, A => n18, ZN => n80);
   U23 : NAND2_X1 port map( A1 => data_in(15), A2 => n101, ZN => n18);
   U24 : OAI21_X1 port map( B1 => n57, B2 => n102, A => n10, ZN => n88);
   U25 : NAND2_X1 port map( A1 => data_in(23), A2 => n100, ZN => n10);
   U26 : OAI21_X1 port map( B1 => n62, B2 => n102, A => n5, ZN => n93);
   U27 : NAND2_X1 port map( A1 => data_in(28), A2 => n99, ZN => n5);
   U28 : OAI21_X1 port map( B1 => n59, B2 => n102, A => n8, ZN => n90);
   U29 : NAND2_X1 port map( A1 => data_in(25), A2 => n100, ZN => n8);
   U30 : OAI21_X1 port map( B1 => n47, B2 => n103, A => n19, ZN => n79);
   U31 : NAND2_X1 port map( A1 => data_in(14), A2 => n100, ZN => n19);
   U32 : OAI21_X1 port map( B1 => n56, B2 => n102, A => n11, ZN => n87);
   U33 : NAND2_X1 port map( A1 => data_in(22), A2 => n101, ZN => n11);
   U34 : OAI21_X1 port map( B1 => n44, B2 => n103, A => n22, ZN => n76);
   U35 : NAND2_X1 port map( A1 => data_in(11), A2 => n100, ZN => n22);
   U36 : OAI21_X1 port map( B1 => n53, B2 => n102, A => n14, ZN => n84);
   U37 : NAND2_X1 port map( A1 => data_in(19), A2 => n101, ZN => n14);
   U38 : OAI21_X1 port map( B1 => n58, B2 => n101, A => n9, ZN => n89);
   U39 : NAND2_X1 port map( A1 => data_in(24), A2 => n100, ZN => n9);
   U40 : OAI21_X1 port map( B1 => n55, B2 => n102, A => n12, ZN => n86);
   U41 : NAND2_X1 port map( A1 => data_in(21), A2 => n100, ZN => n12);
   U42 : OAI21_X1 port map( B1 => n46, B2 => n103, A => n20, ZN => n78);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n100, ZN => n20);
   U44 : OAI21_X1 port map( B1 => n43, B2 => n103, A => n23, ZN => n75);
   U45 : NAND2_X1 port map( A1 => data_in(10), A2 => n100, ZN => n23);
   U46 : OAI21_X1 port map( B1 => n52, B2 => n102, A => n15, ZN => n83);
   U47 : NAND2_X1 port map( A1 => data_in(18), A2 => n101, ZN => n15);
   U48 : OAI21_X1 port map( B1 => n40, B2 => n103, A => n26, ZN => n72);
   U49 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n26);
   U50 : OAI21_X1 port map( B1 => n54, B2 => n102, A => n13, ZN => n85);
   U51 : NAND2_X1 port map( A1 => data_in(20), A2 => n101, ZN => n13);
   U52 : OAI21_X1 port map( B1 => n51, B2 => n102, A => n16, ZN => n82);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n101, ZN => n16);
   U54 : OAI21_X1 port map( B1 => n39, B2 => n103, A => n27, ZN => n71);
   U55 : NAND2_X1 port map( A1 => data_in(6), A2 => n99, ZN => n27);
   U56 : OAI21_X1 port map( B1 => n45, B2 => n103, A => n21, ZN => n77);
   U57 : NAND2_X1 port map( A1 => data_in(12), A2 => n100, ZN => n21);
   U58 : OAI21_X1 port map( B1 => n42, B2 => n103, A => n24, ZN => n74);
   U59 : NAND2_X1 port map( A1 => data_in(9), A2 => n100, ZN => n24);
   U60 : OAI21_X1 port map( B1 => n50, B2 => n102, A => n17, ZN => n81);
   U61 : NAND2_X1 port map( A1 => data_in(16), A2 => n101, ZN => n17);
   U62 : OAI21_X1 port map( B1 => n41, B2 => n103, A => n25, ZN => n73);
   U63 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n25);
   U64 : OAI21_X1 port map( B1 => n38, B2 => n103, A => n28, ZN => n70);
   U65 : NAND2_X1 port map( A1 => data_in(5), A2 => n99, ZN => n28);
   U66 : OAI21_X1 port map( B1 => n36, B2 => n104, A => n30, ZN => n68);
   U67 : NAND2_X1 port map( A1 => data_in(3), A2 => n99, ZN => n30);
   U68 : OAI21_X1 port map( B1 => n37, B2 => n103, A => n29, ZN => n69);
   U69 : NAND2_X1 port map( A1 => data_in(4), A2 => n99, ZN => n29);
   U70 : OAI21_X1 port map( B1 => n34, B2 => n104, A => n32, ZN => n66);
   U71 : NAND2_X1 port map( A1 => data_in(1), A2 => n99, ZN => n32);
   U72 : OAI21_X1 port map( B1 => n35, B2 => n104, A => n31, ZN => n67);
   U73 : NAND2_X1 port map( A1 => data_in(2), A2 => n99, ZN => n31);
   U74 : OAI21_X1 port map( B1 => n33, B2 => n102, A => n49, ZN => n65);
   U75 : NAND2_X1 port map( A1 => data_in(0), A2 => n99, ZN => n49);
   U76 : OAI21_X1 port map( B1 => n96, B2 => n102, A => n2, ZN => n97);
   U77 : NAND2_X1 port map( A1 => data_in(27), A2 => n99, ZN => n6);
   U78 : NAND2_X1 port map( A1 => n104, A2 => data_in(31), ZN => n2);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector (31 
         downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out std_logic_vector (31 
         downto 0);  BMP : inout std_logic;  STALL : out std_logic_vector (1 
         downto 0);  ID_EN, RF_RD, SIGND, IMM_SEL, BPR_EN : in std_logic;  
         ALU_OPCODE : in std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, ALUB_SEL,
         UCB_EN, MEM_EN, MEM_DATA_SEL : in std_logic;  LD_SEL : in 
         std_logic_vector (2 downto 0);  ALR2_SEL : in std_logic;  CWB_SEL : in
         std_logic_vector (1 downto 0);  WB_SEL, RF_WR : in std_logic;  
         RF_MUX_SEL : in std_logic_vector (1 downto 0));

end Datapath;

architecture SYN_BEHAVIORAL of Datapath is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component RF_NBIT32_NREG32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component CWBU
      port( CLOCK : in std_logic;  ALU_OP : in std_logic_vector (0 to 4);  PSW 
            : in std_logic_vector (6 downto 0);  COND_SEL : out 
            std_logic_vector (1 downto 0);  CWB_SEL : in std_logic_vector (1 
            downto 0);  CWB_MUW_SEL : out std_logic_vector (1 downto 0));
   end component;
   
   component BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0
      port( clock, rst : in std_logic;  address : in std_logic_vector (31 
            downto 0);  d_in, w_en : in std_logic;  d_out : out std_logic);
   end component;
   
   component HDU_IR_SIZE32
      port( clk, rst : in std_logic;  IR : in std_logic_vector (31 downto 0);  
            STALL_CODE : out std_logic_vector (1 downto 0);  IF_STALL, ID_STALL
            , EX_STALL, MEM_STALL, WB_STALL : out std_logic);
   end component;
   
   component FWDU_IR_SIZE32
      port( CLOCK, RESET, EN : in std_logic;  IR : in std_logic_vector (31 
            downto 0);  FWD_A, FWD_B : out std_logic_vector (1 downto 0);  
            FWD_B2 : out std_logic;  ZDU_SEL : out std_logic_vector (1 downto 
            0));
   end component;
   
   component ALU_NBIT32
      port( CLOCK : in std_logic;  AluOpcode : in std_logic_vector (0 to 4);  A
            , B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            ALU_out : out std_logic_vector (31 downto 0);  Cout : out std_logic
            ;  COND : out std_logic_vector (5 downto 0));
   end component;
   
   component MUX3to1_NBIT5
      port( A, B, C : in std_logic_vector (4 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (4 downto 
            0));
   end component;
   
   component MUX2to1_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX4to1_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT2
      port( A, B, C, SEL : in std_logic_vector (1 downto 0);  Y : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component MUX2to1_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX5to1_NBIT32_0
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX2to1_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX3to1_NBIT32_1
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT32_2
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT32_3
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX2to1_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_8
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX3to1_NBIT32_0
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component PC_adder_1
      port( A, B : in std_logic_vector (31 downto 0);  Sum : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component PC_adder_0
      port( A, B : in std_logic_vector (31 downto 0);  Sum : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_4
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_5
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT7
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (6 downto 0);  data_out : out std_logic_vector (6 downto 0));
   end component;
   
   component REG_NBIT32_6
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_7
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_8
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_9
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_10
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component FFD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component REG_NBIT32_11
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_12
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component FFD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component REG_NBIT32_13
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_14
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_15
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_16
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_17
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_0
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IRAM_ADDR_31_port, IRAM_ADDR_30_port, 
      IRAM_ADDR_29_port, IRAM_ADDR_28_port, IRAM_ADDR_27_port, 
      IRAM_ADDR_26_port, IRAM_ADDR_25_port, IRAM_ADDR_24_port, 
      IRAM_ADDR_23_port, IRAM_ADDR_22_port, IRAM_ADDR_21_port, 
      IRAM_ADDR_20_port, IRAM_ADDR_19_port, IRAM_ADDR_18_port, 
      IRAM_ADDR_17_port, IRAM_ADDR_16_port, IRAM_ADDR_15_port, 
      IRAM_ADDR_14_port, IRAM_ADDR_13_port, IRAM_ADDR_12_port, 
      IRAM_ADDR_11_port, IRAM_ADDR_10_port, IRAM_ADDR_9_port, IRAM_ADDR_8_port,
      IRAM_ADDR_7_port, IRAM_ADDR_6_port, IRAM_ADDR_5_port, IRAM_ADDR_4_port, 
      IRAM_ADDR_3_port, IRAM_ADDR_2_port, IRAM_ADDR_1_port, IRAM_ADDR_0_port, 
      DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port, NPC_in_31_port, 
      NPC_in_30_port, NPC_in_29_port, NPC_in_28_port, NPC_in_27_port, 
      NPC_in_26_port, NPC_in_25_port, NPC_in_24_port, NPC_in_23_port, 
      NPC_in_22_port, NPC_in_21_port, NPC_in_20_port, NPC_in_19_port, 
      NPC_in_18_port, NPC_in_17_port, NPC_in_16_port, NPC_in_15_port, 
      NPC_in_14_port, NPC_in_13_port, NPC_in_12_port, NPC_in_11_port, 
      NPC_in_10_port, NPC_in_9_port, NPC_in_8_port, NPC_in_7_port, 
      NPC_in_6_port, NPC_in_5_port, NPC_in_4_port, NPC_in_3_port, NPC_in_2_port
      , NPC_in_1_port, NPC_in_0_port, PC_out_31_port, PC_out_30_port, 
      PC_out_29_port, PC_out_28_port, PC_out_27_port, PC_out_26_port, 
      PC_out_25_port, PC_out_24_port, PC_out_23_port, PC_out_22_port, 
      PC_out_21_port, PC_out_20_port, PC_out_19_port, PC_out_18_port, 
      PC_out_17_port, PC_out_16_port, PC_out_15_port, PC_out_14_port, 
      PC_out_13_port, PC_out_12_port, PC_out_11_port, PC_out_10_port, 
      PC_out_9_port, PC_out_8_port, PC_out_7_port, PC_out_6_port, PC_out_5_port
      , PC_out_4_port, PC_out_3_port, PC_out_2_port, PC_out_1_port, 
      PC_out_0_port, IR_out_31_port, IR_out_30_port, IR_out_29_port, 
      IR_out_28_port, IR_out_27_port, IR_out_26_port, IR_out_25_port, 
      IR_out_24_port, IR_out_23_port, IR_out_22_port, IR_out_21_port, 
      IR_out_20_port, IR_out_19_port, IR_out_18_port, IR_out_17_port, 
      IR_out_16_port, IR_out_15_port, IR_out_14_port, IR_out_13_port, 
      IR_out_12_port, IR_out_11_port, IR_out_10_port, IR_out_9_port, 
      IR_out_8_port, IR_out_7_port, IR_out_6_port, IR_out_5_port, IR_out_4_port
      , IR_out_3_port, IR_out_2_port, IR_out_1_port, IR_out_0_port, 
      NPC_out_31_port, NPC_out_30_port, NPC_out_29_port, NPC_out_28_port, 
      NPC_out_27_port, NPC_out_26_port, NPC_out_25_port, NPC_out_24_port, 
      NPC_out_23_port, NPC_out_22_port, NPC_out_21_port, NPC_out_20_port, 
      NPC_out_19_port, NPC_out_18_port, NPC_out_17_port, NPC_out_16_port, 
      NPC_out_15_port, NPC_out_14_port, NPC_out_13_port, NPC_out_12_port, 
      NPC_out_11_port, NPC_out_10_port, NPC_out_9_port, NPC_out_8_port, 
      NPC_out_7_port, NPC_out_6_port, NPC_out_5_port, NPC_out_4_port, 
      NPC_out_3_port, NPC_out_2_port, NPC_out_1_port, NPC_out_0_port, ID_ENABLE
      , PC2_out_31_port, PC2_out_30_port, PC2_out_29_port, PC2_out_28_port, 
      PC2_out_27_port, PC2_out_26_port, PC2_out_25_port, PC2_out_24_port, 
      PC2_out_23_port, PC2_out_22_port, PC2_out_21_port, PC2_out_20_port, 
      PC2_out_19_port, PC2_out_18_port, PC2_out_17_port, PC2_out_16_port, 
      PC2_out_15_port, PC2_out_14_port, PC2_out_13_port, PC2_out_12_port, 
      PC2_out_11_port, PC2_out_10_port, PC2_out_9_port, PC2_out_8_port, 
      PC2_out_7_port, PC2_out_6_port, PC2_out_5_port, PC2_out_4_port, 
      PC2_out_3_port, PC2_out_2_port, PC2_out_1_port, PC2_out_0_port, 
      RIMM_out_31_port, RIMM_out_30_port, RIMM_out_29_port, RIMM_out_28_port, 
      RIMM_out_27_port, RIMM_out_26_port, RIMM_out_25_port, RIMM_out_24_port, 
      RIMM_out_23_port, RIMM_out_22_port, RIMM_out_21_port, RIMM_out_20_port, 
      RIMM_out_19_port, RIMM_out_18_port, RIMM_out_17_port, RIMM_out_16_port, 
      RIMM_out_15_port, RIMM_out_14_port, RIMM_out_13_port, RIMM_out_12_port, 
      RIMM_out_11_port, RIMM_out_10_port, RIMM_out_9_port, RIMM_out_8_port, 
      RIMM_out_7_port, RIMM_out_6_port, RIMM_out_5_port, RIMM_out_4_port, 
      RIMM_out_3_port, RIMM_out_2_port, RIMM_out_1_port, RIMM_out_0_port, 
      RWB1_out_31_port, RWB1_out_30_port, RWB1_out_29_port, RWB1_out_28_port, 
      RWB1_out_27_port, RWB1_out_26_port, RWB1_out_25_port, RWB1_out_24_port, 
      RWB1_out_23_port, RWB1_out_22_port, RWB1_out_21_port, RWB1_out_20_port, 
      RWB1_out_19_port, RWB1_out_18_port, RWB1_out_17_port, RWB1_out_16_port, 
      RWB1_out_15_port, RWB1_out_14_port, RWB1_out_13_port, RWB1_out_12_port, 
      RWB1_out_11_port, RWB1_out_10_port, RWB1_out_9_port, RWB1_out_8_port, 
      RWB1_out_7_port, RWB1_out_6_port, RWB1_out_5_port, RWB1_out_4_port, 
      RWB1_out_3_port, RWB1_out_2_port, RWB1_out_1_port, RWB1_out_0_port, 
      BHT_out, PRD_OUT, NPC2_out_31_port, NPC2_out_30_port, NPC2_out_29_port, 
      NPC2_out_28_port, NPC2_out_27_port, NPC2_out_26_port, NPC2_out_25_port, 
      NPC2_out_24_port, NPC2_out_23_port, NPC2_out_22_port, NPC2_out_21_port, 
      NPC2_out_20_port, NPC2_out_19_port, NPC2_out_18_port, NPC2_out_17_port, 
      NPC2_out_16_port, NPC2_out_15_port, NPC2_out_14_port, NPC2_out_13_port, 
      NPC2_out_12_port, NPC2_out_11_port, NPC2_out_10_port, NPC2_out_9_port, 
      NPC2_out_8_port, NPC2_out_7_port, NPC2_out_6_port, NPC2_out_5_port, 
      NPC2_out_4_port, NPC2_out_3_port, NPC2_out_2_port, NPC2_out_1_port, 
      NPC2_out_0_port, JADDER_out_31_port, JADDER_out_30_port, 
      JADDER_out_29_port, JADDER_out_28_port, JADDER_out_27_port, 
      JADDER_out_26_port, JADDER_out_25_port, JADDER_out_24_port, 
      JADDER_out_23_port, JADDER_out_22_port, JADDER_out_21_port, 
      JADDER_out_20_port, JADDER_out_19_port, JADDER_out_18_port, 
      JADDER_out_17_port, JADDER_out_16_port, JADDER_out_15_port, 
      JADDER_out_14_port, JADDER_out_13_port, JADDER_out_12_port, 
      JADDER_out_11_port, JADDER_out_10_port, JADDER_out_9_port, 
      JADDER_out_8_port, JADDER_out_7_port, JADDER_out_6_port, 
      JADDER_out_5_port, JADDER_out_4_port, JADDER_out_3_port, 
      JADDER_out_2_port, JADDER_out_1_port, JADDER_out_0_port, 
      JADDER2_out_31_port, JADDER2_out_30_port, JADDER2_out_29_port, 
      JADDER2_out_28_port, JADDER2_out_27_port, JADDER2_out_26_port, 
      JADDER2_out_25_port, JADDER2_out_24_port, JADDER2_out_23_port, 
      JADDER2_out_22_port, JADDER2_out_21_port, JADDER2_out_20_port, 
      JADDER2_out_19_port, JADDER2_out_18_port, JADDER2_out_17_port, 
      JADDER2_out_16_port, JADDER2_out_15_port, JADDER2_out_14_port, 
      JADDER2_out_13_port, JADDER2_out_12_port, JADDER2_out_11_port, 
      JADDER2_out_10_port, JADDER2_out_9_port, JADDER2_out_8_port, 
      JADDER2_out_7_port, JADDER2_out_6_port, JADDER2_out_5_port, 
      JADDER2_out_4_port, JADDER2_out_3_port, JADDER2_out_2_port, 
      JADDER2_out_1_port, JADDER2_out_0_port, BPR_EN2, EX_ENABLE, 
      PC3_out_31_port, PC3_out_30_port, PC3_out_29_port, PC3_out_28_port, 
      PC3_out_27_port, PC3_out_26_port, PC3_out_25_port, PC3_out_24_port, 
      PC3_out_23_port, PC3_out_22_port, PC3_out_21_port, PC3_out_20_port, 
      PC3_out_19_port, PC3_out_18_port, PC3_out_17_port, PC3_out_16_port, 
      PC3_out_15_port, PC3_out_14_port, PC3_out_13_port, PC3_out_12_port, 
      PC3_out_11_port, PC3_out_10_port, PC3_out_9_port, PC3_out_8_port, 
      PC3_out_7_port, PC3_out_6_port, PC3_out_5_port, PC3_out_4_port, 
      PC3_out_3_port, PC3_out_2_port, PC3_out_1_port, PC3_out_0_port, 
      RWB2_out_31_port, RWB2_out_30_port, RWB2_out_29_port, RWB2_out_28_port, 
      RWB2_out_27_port, RWB2_out_26_port, RWB2_out_25_port, RWB2_out_24_port, 
      RWB2_out_23_port, RWB2_out_22_port, RWB2_out_21_port, RWB2_out_20_port, 
      RWB2_out_19_port, RWB2_out_18_port, RWB2_out_17_port, RWB2_out_16_port, 
      RWB2_out_15_port, RWB2_out_14_port, RWB2_out_13_port, RWB2_out_12_port, 
      RWB2_out_11_port, RWB2_out_10_port, RWB2_out_9_port, RWB2_out_8_port, 
      RWB2_out_7_port, RWB2_out_6_port, RWB2_out_5_port, RWB2_out_4_port, 
      RWB2_out_3_port, RWB2_out_2_port, RWB2_out_1_port, RWB2_out_0_port, 
      RB_out_31_port, RB_out_30_port, RB_out_29_port, RB_out_28_port, 
      RB_out_27_port, RB_out_26_port, RB_out_25_port, RB_out_24_port, 
      RB_out_23_port, RB_out_22_port, RB_out_21_port, RB_out_20_port, 
      RB_out_19_port, RB_out_18_port, RB_out_17_port, RB_out_16_port, 
      RB_out_15_port, RB_out_14_port, RB_out_13_port, RB_out_12_port, 
      RB_out_11_port, RB_out_10_port, RB_out_9_port, RB_out_8_port, 
      RB_out_7_port, RB_out_6_port, RB_out_5_port, RB_out_4_port, RB_out_3_port
      , RB_out_2_port, RB_out_1_port, RB_out_0_port, B2_out_31_port, 
      B2_out_30_port, B2_out_29_port, B2_out_28_port, B2_out_27_port, 
      B2_out_26_port, B2_out_25_port, B2_out_24_port, B2_out_23_port, 
      B2_out_22_port, B2_out_21_port, B2_out_20_port, B2_out_19_port, 
      B2_out_18_port, B2_out_17_port, B2_out_16_port, B2_out_15_port, 
      B2_out_14_port, B2_out_13_port, B2_out_12_port, B2_out_11_port, 
      B2_out_10_port, B2_out_9_port, B2_out_8_port, B2_out_7_port, 
      B2_out_6_port, B2_out_5_port, B2_out_4_port, B2_out_3_port, B2_out_2_port
      , B2_out_1_port, B2_out_0_port, ALR_in_31_port, ALR_in_30_port, 
      ALR_in_29_port, ALR_in_28_port, ALR_in_27_port, ALR_in_26_port, 
      ALR_in_25_port, ALR_in_24_port, ALR_in_23_port, ALR_in_22_port, 
      ALR_in_21_port, ALR_in_20_port, ALR_in_19_port, ALR_in_18_port, 
      ALR_in_17_port, ALR_in_16_port, ALR_in_15_port, ALR_in_14_port, 
      ALR_in_13_port, ALR_in_12_port, ALR_in_11_port, ALR_in_10_port, 
      ALR_in_9_port, ALR_in_8_port, ALR_in_7_port, ALR_in_6_port, ALR_in_5_port
      , ALR_in_4_port, ALR_in_3_port, ALR_in_2_port, ALR_in_1_port, 
      ALR_in_0_port, NPC3_out_31_port, NPC3_out_30_port, NPC3_out_29_port, 
      NPC3_out_28_port, NPC3_out_27_port, NPC3_out_26_port, NPC3_out_25_port, 
      NPC3_out_24_port, NPC3_out_23_port, NPC3_out_22_port, NPC3_out_21_port, 
      NPC3_out_20_port, NPC3_out_19_port, NPC3_out_18_port, NPC3_out_17_port, 
      NPC3_out_16_port, NPC3_out_15_port, NPC3_out_14_port, NPC3_out_13_port, 
      NPC3_out_12_port, NPC3_out_11_port, NPC3_out_10_port, NPC3_out_9_port, 
      NPC3_out_8_port, NPC3_out_7_port, NPC3_out_6_port, NPC3_out_5_port, 
      NPC3_out_4_port, NPC3_out_3_port, NPC3_out_2_port, NPC3_out_1_port, 
      NPC3_out_0_port, PSW_in_6_port, PSW_in_5_port, PSW_in_4_port, 
      PSW_in_3_port, PSW_in_2_port, PSW_in_1_port, PSW_in_0_port, 
      PSW_out_6_port, PSW_out_5_port, PSW_out_4_port, PSW_out_3_port, 
      PSW_out_2_port, PSW_out_1_port, PSW_out_0_port, MEM_ENABLE, 
      ALR2_in_31_port, ALR2_in_30_port, ALR2_in_29_port, ALR2_in_28_port, 
      ALR2_in_27_port, ALR2_in_26_port, ALR2_in_25_port, ALR2_in_24_port, 
      ALR2_in_23_port, ALR2_in_22_port, ALR2_in_21_port, ALR2_in_20_port, 
      ALR2_in_19_port, ALR2_in_18_port, ALR2_in_17_port, ALR2_in_16_port, 
      ALR2_in_15_port, ALR2_in_14_port, ALR2_in_13_port, ALR2_in_12_port, 
      ALR2_in_11_port, ALR2_in_10_port, ALR2_in_9_port, ALR2_in_8_port, 
      ALR2_in_7_port, ALR2_in_6_port, ALR2_in_5_port, ALR2_in_4_port, 
      ALR2_in_3_port, ALR2_in_2_port, ALR2_in_1_port, ALR2_in_0_port, 
      ALR2_out_31_port, ALR2_out_30_port, ALR2_out_29_port, ALR2_out_28_port, 
      ALR2_out_27_port, ALR2_out_26_port, ALR2_out_25_port, ALR2_out_24_port, 
      ALR2_out_23_port, ALR2_out_22_port, ALR2_out_21_port, ALR2_out_20_port, 
      ALR2_out_19_port, ALR2_out_18_port, ALR2_out_17_port, ALR2_out_16_port, 
      ALR2_out_15_port, ALR2_out_14_port, ALR2_out_13_port, ALR2_out_12_port, 
      ALR2_out_11_port, ALR2_out_10_port, ALR2_out_9_port, ALR2_out_8_port, 
      ALR2_out_7_port, ALR2_out_6_port, ALR2_out_5_port, ALR2_out_4_port, 
      ALR2_out_3_port, ALR2_out_2_port, ALR2_out_1_port, ALR2_out_0_port, 
      RWB3_out_20_port, RWB3_out_19_port, RWB3_out_18_port, RWB3_out_17_port, 
      RWB3_out_16_port, RWB3_out_15_port, RWB3_out_14_port, RWB3_out_13_port, 
      RWB3_out_12_port, RWB3_out_11_port, IMM_out_31_port, IMM_out_30_port, 
      IMM_out_29_port, IMM_out_28_port, IMM_out_27_port, IMM_out_26_port, 
      IMM_out_25_port, IMM_out_24_port, IMM_out_23_port, IMM_out_22_port, 
      IMM_out_21_port, IMM_out_20_port, IMM_out_19_port, IMM_out_18_port, 
      IMM_out_17_port, IMM_out_16_port, IMM_out_15_port, IMM_out_14_port, 
      IMM_out_13_port, IMM_out_12_port, IMM_out_11_port, IMM_out_10_port, 
      IMM_out_9_port, IMM_out_8_port, IMM_out_7_port, IMM_out_6_port, 
      IMM_out_5_port, IMM_out_4_port, IMM_out_3_port, IMM_out_2_port, 
      IMM_out_1_port, IMM_out_0_port, PC_SEL_1_port, PC_MUX_out_31_port, 
      PC_MUX_out_30_port, PC_MUX_out_29_port, PC_MUX_out_28_port, 
      PC_MUX_out_27_port, PC_MUX_out_26_port, PC_MUX_out_25_port, 
      PC_MUX_out_24_port, PC_MUX_out_23_port, PC_MUX_out_22_port, 
      PC_MUX_out_21_port, PC_MUX_out_20_port, PC_MUX_out_19_port, 
      PC_MUX_out_18_port, PC_MUX_out_17_port, PC_MUX_out_16_port, 
      PC_MUX_out_15_port, PC_MUX_out_14_port, PC_MUX_out_13_port, 
      PC_MUX_out_12_port, PC_MUX_out_11_port, PC_MUX_out_10_port, 
      PC_MUX_out_9_port, PC_MUX_out_8_port, PC_MUX_out_7_port, 
      PC_MUX_out_6_port, PC_MUX_out_5_port, PC_MUX_out_4_port, 
      PC_MUX_out_3_port, PC_MUX_out_2_port, PC_MUX_out_1_port, 
      PC_MUX_out_0_port, IRAMMUX_SEL, BHT_in_31_port, BHT_in_30_port, 
      BHT_in_29_port, BHT_in_28_port, BHT_in_27_port, BHT_in_26_port, 
      BHT_in_25_port, BHT_in_24_port, BHT_in_23_port, BHT_in_22_port, 
      BHT_in_21_port, BHT_in_20_port, BHT_in_19_port, BHT_in_18_port, 
      BHT_in_17_port, BHT_in_16_port, BHT_in_15_port, BHT_in_14_port, 
      BHT_in_13_port, BHT_in_12_port, BHT_in_11_port, BHT_in_10_port, 
      BHT_in_9_port, BHT_in_8_port, BHT_in_7_port, BHT_in_6_port, BHT_in_5_port
      , BHT_in_4_port, BHT_in_3_port, BHT_in_2_port, BHT_in_1_port, 
      BHT_in_0_port, FWDA_OUT_31_port, FWDA_OUT_30_port, FWDA_OUT_29_port, 
      FWDA_OUT_28_port, FWDA_OUT_27_port, FWDA_OUT_26_port, FWDA_OUT_25_port, 
      FWDA_OUT_24_port, FWDA_OUT_23_port, FWDA_OUT_22_port, FWDA_OUT_21_port, 
      FWDA_OUT_20_port, FWDA_OUT_19_port, FWDA_OUT_18_port, FWDA_OUT_17_port, 
      FWDA_OUT_16_port, FWDA_OUT_15_port, FWDA_OUT_14_port, FWDA_OUT_13_port, 
      FWDA_OUT_12_port, FWDA_OUT_11_port, FWDA_OUT_10_port, FWDA_OUT_9_port, 
      FWDA_OUT_8_port, FWDA_OUT_7_port, FWDA_OUT_6_port, FWDA_OUT_5_port, 
      FWDA_OUT_4_port, FWDA_OUT_3_port, FWDA_OUT_2_port, FWDA_OUT_1_port, 
      FWDA_OUT_0_port, A_in_31_port, A_in_30_port, A_in_29_port, A_in_28_port, 
      A_in_27_port, A_in_26_port, A_in_25_port, A_in_24_port, A_in_23_port, 
      A_in_22_port, A_in_21_port, A_in_20_port, A_in_19_port, A_in_18_port, 
      A_in_17_port, A_in_16_port, A_in_15_port, A_in_14_port, A_in_13_port, 
      A_in_12_port, A_in_11_port, A_in_10_port, A_in_9_port, A_in_8_port, 
      A_in_7_port, A_in_6_port, A_in_5_port, A_in_4_port, A_in_3_port, 
      A_in_2_port, A_in_1_port, A_in_0_port, FWDB_OUT_31_port, FWDB_OUT_30_port
      , FWDB_OUT_29_port, FWDB_OUT_28_port, FWDB_OUT_27_port, FWDB_OUT_26_port,
      FWDB_OUT_25_port, FWDB_OUT_24_port, FWDB_OUT_23_port, FWDB_OUT_22_port, 
      FWDB_OUT_21_port, FWDB_OUT_20_port, FWDB_OUT_19_port, FWDB_OUT_18_port, 
      FWDB_OUT_17_port, FWDB_OUT_16_port, FWDB_OUT_15_port, FWDB_OUT_14_port, 
      FWDB_OUT_13_port, FWDB_OUT_12_port, FWDB_OUT_11_port, FWDB_OUT_10_port, 
      FWDB_OUT_9_port, FWDB_OUT_8_port, FWDB_OUT_7_port, FWDB_OUT_6_port, 
      FWDB_OUT_5_port, FWDB_OUT_4_port, FWDB_OUT_3_port, FWDB_OUT_2_port, 
      FWDB_OUT_1_port, FWDB_OUT_0_port, B_in_31_port, B_in_30_port, 
      B_in_29_port, B_in_28_port, B_in_27_port, B_in_26_port, B_in_25_port, 
      B_in_24_port, B_in_23_port, B_in_22_port, B_in_21_port, B_in_20_port, 
      B_in_19_port, B_in_18_port, B_in_17_port, B_in_16_port, B_in_15_port, 
      B_in_14_port, B_in_13_port, B_in_12_port, B_in_11_port, B_in_10_port, 
      B_in_9_port, B_in_8_port, B_in_7_port, B_in_6_port, B_in_5_port, 
      B_in_4_port, B_in_3_port, B_in_2_port, B_in_1_port, B_in_0_port, 
      RA_out_31_port, RA_out_30_port, RA_out_29_port, RA_out_28_port, 
      RA_out_27_port, RA_out_26_port, RA_out_25_port, RA_out_24_port, 
      RA_out_23_port, RA_out_22_port, RA_out_21_port, RA_out_20_port, 
      RA_out_19_port, RA_out_18_port, RA_out_17_port, RA_out_16_port, 
      RA_out_15_port, RA_out_14_port, RA_out_13_port, RA_out_12_port, 
      RA_out_11_port, RA_out_10_port, RA_out_9_port, RA_out_8_port, 
      RA_out_7_port, RA_out_6_port, RA_out_5_port, RA_out_4_port, RA_out_3_port
      , RA_out_2_port, RA_out_1_port, RA_out_0_port, WB_in_31_port, 
      WB_in_30_port, WB_in_29_port, WB_in_28_port, WB_in_27_port, WB_in_26_port
      , WB_in_25_port, WB_in_24_port, WB_in_23_port, WB_in_22_port, 
      WB_in_21_port, WB_in_20_port, WB_in_19_port, WB_in_18_port, WB_in_17_port
      , WB_in_16_port, WB_in_15_port, WB_in_14_port, WB_in_13_port, 
      WB_in_12_port, WB_in_11_port, WB_in_10_port, WB_in_9_port, WB_in_8_port, 
      WB_in_7_port, WB_in_6_port, WB_in_5_port, WB_in_4_port, WB_in_3_port, 
      WB_in_2_port, WB_in_1_port, WB_in_0_port, FWDA_SEL_1_port, 
      FWDA_SEL_0_port, FWDB_SEL_1_port, FWDB_SEL_0_port, CWB_MUX2_out_31_port, 
      CWB_MUX2_out_30_port, CWB_MUX2_out_29_port, CWB_MUX2_out_28_port, 
      CWB_MUX2_out_27_port, CWB_MUX2_out_26_port, CWB_MUX2_out_25_port, 
      CWB_MUX2_out_24_port, CWB_MUX2_out_23_port, CWB_MUX2_out_22_port, 
      CWB_MUX2_out_21_port, CWB_MUX2_out_20_port, CWB_MUX2_out_19_port, 
      CWB_MUX2_out_18_port, CWB_MUX2_out_17_port, CWB_MUX2_out_16_port, 
      CWB_MUX2_out_15_port, CWB_MUX2_out_14_port, CWB_MUX2_out_13_port, 
      CWB_MUX2_out_12_port, CWB_MUX2_out_11_port, CWB_MUX2_out_10_port, 
      CWB_MUX2_out_9_port, CWB_MUX2_out_8_port, CWB_MUX2_out_7_port, 
      CWB_MUX2_out_6_port, CWB_MUX2_out_5_port, CWB_MUX2_out_4_port, 
      CWB_MUX2_out_3_port, CWB_MUX2_out_2_port, CWB_MUX2_out_1_port, 
      CWB_MUX2_out_0_port, ZDU_SEL_1_port, ZDU_SEL_0_port, ZDU_MUX_out_30_port,
      ZDU_MUX_out_29_port, ZDU_MUX_out_28_port, ZDU_MUX_out_27_port, 
      ZDU_MUX_out_26_port, ZDU_MUX_out_25_port, ZDU_MUX_out_24_port, 
      ZDU_MUX_out_23_port, ZDU_MUX_out_22_port, ZDU_MUX_out_21_port, 
      ZDU_MUX_out_20_port, ZDU_MUX_out_19_port, ZDU_MUX_out_18_port, 
      ZDU_MUX_out_17_port, ZDU_MUX_out_16_port, ZDU_MUX_out_15_port, 
      ZDU_MUX_out_14_port, ZDU_MUX_out_13_port, ZDU_MUX_out_12_port, 
      ZDU_MUX_out_11_port, ZDU_MUX_out_10_port, ZDU_MUX_out_9_port, 
      ZDU_MUX_out_8_port, ZDU_MUX_out_7_port, ZDU_MUX_out_6_port, 
      ZDU_MUX_out_5_port, ZDU_MUX_out_4_port, ZDU_MUX_out_3_port, 
      ZDU_MUX_out_2_port, ZDU_MUX_out_1_port, ZDU_MUX_out_0_port, 
      B2_MUX_out_31_port, B2_MUX_out_30_port, B2_MUX_out_29_port, 
      B2_MUX_out_28_port, B2_MUX_out_27_port, B2_MUX_out_26_port, 
      B2_MUX_out_25_port, B2_MUX_out_24_port, B2_MUX_out_23_port, 
      B2_MUX_out_22_port, B2_MUX_out_21_port, B2_MUX_out_20_port, 
      B2_MUX_out_19_port, B2_MUX_out_18_port, B2_MUX_out_17_port, 
      B2_MUX_out_16_port, B2_MUX_out_15_port, B2_MUX_out_14_port, 
      B2_MUX_out_13_port, B2_MUX_out_12_port, B2_MUX_out_11_port, 
      B2_MUX_out_10_port, B2_MUX_out_9_port, B2_MUX_out_8_port, 
      B2_MUX_out_7_port, B2_MUX_out_6_port, B2_MUX_out_5_port, 
      B2_MUX_out_4_port, B2_MUX_out_3_port, B2_MUX_out_2_port, 
      B2_MUX_out_1_port, B2_MUX_out_0_port, LMD_out_31_port, LMD_out_30_port, 
      LMD_out_29_port, LMD_out_28_port, LMD_out_27_port, LMD_out_26_port, 
      LMD_out_25_port, LMD_out_24_port, LMD_out_23_port, LMD_out_22_port, 
      LMD_out_21_port, LMD_out_20_port, LMD_out_19_port, LMD_out_18_port, 
      LMD_out_17_port, LMD_out_16_port, LMD_out_15_port, LMD_out_14_port, 
      LMD_out_13_port, LMD_out_12_port, LMD_out_11_port, LMD_out_10_port, 
      LMD_out_9_port, LMD_out_8_port, LMD_out_7_port, LMD_out_6_port, 
      LMD_out_5_port, LMD_out_4_port, LMD_out_3_port, LMD_out_2_port, 
      LMD_out_1_port, LMD_out_0_port, CWB_out_1_port, CWB_out_0_port, 
      CWB_MUX_SEL_1_port, CWB_MUX_SEL_0_port, CWB2_SEL_1_port, CWB2_SEL_0_port,
      FWDB2_SEL, RF_MUX_out_4_port, RF_MUX_out_3_port, RF_MUX_out_2_port, 
      RF_MUX_out_1_port, RF_MUX_out_0_port, IF_STALL, EX_STALL, MEM_STALL, 
      RF_RD_en, N14, n3, n7, n8, n9, n10, n11, n12, n13, n14_port, n15, n16, 
      n17, n18, n19, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n_1586, n_1587, n_1588, n_1589,
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610 : std_logic;

begin
   IRAM_ADDR <= ( IRAM_ADDR_31_port, IRAM_ADDR_30_port, IRAM_ADDR_29_port, 
      IRAM_ADDR_28_port, IRAM_ADDR_27_port, IRAM_ADDR_26_port, 
      IRAM_ADDR_25_port, IRAM_ADDR_24_port, IRAM_ADDR_23_port, 
      IRAM_ADDR_22_port, IRAM_ADDR_21_port, IRAM_ADDR_20_port, 
      IRAM_ADDR_19_port, IRAM_ADDR_18_port, IRAM_ADDR_17_port, 
      IRAM_ADDR_16_port, IRAM_ADDR_15_port, IRAM_ADDR_14_port, 
      IRAM_ADDR_13_port, IRAM_ADDR_12_port, IRAM_ADDR_11_port, 
      IRAM_ADDR_10_port, IRAM_ADDR_9_port, IRAM_ADDR_8_port, IRAM_ADDR_7_port, 
      IRAM_ADDR_6_port, IRAM_ADDR_5_port, IRAM_ADDR_4_port, IRAM_ADDR_3_port, 
      IRAM_ADDR_2_port, IRAM_ADDR_1_port, IRAM_ADDR_0_port );
   DATA_ADDR <= ( DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U28 : XOR2_X1 port map( A => PRD_OUT, B => n19, Z => n3);
   RegPC : REG_NBIT32_0 port map( clk => CLK, reset => n50, enable => n38, 
                           data_in(31) => NPC_in_31_port, data_in(30) => 
                           NPC_in_30_port, data_in(29) => NPC_in_29_port, 
                           data_in(28) => NPC_in_28_port, data_in(27) => 
                           NPC_in_27_port, data_in(26) => NPC_in_26_port, 
                           data_in(25) => NPC_in_25_port, data_in(24) => 
                           NPC_in_24_port, data_in(23) => NPC_in_23_port, 
                           data_in(22) => NPC_in_22_port, data_in(21) => 
                           NPC_in_21_port, data_in(20) => NPC_in_20_port, 
                           data_in(19) => NPC_in_19_port, data_in(18) => 
                           NPC_in_18_port, data_in(17) => NPC_in_17_port, 
                           data_in(16) => NPC_in_16_port, data_in(15) => 
                           NPC_in_15_port, data_in(14) => NPC_in_14_port, 
                           data_in(13) => NPC_in_13_port, data_in(12) => 
                           NPC_in_12_port, data_in(11) => NPC_in_11_port, 
                           data_in(10) => NPC_in_10_port, data_in(9) => 
                           NPC_in_9_port, data_in(8) => NPC_in_8_port, 
                           data_in(7) => NPC_in_7_port, data_in(6) => 
                           NPC_in_6_port, data_in(5) => NPC_in_5_port, 
                           data_in(4) => NPC_in_4_port, data_in(3) => 
                           NPC_in_3_port, data_in(2) => NPC_in_2_port, 
                           data_in(1) => NPC_in_1_port, data_in(0) => 
                           NPC_in_0_port, data_out(31) => PC_out_31_port, 
                           data_out(30) => PC_out_30_port, data_out(29) => 
                           PC_out_29_port, data_out(28) => PC_out_28_port, 
                           data_out(27) => PC_out_27_port, data_out(26) => 
                           PC_out_26_port, data_out(25) => PC_out_25_port, 
                           data_out(24) => PC_out_24_port, data_out(23) => 
                           PC_out_23_port, data_out(22) => PC_out_22_port, 
                           data_out(21) => PC_out_21_port, data_out(20) => 
                           PC_out_20_port, data_out(19) => PC_out_19_port, 
                           data_out(18) => PC_out_18_port, data_out(17) => 
                           PC_out_17_port, data_out(16) => PC_out_16_port, 
                           data_out(15) => PC_out_15_port, data_out(14) => 
                           PC_out_14_port, data_out(13) => PC_out_13_port, 
                           data_out(12) => PC_out_12_port, data_out(11) => 
                           PC_out_11_port, data_out(10) => PC_out_10_port, 
                           data_out(9) => PC_out_9_port, data_out(8) => 
                           PC_out_8_port, data_out(7) => PC_out_7_port, 
                           data_out(6) => PC_out_6_port, data_out(5) => 
                           PC_out_5_port, data_out(4) => PC_out_4_port, 
                           data_out(3) => PC_out_3_port, data_out(2) => 
                           PC_out_2_port, data_out(1) => PC_out_1_port, 
                           data_out(0) => PC_out_0_port);
   RegIR : REG_NBIT32_17 port map( clk => CLK, reset => n50, enable => n38, 
                           data_in(31) => IRAM_OUT(31), data_in(30) => 
                           IRAM_OUT(30), data_in(29) => IRAM_OUT(29), 
                           data_in(28) => IRAM_OUT(28), data_in(27) => 
                           IRAM_OUT(27), data_in(26) => IRAM_OUT(26), 
                           data_in(25) => IRAM_OUT(25), data_in(24) => 
                           IRAM_OUT(24), data_in(23) => IRAM_OUT(23), 
                           data_in(22) => IRAM_OUT(22), data_in(21) => 
                           IRAM_OUT(21), data_in(20) => IRAM_OUT(20), 
                           data_in(19) => IRAM_OUT(19), data_in(18) => 
                           IRAM_OUT(18), data_in(17) => IRAM_OUT(17), 
                           data_in(16) => IRAM_OUT(16), data_in(15) => 
                           IRAM_OUT(15), data_in(14) => IRAM_OUT(14), 
                           data_in(13) => IRAM_OUT(13), data_in(12) => 
                           IRAM_OUT(12), data_in(11) => IRAM_OUT(11), 
                           data_in(10) => IRAM_OUT(10), data_in(9) => 
                           IRAM_OUT(9), data_in(8) => IRAM_OUT(8), data_in(7) 
                           => IRAM_OUT(7), data_in(6) => IRAM_OUT(6), 
                           data_in(5) => IRAM_OUT(5), data_in(4) => IRAM_OUT(4)
                           , data_in(3) => IRAM_OUT(3), data_in(2) => 
                           IRAM_OUT(2), data_in(1) => IRAM_OUT(1), data_in(0) 
                           => IRAM_OUT(0), data_out(31) => IR_out_31_port, 
                           data_out(30) => IR_out_30_port, data_out(29) => 
                           IR_out_29_port, data_out(28) => IR_out_28_port, 
                           data_out(27) => IR_out_27_port, data_out(26) => 
                           IR_out_26_port, data_out(25) => IR_out_25_port, 
                           data_out(24) => IR_out_24_port, data_out(23) => 
                           IR_out_23_port, data_out(22) => IR_out_22_port, 
                           data_out(21) => IR_out_21_port, data_out(20) => 
                           IR_out_20_port, data_out(19) => IR_out_19_port, 
                           data_out(18) => IR_out_18_port, data_out(17) => 
                           IR_out_17_port, data_out(16) => IR_out_16_port, 
                           data_out(15) => IR_out_15_port, data_out(14) => 
                           IR_out_14_port, data_out(13) => IR_out_13_port, 
                           data_out(12) => IR_out_12_port, data_out(11) => 
                           IR_out_11_port, data_out(10) => IR_out_10_port, 
                           data_out(9) => IR_out_9_port, data_out(8) => 
                           IR_out_8_port, data_out(7) => IR_out_7_port, 
                           data_out(6) => IR_out_6_port, data_out(5) => 
                           IR_out_5_port, data_out(4) => IR_out_4_port, 
                           data_out(3) => IR_out_3_port, data_out(2) => 
                           IR_out_2_port, data_out(1) => IR_out_1_port, 
                           data_out(0) => IR_out_0_port);
   RegNPC : REG_NBIT32_16 port map( clk => CLK, reset => n50, enable => n38, 
                           data_in(31) => NPC_in_31_port, data_in(30) => 
                           NPC_in_30_port, data_in(29) => NPC_in_29_port, 
                           data_in(28) => NPC_in_28_port, data_in(27) => 
                           NPC_in_27_port, data_in(26) => NPC_in_26_port, 
                           data_in(25) => NPC_in_25_port, data_in(24) => 
                           NPC_in_24_port, data_in(23) => NPC_in_23_port, 
                           data_in(22) => NPC_in_22_port, data_in(21) => 
                           NPC_in_21_port, data_in(20) => NPC_in_20_port, 
                           data_in(19) => NPC_in_19_port, data_in(18) => 
                           NPC_in_18_port, data_in(17) => NPC_in_17_port, 
                           data_in(16) => NPC_in_16_port, data_in(15) => 
                           NPC_in_15_port, data_in(14) => NPC_in_14_port, 
                           data_in(13) => NPC_in_13_port, data_in(12) => 
                           NPC_in_12_port, data_in(11) => NPC_in_11_port, 
                           data_in(10) => NPC_in_10_port, data_in(9) => 
                           NPC_in_9_port, data_in(8) => NPC_in_8_port, 
                           data_in(7) => NPC_in_7_port, data_in(6) => 
                           NPC_in_6_port, data_in(5) => NPC_in_5_port, 
                           data_in(4) => NPC_in_4_port, data_in(3) => 
                           NPC_in_3_port, data_in(2) => NPC_in_2_port, 
                           data_in(1) => NPC_in_1_port, data_in(0) => 
                           NPC_in_0_port, data_out(31) => NPC_out_31_port, 
                           data_out(30) => NPC_out_30_port, data_out(29) => 
                           NPC_out_29_port, data_out(28) => NPC_out_28_port, 
                           data_out(27) => NPC_out_27_port, data_out(26) => 
                           NPC_out_26_port, data_out(25) => NPC_out_25_port, 
                           data_out(24) => NPC_out_24_port, data_out(23) => 
                           NPC_out_23_port, data_out(22) => NPC_out_22_port, 
                           data_out(21) => NPC_out_21_port, data_out(20) => 
                           NPC_out_20_port, data_out(19) => NPC_out_19_port, 
                           data_out(18) => NPC_out_18_port, data_out(17) => 
                           NPC_out_17_port, data_out(16) => NPC_out_16_port, 
                           data_out(15) => NPC_out_15_port, data_out(14) => 
                           NPC_out_14_port, data_out(13) => NPC_out_13_port, 
                           data_out(12) => NPC_out_12_port, data_out(11) => 
                           NPC_out_11_port, data_out(10) => NPC_out_10_port, 
                           data_out(9) => NPC_out_9_port, data_out(8) => 
                           NPC_out_8_port, data_out(7) => NPC_out_7_port, 
                           data_out(6) => NPC_out_6_port, data_out(5) => 
                           NPC_out_5_port, data_out(4) => NPC_out_4_port, 
                           data_out(3) => NPC_out_3_port, data_out(2) => 
                           NPC_out_2_port, data_out(1) => NPC_out_1_port, 
                           data_out(0) => NPC_out_0_port);
   RegPC2 : REG_NBIT32_15 port map( clk => CLK, reset => n50, enable => n41, 
                           data_in(31) => PC_out_31_port, data_in(30) => 
                           PC_out_30_port, data_in(29) => PC_out_29_port, 
                           data_in(28) => PC_out_28_port, data_in(27) => 
                           PC_out_27_port, data_in(26) => PC_out_26_port, 
                           data_in(25) => PC_out_25_port, data_in(24) => 
                           PC_out_24_port, data_in(23) => PC_out_23_port, 
                           data_in(22) => PC_out_22_port, data_in(21) => 
                           PC_out_21_port, data_in(20) => PC_out_20_port, 
                           data_in(19) => PC_out_19_port, data_in(18) => 
                           PC_out_18_port, data_in(17) => PC_out_17_port, 
                           data_in(16) => PC_out_16_port, data_in(15) => 
                           PC_out_15_port, data_in(14) => PC_out_14_port, 
                           data_in(13) => PC_out_13_port, data_in(12) => 
                           PC_out_12_port, data_in(11) => PC_out_11_port, 
                           data_in(10) => PC_out_10_port, data_in(9) => 
                           PC_out_9_port, data_in(8) => PC_out_8_port, 
                           data_in(7) => PC_out_7_port, data_in(6) => 
                           PC_out_6_port, data_in(5) => PC_out_5_port, 
                           data_in(4) => PC_out_4_port, data_in(3) => 
                           PC_out_3_port, data_in(2) => PC_out_2_port, 
                           data_in(1) => PC_out_1_port, data_in(0) => 
                           PC_out_0_port, data_out(31) => PC2_out_31_port, 
                           data_out(30) => PC2_out_30_port, data_out(29) => 
                           PC2_out_29_port, data_out(28) => PC2_out_28_port, 
                           data_out(27) => PC2_out_27_port, data_out(26) => 
                           PC2_out_26_port, data_out(25) => PC2_out_25_port, 
                           data_out(24) => PC2_out_24_port, data_out(23) => 
                           PC2_out_23_port, data_out(22) => PC2_out_22_port, 
                           data_out(21) => PC2_out_21_port, data_out(20) => 
                           PC2_out_20_port, data_out(19) => PC2_out_19_port, 
                           data_out(18) => PC2_out_18_port, data_out(17) => 
                           PC2_out_17_port, data_out(16) => PC2_out_16_port, 
                           data_out(15) => PC2_out_15_port, data_out(14) => 
                           PC2_out_14_port, data_out(13) => PC2_out_13_port, 
                           data_out(12) => PC2_out_12_port, data_out(11) => 
                           PC2_out_11_port, data_out(10) => PC2_out_10_port, 
                           data_out(9) => PC2_out_9_port, data_out(8) => 
                           PC2_out_8_port, data_out(7) => PC2_out_7_port, 
                           data_out(6) => PC2_out_6_port, data_out(5) => 
                           PC2_out_5_port, data_out(4) => PC2_out_4_port, 
                           data_out(3) => PC2_out_3_port, data_out(2) => 
                           PC2_out_2_port, data_out(1) => PC2_out_1_port, 
                           data_out(0) => PC2_out_0_port);
   RegIMM : REG_NBIT32_14 port map( clk => CLK, reset => n50, enable => n41, 
                           data_in(31) => N14, data_in(30) => N14, data_in(29) 
                           => N14, data_in(28) => N14, data_in(27) => N14, 
                           data_in(26) => N14, data_in(25) => N14, data_in(24) 
                           => N14, data_in(23) => N14, data_in(22) => N14, 
                           data_in(21) => N14, data_in(20) => N14, data_in(19) 
                           => N14, data_in(18) => N14, data_in(17) => N14, 
                           data_in(16) => N14, data_in(15) => IR_out_15_port, 
                           data_in(14) => IR_out_14_port, data_in(13) => 
                           IR_out_13_port, data_in(12) => IR_out_12_port, 
                           data_in(11) => IR_out_11_port, data_in(10) => 
                           IR_out_10_port, data_in(9) => IR_out_9_port, 
                           data_in(8) => IR_out_8_port, data_in(7) => 
                           IR_out_7_port, data_in(6) => IR_out_6_port, 
                           data_in(5) => IR_out_5_port, data_in(4) => 
                           IR_out_4_port, data_in(3) => IR_out_3_port, 
                           data_in(2) => IR_out_2_port, data_in(1) => 
                           IR_out_1_port, data_in(0) => IR_out_0_port, 
                           data_out(31) => RIMM_out_31_port, data_out(30) => 
                           RIMM_out_30_port, data_out(29) => RIMM_out_29_port, 
                           data_out(28) => RIMM_out_28_port, data_out(27) => 
                           RIMM_out_27_port, data_out(26) => RIMM_out_26_port, 
                           data_out(25) => RIMM_out_25_port, data_out(24) => 
                           RIMM_out_24_port, data_out(23) => RIMM_out_23_port, 
                           data_out(22) => RIMM_out_22_port, data_out(21) => 
                           RIMM_out_21_port, data_out(20) => RIMM_out_20_port, 
                           data_out(19) => RIMM_out_19_port, data_out(18) => 
                           RIMM_out_18_port, data_out(17) => RIMM_out_17_port, 
                           data_out(16) => RIMM_out_16_port, data_out(15) => 
                           RIMM_out_15_port, data_out(14) => RIMM_out_14_port, 
                           data_out(13) => RIMM_out_13_port, data_out(12) => 
                           RIMM_out_12_port, data_out(11) => RIMM_out_11_port, 
                           data_out(10) => RIMM_out_10_port, data_out(9) => 
                           RIMM_out_9_port, data_out(8) => RIMM_out_8_port, 
                           data_out(7) => RIMM_out_7_port, data_out(6) => 
                           RIMM_out_6_port, data_out(5) => RIMM_out_5_port, 
                           data_out(4) => RIMM_out_4_port, data_out(3) => 
                           RIMM_out_3_port, data_out(2) => RIMM_out_2_port, 
                           data_out(1) => RIMM_out_1_port, data_out(0) => 
                           RIMM_out_0_port);
   RegWB1 : REG_NBIT32_13 port map( clk => CLK, reset => n50, enable => n41, 
                           data_in(31) => IR_out_31_port, data_in(30) => 
                           IR_out_30_port, data_in(29) => IR_out_29_port, 
                           data_in(28) => IR_out_28_port, data_in(27) => 
                           IR_out_27_port, data_in(26) => IR_out_26_port, 
                           data_in(25) => IR_out_25_port, data_in(24) => 
                           IR_out_24_port, data_in(23) => IR_out_23_port, 
                           data_in(22) => IR_out_22_port, data_in(21) => 
                           IR_out_21_port, data_in(20) => IR_out_20_port, 
                           data_in(19) => IR_out_19_port, data_in(18) => n36, 
                           data_in(17) => IR_out_17_port, data_in(16) => 
                           IR_out_16_port, data_in(15) => IR_out_15_port, 
                           data_in(14) => IR_out_14_port, data_in(13) => 
                           IR_out_13_port, data_in(12) => IR_out_12_port, 
                           data_in(11) => IR_out_11_port, data_in(10) => 
                           IR_out_10_port, data_in(9) => IR_out_9_port, 
                           data_in(8) => IR_out_8_port, data_in(7) => 
                           IR_out_7_port, data_in(6) => IR_out_6_port, 
                           data_in(5) => IR_out_5_port, data_in(4) => 
                           IR_out_4_port, data_in(3) => IR_out_3_port, 
                           data_in(2) => IR_out_2_port, data_in(1) => 
                           IR_out_1_port, data_in(0) => IR_out_0_port, 
                           data_out(31) => RWB1_out_31_port, data_out(30) => 
                           RWB1_out_30_port, data_out(29) => RWB1_out_29_port, 
                           data_out(28) => RWB1_out_28_port, data_out(27) => 
                           RWB1_out_27_port, data_out(26) => RWB1_out_26_port, 
                           data_out(25) => RWB1_out_25_port, data_out(24) => 
                           RWB1_out_24_port, data_out(23) => RWB1_out_23_port, 
                           data_out(22) => RWB1_out_22_port, data_out(21) => 
                           RWB1_out_21_port, data_out(20) => RWB1_out_20_port, 
                           data_out(19) => RWB1_out_19_port, data_out(18) => 
                           RWB1_out_18_port, data_out(17) => RWB1_out_17_port, 
                           data_out(16) => RWB1_out_16_port, data_out(15) => 
                           RWB1_out_15_port, data_out(14) => RWB1_out_14_port, 
                           data_out(13) => RWB1_out_13_port, data_out(12) => 
                           RWB1_out_12_port, data_out(11) => RWB1_out_11_port, 
                           data_out(10) => RWB1_out_10_port, data_out(9) => 
                           RWB1_out_9_port, data_out(8) => RWB1_out_8_port, 
                           data_out(7) => RWB1_out_7_port, data_out(6) => 
                           RWB1_out_6_port, data_out(5) => RWB1_out_5_port, 
                           data_out(4) => RWB1_out_4_port, data_out(3) => 
                           RWB1_out_3_port, data_out(2) => RWB1_out_2_port, 
                           data_out(1) => RWB1_out_1_port, data_out(0) => 
                           RWB1_out_0_port);
   F_PRD : FFD_0 port map( D => BHT_out, CK => CLK, RESET => n50, ENABLE => n41
                           , Q => PRD_OUT);
   RegNPC2 : REG_NBIT32_12 port map( clk => CLK, reset => n50, enable => n41, 
                           data_in(31) => NPC_out_31_port, data_in(30) => 
                           NPC_out_30_port, data_in(29) => NPC_out_29_port, 
                           data_in(28) => NPC_out_28_port, data_in(27) => 
                           NPC_out_27_port, data_in(26) => NPC_out_26_port, 
                           data_in(25) => NPC_out_25_port, data_in(24) => 
                           NPC_out_24_port, data_in(23) => NPC_out_23_port, 
                           data_in(22) => NPC_out_22_port, data_in(21) => 
                           NPC_out_21_port, data_in(20) => NPC_out_20_port, 
                           data_in(19) => NPC_out_19_port, data_in(18) => 
                           NPC_out_18_port, data_in(17) => NPC_out_17_port, 
                           data_in(16) => NPC_out_16_port, data_in(15) => 
                           NPC_out_15_port, data_in(14) => NPC_out_14_port, 
                           data_in(13) => NPC_out_13_port, data_in(12) => 
                           NPC_out_12_port, data_in(11) => NPC_out_11_port, 
                           data_in(10) => NPC_out_10_port, data_in(9) => 
                           NPC_out_9_port, data_in(8) => NPC_out_8_port, 
                           data_in(7) => NPC_out_7_port, data_in(6) => 
                           NPC_out_6_port, data_in(5) => NPC_out_5_port, 
                           data_in(4) => NPC_out_4_port, data_in(3) => 
                           NPC_out_3_port, data_in(2) => NPC_out_2_port, 
                           data_in(1) => NPC_out_1_port, data_in(0) => 
                           NPC_out_0_port, data_out(31) => NPC2_out_31_port, 
                           data_out(30) => NPC2_out_30_port, data_out(29) => 
                           NPC2_out_29_port, data_out(28) => NPC2_out_28_port, 
                           data_out(27) => NPC2_out_27_port, data_out(26) => 
                           NPC2_out_26_port, data_out(25) => NPC2_out_25_port, 
                           data_out(24) => NPC2_out_24_port, data_out(23) => 
                           NPC2_out_23_port, data_out(22) => NPC2_out_22_port, 
                           data_out(21) => NPC2_out_21_port, data_out(20) => 
                           NPC2_out_20_port, data_out(19) => NPC2_out_19_port, 
                           data_out(18) => NPC2_out_18_port, data_out(17) => 
                           NPC2_out_17_port, data_out(16) => NPC2_out_16_port, 
                           data_out(15) => NPC2_out_15_port, data_out(14) => 
                           NPC2_out_14_port, data_out(13) => NPC2_out_13_port, 
                           data_out(12) => NPC2_out_12_port, data_out(11) => 
                           NPC2_out_11_port, data_out(10) => NPC2_out_10_port, 
                           data_out(9) => NPC2_out_9_port, data_out(8) => 
                           NPC2_out_8_port, data_out(7) => NPC2_out_7_port, 
                           data_out(6) => NPC2_out_6_port, data_out(5) => 
                           NPC2_out_5_port, data_out(4) => NPC2_out_4_port, 
                           data_out(3) => NPC2_out_3_port, data_out(2) => 
                           NPC2_out_2_port, data_out(1) => NPC2_out_1_port, 
                           data_out(0) => NPC2_out_0_port);
   RegJADD2 : REG_NBIT32_11 port map( clk => CLK, reset => n50, enable => n41, 
                           data_in(31) => JADDER_out_31_port, data_in(30) => 
                           JADDER_out_30_port, data_in(29) => 
                           JADDER_out_29_port, data_in(28) => 
                           JADDER_out_28_port, data_in(27) => 
                           JADDER_out_27_port, data_in(26) => 
                           JADDER_out_26_port, data_in(25) => 
                           JADDER_out_25_port, data_in(24) => 
                           JADDER_out_24_port, data_in(23) => 
                           JADDER_out_23_port, data_in(22) => 
                           JADDER_out_22_port, data_in(21) => 
                           JADDER_out_21_port, data_in(20) => 
                           JADDER_out_20_port, data_in(19) => 
                           JADDER_out_19_port, data_in(18) => 
                           JADDER_out_18_port, data_in(17) => 
                           JADDER_out_17_port, data_in(16) => 
                           JADDER_out_16_port, data_in(15) => 
                           JADDER_out_15_port, data_in(14) => 
                           JADDER_out_14_port, data_in(13) => 
                           JADDER_out_13_port, data_in(12) => 
                           JADDER_out_12_port, data_in(11) => 
                           JADDER_out_11_port, data_in(10) => 
                           JADDER_out_10_port, data_in(9) => JADDER_out_9_port,
                           data_in(8) => JADDER_out_8_port, data_in(7) => 
                           JADDER_out_7_port, data_in(6) => JADDER_out_6_port, 
                           data_in(5) => JADDER_out_5_port, data_in(4) => 
                           JADDER_out_4_port, data_in(3) => JADDER_out_3_port, 
                           data_in(2) => JADDER_out_2_port, data_in(1) => 
                           JADDER_out_1_port, data_in(0) => JADDER_out_0_port, 
                           data_out(31) => JADDER2_out_31_port, data_out(30) =>
                           JADDER2_out_30_port, data_out(29) => 
                           JADDER2_out_29_port, data_out(28) => 
                           JADDER2_out_28_port, data_out(27) => 
                           JADDER2_out_27_port, data_out(26) => 
                           JADDER2_out_26_port, data_out(25) => 
                           JADDER2_out_25_port, data_out(24) => 
                           JADDER2_out_24_port, data_out(23) => 
                           JADDER2_out_23_port, data_out(22) => 
                           JADDER2_out_22_port, data_out(21) => 
                           JADDER2_out_21_port, data_out(20) => 
                           JADDER2_out_20_port, data_out(19) => 
                           JADDER2_out_19_port, data_out(18) => 
                           JADDER2_out_18_port, data_out(17) => 
                           JADDER2_out_17_port, data_out(16) => 
                           JADDER2_out_16_port, data_out(15) => 
                           JADDER2_out_15_port, data_out(14) => 
                           JADDER2_out_14_port, data_out(13) => 
                           JADDER2_out_13_port, data_out(12) => 
                           JADDER2_out_12_port, data_out(11) => 
                           JADDER2_out_11_port, data_out(10) => 
                           JADDER2_out_10_port, data_out(9) => 
                           JADDER2_out_9_port, data_out(8) => 
                           JADDER2_out_8_port, data_out(7) => 
                           JADDER2_out_7_port, data_out(6) => 
                           JADDER2_out_6_port, data_out(5) => 
                           JADDER2_out_5_port, data_out(4) => 
                           JADDER2_out_4_port, data_out(3) => 
                           JADDER2_out_3_port, data_out(2) => 
                           JADDER2_out_2_port, data_out(1) => 
                           JADDER2_out_1_port, data_out(0) => 
                           JADDER2_out_0_port);
   F_JR : FFD_1 port map( D => BPR_EN, CK => CLK, RESET => n50, ENABLE => n41, 
                           Q => BPR_EN2);
   RegPC3 : REG_NBIT32_10 port map( clk => CLK, reset => n50, enable => n40, 
                           data_in(31) => PC2_out_31_port, data_in(30) => 
                           PC2_out_30_port, data_in(29) => PC2_out_29_port, 
                           data_in(28) => PC2_out_28_port, data_in(27) => 
                           PC2_out_27_port, data_in(26) => PC2_out_26_port, 
                           data_in(25) => PC2_out_25_port, data_in(24) => 
                           PC2_out_24_port, data_in(23) => PC2_out_23_port, 
                           data_in(22) => PC2_out_22_port, data_in(21) => 
                           PC2_out_21_port, data_in(20) => PC2_out_20_port, 
                           data_in(19) => PC2_out_19_port, data_in(18) => 
                           PC2_out_18_port, data_in(17) => PC2_out_17_port, 
                           data_in(16) => PC2_out_16_port, data_in(15) => 
                           PC2_out_15_port, data_in(14) => PC2_out_14_port, 
                           data_in(13) => PC2_out_13_port, data_in(12) => 
                           PC2_out_12_port, data_in(11) => PC2_out_11_port, 
                           data_in(10) => PC2_out_10_port, data_in(9) => 
                           PC2_out_9_port, data_in(8) => PC2_out_8_port, 
                           data_in(7) => PC2_out_7_port, data_in(6) => 
                           PC2_out_6_port, data_in(5) => PC2_out_5_port, 
                           data_in(4) => PC2_out_4_port, data_in(3) => 
                           PC2_out_3_port, data_in(2) => PC2_out_2_port, 
                           data_in(1) => PC2_out_1_port, data_in(0) => 
                           PC2_out_0_port, data_out(31) => PC3_out_31_port, 
                           data_out(30) => PC3_out_30_port, data_out(29) => 
                           PC3_out_29_port, data_out(28) => PC3_out_28_port, 
                           data_out(27) => PC3_out_27_port, data_out(26) => 
                           PC3_out_26_port, data_out(25) => PC3_out_25_port, 
                           data_out(24) => PC3_out_24_port, data_out(23) => 
                           PC3_out_23_port, data_out(22) => PC3_out_22_port, 
                           data_out(21) => PC3_out_21_port, data_out(20) => 
                           PC3_out_20_port, data_out(19) => PC3_out_19_port, 
                           data_out(18) => PC3_out_18_port, data_out(17) => 
                           PC3_out_17_port, data_out(16) => PC3_out_16_port, 
                           data_out(15) => PC3_out_15_port, data_out(14) => 
                           PC3_out_14_port, data_out(13) => PC3_out_13_port, 
                           data_out(12) => PC3_out_12_port, data_out(11) => 
                           PC3_out_11_port, data_out(10) => PC3_out_10_port, 
                           data_out(9) => PC3_out_9_port, data_out(8) => 
                           PC3_out_8_port, data_out(7) => PC3_out_7_port, 
                           data_out(6) => PC3_out_6_port, data_out(5) => 
                           PC3_out_5_port, data_out(4) => PC3_out_4_port, 
                           data_out(3) => PC3_out_3_port, data_out(2) => 
                           PC3_out_2_port, data_out(1) => PC3_out_1_port, 
                           data_out(0) => PC3_out_0_port);
   RegWB2 : REG_NBIT32_9 port map( clk => CLK, reset => n51, enable => n40, 
                           data_in(31) => RWB1_out_31_port, data_in(30) => 
                           RWB1_out_30_port, data_in(29) => RWB1_out_29_port, 
                           data_in(28) => RWB1_out_28_port, data_in(27) => 
                           RWB1_out_27_port, data_in(26) => RWB1_out_26_port, 
                           data_in(25) => RWB1_out_25_port, data_in(24) => 
                           RWB1_out_24_port, data_in(23) => RWB1_out_23_port, 
                           data_in(22) => RWB1_out_22_port, data_in(21) => 
                           RWB1_out_21_port, data_in(20) => RWB1_out_20_port, 
                           data_in(19) => RWB1_out_19_port, data_in(18) => 
                           RWB1_out_18_port, data_in(17) => RWB1_out_17_port, 
                           data_in(16) => RWB1_out_16_port, data_in(15) => 
                           RWB1_out_15_port, data_in(14) => RWB1_out_14_port, 
                           data_in(13) => RWB1_out_13_port, data_in(12) => 
                           RWB1_out_12_port, data_in(11) => RWB1_out_11_port, 
                           data_in(10) => RWB1_out_10_port, data_in(9) => 
                           RWB1_out_9_port, data_in(8) => RWB1_out_8_port, 
                           data_in(7) => RWB1_out_7_port, data_in(6) => 
                           RWB1_out_6_port, data_in(5) => RWB1_out_5_port, 
                           data_in(4) => RWB1_out_4_port, data_in(3) => 
                           RWB1_out_3_port, data_in(2) => RWB1_out_2_port, 
                           data_in(1) => RWB1_out_1_port, data_in(0) => 
                           RWB1_out_0_port, data_out(31) => RWB2_out_31_port, 
                           data_out(30) => RWB2_out_30_port, data_out(29) => 
                           RWB2_out_29_port, data_out(28) => RWB2_out_28_port, 
                           data_out(27) => RWB2_out_27_port, data_out(26) => 
                           RWB2_out_26_port, data_out(25) => RWB2_out_25_port, 
                           data_out(24) => RWB2_out_24_port, data_out(23) => 
                           RWB2_out_23_port, data_out(22) => RWB2_out_22_port, 
                           data_out(21) => RWB2_out_21_port, data_out(20) => 
                           RWB2_out_20_port, data_out(19) => RWB2_out_19_port, 
                           data_out(18) => RWB2_out_18_port, data_out(17) => 
                           RWB2_out_17_port, data_out(16) => RWB2_out_16_port, 
                           data_out(15) => RWB2_out_15_port, data_out(14) => 
                           RWB2_out_14_port, data_out(13) => RWB2_out_13_port, 
                           data_out(12) => RWB2_out_12_port, data_out(11) => 
                           RWB2_out_11_port, data_out(10) => RWB2_out_10_port, 
                           data_out(9) => RWB2_out_9_port, data_out(8) => 
                           RWB2_out_8_port, data_out(7) => RWB2_out_7_port, 
                           data_out(6) => RWB2_out_6_port, data_out(5) => 
                           RWB2_out_5_port, data_out(4) => RWB2_out_4_port, 
                           data_out(3) => RWB2_out_3_port, data_out(2) => 
                           RWB2_out_2_port, data_out(1) => RWB2_out_1_port, 
                           data_out(0) => RWB2_out_0_port);
   RegB2 : REG_NBIT32_8 port map( clk => CLK, reset => n51, enable => n40, 
                           data_in(31) => RB_out_31_port, data_in(30) => 
                           RB_out_30_port, data_in(29) => RB_out_29_port, 
                           data_in(28) => RB_out_28_port, data_in(27) => 
                           RB_out_27_port, data_in(26) => RB_out_26_port, 
                           data_in(25) => RB_out_25_port, data_in(24) => 
                           RB_out_24_port, data_in(23) => RB_out_23_port, 
                           data_in(22) => RB_out_22_port, data_in(21) => 
                           RB_out_21_port, data_in(20) => RB_out_20_port, 
                           data_in(19) => RB_out_19_port, data_in(18) => 
                           RB_out_18_port, data_in(17) => RB_out_17_port, 
                           data_in(16) => RB_out_16_port, data_in(15) => 
                           RB_out_15_port, data_in(14) => RB_out_14_port, 
                           data_in(13) => RB_out_13_port, data_in(12) => 
                           RB_out_12_port, data_in(11) => RB_out_11_port, 
                           data_in(10) => RB_out_10_port, data_in(9) => 
                           RB_out_9_port, data_in(8) => RB_out_8_port, 
                           data_in(7) => RB_out_7_port, data_in(6) => 
                           RB_out_6_port, data_in(5) => RB_out_5_port, 
                           data_in(4) => RB_out_4_port, data_in(3) => 
                           RB_out_3_port, data_in(2) => RB_out_2_port, 
                           data_in(1) => RB_out_1_port, data_in(0) => 
                           RB_out_0_port, data_out(31) => B2_out_31_port, 
                           data_out(30) => B2_out_30_port, data_out(29) => 
                           B2_out_29_port, data_out(28) => B2_out_28_port, 
                           data_out(27) => B2_out_27_port, data_out(26) => 
                           B2_out_26_port, data_out(25) => B2_out_25_port, 
                           data_out(24) => B2_out_24_port, data_out(23) => 
                           B2_out_23_port, data_out(22) => B2_out_22_port, 
                           data_out(21) => B2_out_21_port, data_out(20) => 
                           B2_out_20_port, data_out(19) => B2_out_19_port, 
                           data_out(18) => B2_out_18_port, data_out(17) => 
                           B2_out_17_port, data_out(16) => B2_out_16_port, 
                           data_out(15) => B2_out_15_port, data_out(14) => 
                           B2_out_14_port, data_out(13) => B2_out_13_port, 
                           data_out(12) => B2_out_12_port, data_out(11) => 
                           B2_out_11_port, data_out(10) => B2_out_10_port, 
                           data_out(9) => B2_out_9_port, data_out(8) => 
                           B2_out_8_port, data_out(7) => B2_out_7_port, 
                           data_out(6) => B2_out_6_port, data_out(5) => 
                           B2_out_5_port, data_out(4) => B2_out_4_port, 
                           data_out(3) => B2_out_3_port, data_out(2) => 
                           B2_out_2_port, data_out(1) => B2_out_1_port, 
                           data_out(0) => B2_out_0_port);
   RegALR : REG_NBIT32_7 port map( clk => CLK, reset => n51, enable => n40, 
                           data_in(31) => ALR_in_31_port, data_in(30) => 
                           ALR_in_30_port, data_in(29) => ALR_in_29_port, 
                           data_in(28) => ALR_in_28_port, data_in(27) => 
                           ALR_in_27_port, data_in(26) => ALR_in_26_port, 
                           data_in(25) => ALR_in_25_port, data_in(24) => 
                           ALR_in_24_port, data_in(23) => ALR_in_23_port, 
                           data_in(22) => ALR_in_22_port, data_in(21) => 
                           ALR_in_21_port, data_in(20) => ALR_in_20_port, 
                           data_in(19) => ALR_in_19_port, data_in(18) => 
                           ALR_in_18_port, data_in(17) => ALR_in_17_port, 
                           data_in(16) => ALR_in_16_port, data_in(15) => 
                           ALR_in_15_port, data_in(14) => ALR_in_14_port, 
                           data_in(13) => ALR_in_13_port, data_in(12) => 
                           ALR_in_12_port, data_in(11) => ALR_in_11_port, 
                           data_in(10) => ALR_in_10_port, data_in(9) => 
                           ALR_in_9_port, data_in(8) => ALR_in_8_port, 
                           data_in(7) => ALR_in_7_port, data_in(6) => 
                           ALR_in_6_port, data_in(5) => ALR_in_5_port, 
                           data_in(4) => ALR_in_4_port, data_in(3) => 
                           ALR_in_3_port, data_in(2) => ALR_in_2_port, 
                           data_in(1) => ALR_in_1_port, data_in(0) => 
                           ALR_in_0_port, data_out(31) => DATA_ADDR_31_port, 
                           data_out(30) => DATA_ADDR_30_port, data_out(29) => 
                           DATA_ADDR_29_port, data_out(28) => DATA_ADDR_28_port
                           , data_out(27) => DATA_ADDR_27_port, data_out(26) =>
                           DATA_ADDR_26_port, data_out(25) => DATA_ADDR_25_port
                           , data_out(24) => DATA_ADDR_24_port, data_out(23) =>
                           DATA_ADDR_23_port, data_out(22) => DATA_ADDR_22_port
                           , data_out(21) => DATA_ADDR_21_port, data_out(20) =>
                           DATA_ADDR_20_port, data_out(19) => DATA_ADDR_19_port
                           , data_out(18) => DATA_ADDR_18_port, data_out(17) =>
                           DATA_ADDR_17_port, data_out(16) => DATA_ADDR_16_port
                           , data_out(15) => DATA_ADDR_15_port, data_out(14) =>
                           DATA_ADDR_14_port, data_out(13) => DATA_ADDR_13_port
                           , data_out(12) => DATA_ADDR_12_port, data_out(11) =>
                           DATA_ADDR_11_port, data_out(10) => DATA_ADDR_10_port
                           , data_out(9) => DATA_ADDR_9_port, data_out(8) => 
                           DATA_ADDR_8_port, data_out(7) => DATA_ADDR_7_port, 
                           data_out(6) => DATA_ADDR_6_port, data_out(5) => 
                           DATA_ADDR_5_port, data_out(4) => DATA_ADDR_4_port, 
                           data_out(3) => DATA_ADDR_3_port, data_out(2) => 
                           DATA_ADDR_2_port, data_out(1) => DATA_ADDR_1_port, 
                           data_out(0) => DATA_ADDR_0_port);
   RegNPC3 : REG_NBIT32_6 port map( clk => CLK, reset => n50, enable => n40, 
                           data_in(31) => NPC2_out_31_port, data_in(30) => 
                           NPC2_out_30_port, data_in(29) => NPC2_out_29_port, 
                           data_in(28) => NPC2_out_28_port, data_in(27) => 
                           NPC2_out_27_port, data_in(26) => NPC2_out_26_port, 
                           data_in(25) => NPC2_out_25_port, data_in(24) => 
                           NPC2_out_24_port, data_in(23) => NPC2_out_23_port, 
                           data_in(22) => NPC2_out_22_port, data_in(21) => 
                           NPC2_out_21_port, data_in(20) => NPC2_out_20_port, 
                           data_in(19) => NPC2_out_19_port, data_in(18) => 
                           NPC2_out_18_port, data_in(17) => NPC2_out_17_port, 
                           data_in(16) => NPC2_out_16_port, data_in(15) => 
                           NPC2_out_15_port, data_in(14) => NPC2_out_14_port, 
                           data_in(13) => NPC2_out_13_port, data_in(12) => 
                           NPC2_out_12_port, data_in(11) => NPC2_out_11_port, 
                           data_in(10) => NPC2_out_10_port, data_in(9) => 
                           NPC2_out_9_port, data_in(8) => NPC2_out_8_port, 
                           data_in(7) => NPC2_out_7_port, data_in(6) => 
                           NPC2_out_6_port, data_in(5) => NPC2_out_5_port, 
                           data_in(4) => NPC2_out_4_port, data_in(3) => 
                           NPC2_out_3_port, data_in(2) => NPC2_out_2_port, 
                           data_in(1) => NPC2_out_1_port, data_in(0) => 
                           NPC2_out_0_port, data_out(31) => NPC3_out_31_port, 
                           data_out(30) => NPC3_out_30_port, data_out(29) => 
                           NPC3_out_29_port, data_out(28) => NPC3_out_28_port, 
                           data_out(27) => NPC3_out_27_port, data_out(26) => 
                           NPC3_out_26_port, data_out(25) => NPC3_out_25_port, 
                           data_out(24) => NPC3_out_24_port, data_out(23) => 
                           NPC3_out_23_port, data_out(22) => NPC3_out_22_port, 
                           data_out(21) => NPC3_out_21_port, data_out(20) => 
                           NPC3_out_20_port, data_out(19) => NPC3_out_19_port, 
                           data_out(18) => NPC3_out_18_port, data_out(17) => 
                           NPC3_out_17_port, data_out(16) => NPC3_out_16_port, 
                           data_out(15) => NPC3_out_15_port, data_out(14) => 
                           NPC3_out_14_port, data_out(13) => NPC3_out_13_port, 
                           data_out(12) => NPC3_out_12_port, data_out(11) => 
                           NPC3_out_11_port, data_out(10) => NPC3_out_10_port, 
                           data_out(9) => NPC3_out_9_port, data_out(8) => 
                           NPC3_out_8_port, data_out(7) => NPC3_out_7_port, 
                           data_out(6) => NPC3_out_6_port, data_out(5) => 
                           NPC3_out_5_port, data_out(4) => NPC3_out_4_port, 
                           data_out(3) => NPC3_out_3_port, data_out(2) => 
                           NPC3_out_2_port, data_out(1) => NPC3_out_1_port, 
                           data_out(0) => NPC3_out_0_port);
   RegPSW : REG_NBIT7 port map( clk => CLK, reset => n51, enable => n40, 
                           data_in(6) => PSW_in_6_port, data_in(5) => 
                           PSW_in_5_port, data_in(4) => PSW_in_4_port, 
                           data_in(3) => PSW_in_3_port, data_in(2) => 
                           PSW_in_2_port, data_in(1) => PSW_in_1_port, 
                           data_in(0) => PSW_in_0_port, data_out(6) => 
                           PSW_out_6_port, data_out(5) => PSW_out_5_port, 
                           data_out(4) => PSW_out_4_port, data_out(3) => 
                           PSW_out_3_port, data_out(2) => PSW_out_2_port, 
                           data_out(1) => PSW_out_1_port, data_out(0) => 
                           PSW_out_0_port);
   RegALR2 : REG_NBIT32_5 port map( clk => CLK, reset => n51, enable => n39, 
                           data_in(31) => ALR2_in_31_port, data_in(30) => 
                           ALR2_in_30_port, data_in(29) => ALR2_in_29_port, 
                           data_in(28) => ALR2_in_28_port, data_in(27) => 
                           ALR2_in_27_port, data_in(26) => ALR2_in_26_port, 
                           data_in(25) => ALR2_in_25_port, data_in(24) => 
                           ALR2_in_24_port, data_in(23) => ALR2_in_23_port, 
                           data_in(22) => ALR2_in_22_port, data_in(21) => 
                           ALR2_in_21_port, data_in(20) => ALR2_in_20_port, 
                           data_in(19) => ALR2_in_19_port, data_in(18) => 
                           ALR2_in_18_port, data_in(17) => ALR2_in_17_port, 
                           data_in(16) => ALR2_in_16_port, data_in(15) => 
                           ALR2_in_15_port, data_in(14) => ALR2_in_14_port, 
                           data_in(13) => ALR2_in_13_port, data_in(12) => 
                           ALR2_in_12_port, data_in(11) => ALR2_in_11_port, 
                           data_in(10) => ALR2_in_10_port, data_in(9) => 
                           ALR2_in_9_port, data_in(8) => ALR2_in_8_port, 
                           data_in(7) => ALR2_in_7_port, data_in(6) => 
                           ALR2_in_6_port, data_in(5) => ALR2_in_5_port, 
                           data_in(4) => ALR2_in_4_port, data_in(3) => 
                           ALR2_in_3_port, data_in(2) => ALR2_in_2_port, 
                           data_in(1) => ALR2_in_1_port, data_in(0) => 
                           ALR2_in_0_port, data_out(31) => ALR2_out_31_port, 
                           data_out(30) => ALR2_out_30_port, data_out(29) => 
                           ALR2_out_29_port, data_out(28) => ALR2_out_28_port, 
                           data_out(27) => ALR2_out_27_port, data_out(26) => 
                           ALR2_out_26_port, data_out(25) => ALR2_out_25_port, 
                           data_out(24) => ALR2_out_24_port, data_out(23) => 
                           ALR2_out_23_port, data_out(22) => ALR2_out_22_port, 
                           data_out(21) => ALR2_out_21_port, data_out(20) => 
                           ALR2_out_20_port, data_out(19) => ALR2_out_19_port, 
                           data_out(18) => ALR2_out_18_port, data_out(17) => 
                           ALR2_out_17_port, data_out(16) => ALR2_out_16_port, 
                           data_out(15) => ALR2_out_15_port, data_out(14) => 
                           ALR2_out_14_port, data_out(13) => ALR2_out_13_port, 
                           data_out(12) => ALR2_out_12_port, data_out(11) => 
                           ALR2_out_11_port, data_out(10) => ALR2_out_10_port, 
                           data_out(9) => ALR2_out_9_port, data_out(8) => 
                           ALR2_out_8_port, data_out(7) => ALR2_out_7_port, 
                           data_out(6) => ALR2_out_6_port, data_out(5) => 
                           ALR2_out_5_port, data_out(4) => ALR2_out_4_port, 
                           data_out(3) => ALR2_out_3_port, data_out(2) => 
                           ALR2_out_2_port, data_out(1) => ALR2_out_1_port, 
                           data_out(0) => ALR2_out_0_port);
   RegWB3 : REG_NBIT32_4 port map( clk => CLK, reset => n51, enable => n39, 
                           data_in(31) => RWB2_out_31_port, data_in(30) => 
                           RWB2_out_30_port, data_in(29) => RWB2_out_29_port, 
                           data_in(28) => RWB2_out_28_port, data_in(27) => 
                           RWB2_out_27_port, data_in(26) => RWB2_out_26_port, 
                           data_in(25) => RWB2_out_25_port, data_in(24) => 
                           RWB2_out_24_port, data_in(23) => RWB2_out_23_port, 
                           data_in(22) => RWB2_out_22_port, data_in(21) => 
                           RWB2_out_21_port, data_in(20) => RWB2_out_20_port, 
                           data_in(19) => RWB2_out_19_port, data_in(18) => 
                           RWB2_out_18_port, data_in(17) => RWB2_out_17_port, 
                           data_in(16) => RWB2_out_16_port, data_in(15) => 
                           RWB2_out_15_port, data_in(14) => RWB2_out_14_port, 
                           data_in(13) => RWB2_out_13_port, data_in(12) => 
                           RWB2_out_12_port, data_in(11) => RWB2_out_11_port, 
                           data_in(10) => RWB2_out_10_port, data_in(9) => 
                           RWB2_out_9_port, data_in(8) => RWB2_out_8_port, 
                           data_in(7) => RWB2_out_7_port, data_in(6) => 
                           RWB2_out_6_port, data_in(5) => RWB2_out_5_port, 
                           data_in(4) => RWB2_out_4_port, data_in(3) => 
                           RWB2_out_3_port, data_in(2) => RWB2_out_2_port, 
                           data_in(1) => RWB2_out_1_port, data_in(0) => 
                           RWB2_out_0_port, data_out(31) => n_1586, 
                           data_out(30) => n_1587, data_out(29) => n_1588, 
                           data_out(28) => n_1589, data_out(27) => n_1590, 
                           data_out(26) => n_1591, data_out(25) => n_1592, 
                           data_out(24) => n_1593, data_out(23) => n_1594, 
                           data_out(22) => n_1595, data_out(21) => n_1596, 
                           data_out(20) => RWB3_out_20_port, data_out(19) => 
                           RWB3_out_19_port, data_out(18) => RWB3_out_18_port, 
                           data_out(17) => RWB3_out_17_port, data_out(16) => 
                           RWB3_out_16_port, data_out(15) => RWB3_out_15_port, 
                           data_out(14) => RWB3_out_14_port, data_out(13) => 
                           RWB3_out_13_port, data_out(12) => RWB3_out_12_port, 
                           data_out(11) => RWB3_out_11_port, data_out(10) => 
                           n_1597, data_out(9) => n_1598, data_out(8) => n_1599
                           , data_out(7) => n_1600, data_out(6) => n_1601, 
                           data_out(5) => n_1602, data_out(4) => n_1603, 
                           data_out(3) => n_1604, data_out(2) => n_1605, 
                           data_out(1) => n_1606, data_out(0) => n_1607);
   AdderPC : PC_adder_0 port map( A(31) => IRAM_ADDR_31_port, A(30) => 
                           IRAM_ADDR_30_port, A(29) => IRAM_ADDR_29_port, A(28)
                           => IRAM_ADDR_28_port, A(27) => IRAM_ADDR_27_port, 
                           A(26) => IRAM_ADDR_26_port, A(25) => 
                           IRAM_ADDR_25_port, A(24) => IRAM_ADDR_24_port, A(23)
                           => IRAM_ADDR_23_port, A(22) => IRAM_ADDR_22_port, 
                           A(21) => IRAM_ADDR_21_port, A(20) => 
                           IRAM_ADDR_20_port, A(19) => IRAM_ADDR_19_port, A(18)
                           => IRAM_ADDR_18_port, A(17) => IRAM_ADDR_17_port, 
                           A(16) => IRAM_ADDR_16_port, A(15) => 
                           IRAM_ADDR_15_port, A(14) => IRAM_ADDR_14_port, A(13)
                           => IRAM_ADDR_13_port, A(12) => IRAM_ADDR_12_port, 
                           A(11) => IRAM_ADDR_11_port, A(10) => 
                           IRAM_ADDR_10_port, A(9) => IRAM_ADDR_9_port, A(8) =>
                           IRAM_ADDR_8_port, A(7) => IRAM_ADDR_7_port, A(6) => 
                           IRAM_ADDR_6_port, A(5) => IRAM_ADDR_5_port, A(4) => 
                           IRAM_ADDR_4_port, A(3) => IRAM_ADDR_3_port, A(2) => 
                           IRAM_ADDR_2_port, A(1) => IRAM_ADDR_1_port, A(0) => 
                           IRAM_ADDR_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, Sum(31) => NPC_in_31_port, Sum(30) =>
                           NPC_in_30_port, Sum(29) => NPC_in_29_port, Sum(28) 
                           => NPC_in_28_port, Sum(27) => NPC_in_27_port, 
                           Sum(26) => NPC_in_26_port, Sum(25) => NPC_in_25_port
                           , Sum(24) => NPC_in_24_port, Sum(23) => 
                           NPC_in_23_port, Sum(22) => NPC_in_22_port, Sum(21) 
                           => NPC_in_21_port, Sum(20) => NPC_in_20_port, 
                           Sum(19) => NPC_in_19_port, Sum(18) => NPC_in_18_port
                           , Sum(17) => NPC_in_17_port, Sum(16) => 
                           NPC_in_16_port, Sum(15) => NPC_in_15_port, Sum(14) 
                           => NPC_in_14_port, Sum(13) => NPC_in_13_port, 
                           Sum(12) => NPC_in_12_port, Sum(11) => NPC_in_11_port
                           , Sum(10) => NPC_in_10_port, Sum(9) => NPC_in_9_port
                           , Sum(8) => NPC_in_8_port, Sum(7) => NPC_in_7_port, 
                           Sum(6) => NPC_in_6_port, Sum(5) => NPC_in_5_port, 
                           Sum(4) => NPC_in_4_port, Sum(3) => NPC_in_3_port, 
                           Sum(2) => NPC_in_2_port, Sum(1) => NPC_in_1_port, 
                           Sum(0) => NPC_in_0_port);
   J_Adder : PC_adder_1 port map( A(31) => PC2_out_31_port, A(30) => 
                           PC2_out_30_port, A(29) => PC2_out_29_port, A(28) => 
                           PC2_out_28_port, A(27) => PC2_out_27_port, A(26) => 
                           PC2_out_26_port, A(25) => PC2_out_25_port, A(24) => 
                           PC2_out_24_port, A(23) => PC2_out_23_port, A(22) => 
                           PC2_out_22_port, A(21) => PC2_out_21_port, A(20) => 
                           PC2_out_20_port, A(19) => PC2_out_19_port, A(18) => 
                           PC2_out_18_port, A(17) => PC2_out_17_port, A(16) => 
                           PC2_out_16_port, A(15) => PC2_out_15_port, A(14) => 
                           PC2_out_14_port, A(13) => PC2_out_13_port, A(12) => 
                           PC2_out_12_port, A(11) => PC2_out_11_port, A(10) => 
                           PC2_out_10_port, A(9) => PC2_out_9_port, A(8) => 
                           PC2_out_8_port, A(7) => PC2_out_7_port, A(6) => 
                           PC2_out_6_port, A(5) => PC2_out_5_port, A(4) => 
                           PC2_out_4_port, A(3) => PC2_out_3_port, A(2) => 
                           PC2_out_2_port, A(1) => PC2_out_1_port, A(0) => 
                           PC2_out_0_port, B(31) => IMM_out_31_port, B(30) => 
                           IMM_out_30_port, B(29) => IMM_out_29_port, B(28) => 
                           IMM_out_28_port, B(27) => IMM_out_27_port, B(26) => 
                           IMM_out_26_port, B(25) => IMM_out_25_port, B(24) => 
                           IMM_out_24_port, B(23) => IMM_out_23_port, B(22) => 
                           IMM_out_22_port, B(21) => IMM_out_21_port, B(20) => 
                           IMM_out_20_port, B(19) => IMM_out_19_port, B(18) => 
                           IMM_out_18_port, B(17) => IMM_out_17_port, B(16) => 
                           IMM_out_16_port, B(15) => IMM_out_15_port, B(14) => 
                           IMM_out_14_port, B(13) => IMM_out_13_port, B(12) => 
                           IMM_out_12_port, B(11) => IMM_out_11_port, B(10) => 
                           IMM_out_10_port, B(9) => IMM_out_9_port, B(8) => 
                           IMM_out_8_port, B(7) => IMM_out_7_port, B(6) => 
                           IMM_out_6_port, B(5) => IMM_out_5_port, B(4) => 
                           IMM_out_4_port, B(3) => IMM_out_3_port, B(2) => 
                           IMM_out_2_port, B(1) => IMM_out_1_port, B(0) => 
                           IMM_out_0_port, Sum(31) => JADDER_out_31_port, 
                           Sum(30) => JADDER_out_30_port, Sum(29) => 
                           JADDER_out_29_port, Sum(28) => JADDER_out_28_port, 
                           Sum(27) => JADDER_out_27_port, Sum(26) => 
                           JADDER_out_26_port, Sum(25) => JADDER_out_25_port, 
                           Sum(24) => JADDER_out_24_port, Sum(23) => 
                           JADDER_out_23_port, Sum(22) => JADDER_out_22_port, 
                           Sum(21) => JADDER_out_21_port, Sum(20) => 
                           JADDER_out_20_port, Sum(19) => JADDER_out_19_port, 
                           Sum(18) => JADDER_out_18_port, Sum(17) => 
                           JADDER_out_17_port, Sum(16) => JADDER_out_16_port, 
                           Sum(15) => JADDER_out_15_port, Sum(14) => 
                           JADDER_out_14_port, Sum(13) => JADDER_out_13_port, 
                           Sum(12) => JADDER_out_12_port, Sum(11) => 
                           JADDER_out_11_port, Sum(10) => JADDER_out_10_port, 
                           Sum(9) => JADDER_out_9_port, Sum(8) => 
                           JADDER_out_8_port, Sum(7) => JADDER_out_7_port, 
                           Sum(6) => JADDER_out_6_port, Sum(5) => 
                           JADDER_out_5_port, Sum(4) => JADDER_out_4_port, 
                           Sum(3) => JADDER_out_3_port, Sum(2) => 
                           JADDER_out_2_port, Sum(1) => JADDER_out_1_port, 
                           Sum(0) => JADDER_out_0_port);
   PCMUX : MUX3to1_NBIT32_0 port map( A(31) => PC_out_31_port, A(30) => 
                           PC_out_30_port, A(29) => PC_out_29_port, A(28) => 
                           PC_out_28_port, A(27) => PC_out_27_port, A(26) => 
                           PC_out_26_port, A(25) => PC_out_25_port, A(24) => 
                           PC_out_24_port, A(23) => PC_out_23_port, A(22) => 
                           PC_out_22_port, A(21) => PC_out_21_port, A(20) => 
                           PC_out_20_port, A(19) => PC_out_19_port, A(18) => 
                           PC_out_18_port, A(17) => PC_out_17_port, A(16) => 
                           PC_out_16_port, A(15) => PC_out_15_port, A(14) => 
                           PC_out_14_port, A(13) => PC_out_13_port, A(12) => 
                           PC_out_12_port, A(11) => PC_out_11_port, A(10) => 
                           PC_out_10_port, A(9) => PC_out_9_port, A(8) => 
                           PC_out_8_port, A(7) => PC_out_7_port, A(6) => 
                           PC_out_6_port, A(5) => PC_out_5_port, A(4) => 
                           PC_out_4_port, A(3) => PC_out_3_port, A(2) => 
                           PC_out_2_port, A(1) => PC_out_1_port, A(0) => 
                           PC_out_0_port, B(31) => JADDER_out_31_port, B(30) =>
                           JADDER_out_30_port, B(29) => JADDER_out_29_port, 
                           B(28) => JADDER_out_28_port, B(27) => 
                           JADDER_out_27_port, B(26) => JADDER_out_26_port, 
                           B(25) => JADDER_out_25_port, B(24) => 
                           JADDER_out_24_port, B(23) => JADDER_out_23_port, 
                           B(22) => JADDER_out_22_port, B(21) => 
                           JADDER_out_21_port, B(20) => JADDER_out_20_port, 
                           B(19) => JADDER_out_19_port, B(18) => 
                           JADDER_out_18_port, B(17) => JADDER_out_17_port, 
                           B(16) => JADDER_out_16_port, B(15) => 
                           JADDER_out_15_port, B(14) => JADDER_out_14_port, 
                           B(13) => JADDER_out_13_port, B(12) => 
                           JADDER_out_12_port, B(11) => JADDER_out_11_port, 
                           B(10) => JADDER_out_10_port, B(9) => 
                           JADDER_out_9_port, B(8) => JADDER_out_8_port, B(7) 
                           => JADDER_out_7_port, B(6) => JADDER_out_6_port, 
                           B(5) => JADDER_out_5_port, B(4) => JADDER_out_4_port
                           , B(3) => JADDER_out_3_port, B(2) => 
                           JADDER_out_2_port, B(1) => JADDER_out_1_port, B(0) 
                           => JADDER_out_0_port, C(31) => JADDER2_out_31_port, 
                           C(30) => JADDER2_out_30_port, C(29) => 
                           JADDER2_out_29_port, C(28) => JADDER2_out_28_port, 
                           C(27) => JADDER2_out_27_port, C(26) => 
                           JADDER2_out_26_port, C(25) => JADDER2_out_25_port, 
                           C(24) => JADDER2_out_24_port, C(23) => 
                           JADDER2_out_23_port, C(22) => JADDER2_out_22_port, 
                           C(21) => JADDER2_out_21_port, C(20) => 
                           JADDER2_out_20_port, C(19) => JADDER2_out_19_port, 
                           C(18) => JADDER2_out_18_port, C(17) => 
                           JADDER2_out_17_port, C(16) => JADDER2_out_16_port, 
                           C(15) => JADDER2_out_15_port, C(14) => 
                           JADDER2_out_14_port, C(13) => JADDER2_out_13_port, 
                           C(12) => JADDER2_out_12_port, C(11) => 
                           JADDER2_out_11_port, C(10) => JADDER2_out_10_port, 
                           C(9) => JADDER2_out_9_port, C(8) => 
                           JADDER2_out_8_port, C(7) => JADDER2_out_7_port, C(6)
                           => JADDER2_out_6_port, C(5) => JADDER2_out_5_port, 
                           C(4) => JADDER2_out_4_port, C(3) => 
                           JADDER2_out_3_port, C(2) => JADDER2_out_2_port, C(1)
                           => JADDER2_out_1_port, C(0) => JADDER2_out_0_port, 
                           SEL(1) => PC_SEL_1_port, SEL(0) => n52, Y(31) => 
                           PC_MUX_out_31_port, Y(30) => PC_MUX_out_30_port, 
                           Y(29) => PC_MUX_out_29_port, Y(28) => 
                           PC_MUX_out_28_port, Y(27) => PC_MUX_out_27_port, 
                           Y(26) => PC_MUX_out_26_port, Y(25) => 
                           PC_MUX_out_25_port, Y(24) => PC_MUX_out_24_port, 
                           Y(23) => PC_MUX_out_23_port, Y(22) => 
                           PC_MUX_out_22_port, Y(21) => PC_MUX_out_21_port, 
                           Y(20) => PC_MUX_out_20_port, Y(19) => 
                           PC_MUX_out_19_port, Y(18) => PC_MUX_out_18_port, 
                           Y(17) => PC_MUX_out_17_port, Y(16) => 
                           PC_MUX_out_16_port, Y(15) => PC_MUX_out_15_port, 
                           Y(14) => PC_MUX_out_14_port, Y(13) => 
                           PC_MUX_out_13_port, Y(12) => PC_MUX_out_12_port, 
                           Y(11) => PC_MUX_out_11_port, Y(10) => 
                           PC_MUX_out_10_port, Y(9) => PC_MUX_out_9_port, Y(8) 
                           => PC_MUX_out_8_port, Y(7) => PC_MUX_out_7_port, 
                           Y(6) => PC_MUX_out_6_port, Y(5) => PC_MUX_out_5_port
                           , Y(4) => PC_MUX_out_4_port, Y(3) => 
                           PC_MUX_out_3_port, Y(2) => PC_MUX_out_2_port, Y(1) 
                           => PC_MUX_out_1_port, Y(0) => PC_MUX_out_0_port);
   IRAMMUX : MUX2to1_NBIT32_0 port map( A(31) => PC_MUX_out_31_port, A(30) => 
                           PC_MUX_out_30_port, A(29) => PC_MUX_out_29_port, 
                           A(28) => PC_MUX_out_28_port, A(27) => 
                           PC_MUX_out_27_port, A(26) => PC_MUX_out_26_port, 
                           A(25) => PC_MUX_out_25_port, A(24) => 
                           PC_MUX_out_24_port, A(23) => PC_MUX_out_23_port, 
                           A(22) => PC_MUX_out_22_port, A(21) => 
                           PC_MUX_out_21_port, A(20) => PC_MUX_out_20_port, 
                           A(19) => PC_MUX_out_19_port, A(18) => 
                           PC_MUX_out_18_port, A(17) => PC_MUX_out_17_port, 
                           A(16) => PC_MUX_out_16_port, A(15) => 
                           PC_MUX_out_15_port, A(14) => PC_MUX_out_14_port, 
                           A(13) => PC_MUX_out_13_port, A(12) => 
                           PC_MUX_out_12_port, A(11) => PC_MUX_out_11_port, 
                           A(10) => PC_MUX_out_10_port, A(9) => 
                           PC_MUX_out_9_port, A(8) => PC_MUX_out_8_port, A(7) 
                           => PC_MUX_out_7_port, A(6) => PC_MUX_out_6_port, 
                           A(5) => PC_MUX_out_5_port, A(4) => PC_MUX_out_4_port
                           , A(3) => PC_MUX_out_3_port, A(2) => 
                           PC_MUX_out_2_port, A(1) => PC_MUX_out_1_port, A(0) 
                           => PC_MUX_out_0_port, B(31) => NPC2_out_31_port, 
                           B(30) => NPC2_out_30_port, B(29) => NPC2_out_29_port
                           , B(28) => NPC2_out_28_port, B(27) => 
                           NPC2_out_27_port, B(26) => NPC2_out_26_port, B(25) 
                           => NPC2_out_25_port, B(24) => NPC2_out_24_port, 
                           B(23) => NPC2_out_23_port, B(22) => NPC2_out_22_port
                           , B(21) => NPC2_out_21_port, B(20) => 
                           NPC2_out_20_port, B(19) => NPC2_out_19_port, B(18) 
                           => NPC2_out_18_port, B(17) => NPC2_out_17_port, 
                           B(16) => NPC2_out_16_port, B(15) => NPC2_out_15_port
                           , B(14) => NPC2_out_14_port, B(13) => 
                           NPC2_out_13_port, B(12) => NPC2_out_12_port, B(11) 
                           => NPC2_out_11_port, B(10) => NPC2_out_10_port, B(9)
                           => NPC2_out_9_port, B(8) => NPC2_out_8_port, B(7) =>
                           NPC2_out_7_port, B(6) => NPC2_out_6_port, B(5) => 
                           NPC2_out_5_port, B(4) => NPC2_out_4_port, B(3) => 
                           NPC2_out_3_port, B(2) => NPC2_out_2_port, B(1) => 
                           NPC2_out_1_port, B(0) => NPC2_out_0_port, SEL => 
                           IRAMMUX_SEL, Y(31) => IRAM_ADDR_31_port, Y(30) => 
                           IRAM_ADDR_30_port, Y(29) => IRAM_ADDR_29_port, Y(28)
                           => IRAM_ADDR_28_port, Y(27) => IRAM_ADDR_27_port, 
                           Y(26) => IRAM_ADDR_26_port, Y(25) => 
                           IRAM_ADDR_25_port, Y(24) => IRAM_ADDR_24_port, Y(23)
                           => IRAM_ADDR_23_port, Y(22) => IRAM_ADDR_22_port, 
                           Y(21) => IRAM_ADDR_21_port, Y(20) => 
                           IRAM_ADDR_20_port, Y(19) => IRAM_ADDR_19_port, Y(18)
                           => IRAM_ADDR_18_port, Y(17) => IRAM_ADDR_17_port, 
                           Y(16) => IRAM_ADDR_16_port, Y(15) => 
                           IRAM_ADDR_15_port, Y(14) => IRAM_ADDR_14_port, Y(13)
                           => IRAM_ADDR_13_port, Y(12) => IRAM_ADDR_12_port, 
                           Y(11) => IRAM_ADDR_11_port, Y(10) => 
                           IRAM_ADDR_10_port, Y(9) => IRAM_ADDR_9_port, Y(8) =>
                           IRAM_ADDR_8_port, Y(7) => IRAM_ADDR_7_port, Y(6) => 
                           IRAM_ADDR_6_port, Y(5) => IRAM_ADDR_5_port, Y(4) => 
                           IRAM_ADDR_4_port, Y(3) => IRAM_ADDR_3_port, Y(2) => 
                           IRAM_ADDR_2_port, Y(1) => IRAM_ADDR_1_port, Y(0) => 
                           IRAM_ADDR_0_port);
   IMMMUX : MUX2to1_NBIT32_8 port map( A(31) => IR_out_15_port, A(30) => 
                           IR_out_15_port, A(29) => IR_out_15_port, A(28) => 
                           IR_out_15_port, A(27) => IR_out_15_port, A(26) => 
                           IR_out_15_port, A(25) => IR_out_15_port, A(24) => 
                           IR_out_15_port, A(23) => IR_out_15_port, A(22) => 
                           IR_out_15_port, A(21) => IR_out_15_port, A(20) => 
                           IR_out_15_port, A(19) => IR_out_15_port, A(18) => 
                           IR_out_15_port, A(17) => IR_out_15_port, A(16) => 
                           IR_out_15_port, A(15) => IR_out_15_port, A(14) => 
                           IR_out_14_port, A(13) => IR_out_13_port, A(12) => 
                           IR_out_12_port, A(11) => IR_out_11_port, A(10) => 
                           IR_out_10_port, A(9) => IR_out_9_port, A(8) => 
                           IR_out_8_port, A(7) => IR_out_7_port, A(6) => 
                           IR_out_6_port, A(5) => IR_out_5_port, A(4) => 
                           IR_out_4_port, A(3) => IR_out_3_port, A(2) => 
                           IR_out_2_port, A(1) => IR_out_1_port, A(0) => 
                           IR_out_0_port, B(31) => IR_out_25_port, B(30) => 
                           IR_out_25_port, B(29) => IR_out_25_port, B(28) => 
                           IR_out_25_port, B(27) => IR_out_25_port, B(26) => 
                           IR_out_25_port, B(25) => IR_out_25_port, B(24) => 
                           IR_out_24_port, B(23) => IR_out_23_port, B(22) => 
                           IR_out_22_port, B(21) => IR_out_21_port, B(20) => 
                           IR_out_20_port, B(19) => IR_out_19_port, B(18) => 
                           n36, B(17) => IR_out_17_port, B(16) => 
                           IR_out_16_port, B(15) => IR_out_15_port, B(14) => 
                           IR_out_14_port, B(13) => IR_out_13_port, B(12) => 
                           IR_out_12_port, B(11) => IR_out_11_port, B(10) => 
                           IR_out_10_port, B(9) => IR_out_9_port, B(8) => 
                           IR_out_8_port, B(7) => IR_out_7_port, B(6) => 
                           IR_out_6_port, B(5) => IR_out_5_port, B(4) => 
                           IR_out_4_port, B(3) => IR_out_3_port, B(2) => 
                           IR_out_2_port, B(1) => IR_out_1_port, B(0) => 
                           IR_out_0_port, SEL => IMM_SEL, Y(31) => 
                           IMM_out_31_port, Y(30) => IMM_out_30_port, Y(29) => 
                           IMM_out_29_port, Y(28) => IMM_out_28_port, Y(27) => 
                           IMM_out_27_port, Y(26) => IMM_out_26_port, Y(25) => 
                           IMM_out_25_port, Y(24) => IMM_out_24_port, Y(23) => 
                           IMM_out_23_port, Y(22) => IMM_out_22_port, Y(21) => 
                           IMM_out_21_port, Y(20) => IMM_out_20_port, Y(19) => 
                           IMM_out_19_port, Y(18) => IMM_out_18_port, Y(17) => 
                           IMM_out_17_port, Y(16) => IMM_out_16_port, Y(15) => 
                           IMM_out_15_port, Y(14) => IMM_out_14_port, Y(13) => 
                           IMM_out_13_port, Y(12) => IMM_out_12_port, Y(11) => 
                           IMM_out_11_port, Y(10) => IMM_out_10_port, Y(9) => 
                           IMM_out_9_port, Y(8) => IMM_out_8_port, Y(7) => 
                           IMM_out_7_port, Y(6) => IMM_out_6_port, Y(5) => 
                           IMM_out_5_port, Y(4) => IMM_out_4_port, Y(3) => 
                           IMM_out_3_port, Y(2) => IMM_out_2_port, Y(1) => 
                           IMM_out_1_port, Y(0) => IMM_out_0_port);
   BHTMUX : MUX2to1_NBIT32_7 port map( A(31) => PC2_out_31_port, A(30) => 
                           PC2_out_30_port, A(29) => PC2_out_29_port, A(28) => 
                           PC2_out_28_port, A(27) => PC2_out_27_port, A(26) => 
                           PC2_out_26_port, A(25) => PC2_out_25_port, A(24) => 
                           PC2_out_24_port, A(23) => PC2_out_23_port, A(22) => 
                           PC2_out_22_port, A(21) => PC2_out_21_port, A(20) => 
                           PC2_out_20_port, A(19) => PC2_out_19_port, A(18) => 
                           PC2_out_18_port, A(17) => PC2_out_17_port, A(16) => 
                           PC2_out_16_port, A(15) => PC2_out_15_port, A(14) => 
                           PC2_out_14_port, A(13) => PC2_out_13_port, A(12) => 
                           PC2_out_12_port, A(11) => PC2_out_11_port, A(10) => 
                           PC2_out_10_port, A(9) => PC2_out_9_port, A(8) => 
                           PC2_out_8_port, A(7) => PC2_out_7_port, A(6) => 
                           PC2_out_6_port, A(5) => PC2_out_5_port, A(4) => 
                           PC2_out_4_port, A(3) => PC2_out_3_port, A(2) => 
                           PC2_out_2_port, A(1) => PC2_out_1_port, A(0) => 
                           PC2_out_0_port, B(31) => PC3_out_31_port, B(30) => 
                           PC3_out_30_port, B(29) => PC3_out_29_port, B(28) => 
                           PC3_out_28_port, B(27) => PC3_out_27_port, B(26) => 
                           PC3_out_26_port, B(25) => PC3_out_25_port, B(24) => 
                           PC3_out_24_port, B(23) => PC3_out_23_port, B(22) => 
                           PC3_out_22_port, B(21) => PC3_out_21_port, B(20) => 
                           PC3_out_20_port, B(19) => PC3_out_19_port, B(18) => 
                           PC3_out_18_port, B(17) => PC3_out_17_port, B(16) => 
                           PC3_out_16_port, B(15) => PC3_out_15_port, B(14) => 
                           PC3_out_14_port, B(13) => PC3_out_13_port, B(12) => 
                           PC3_out_12_port, B(11) => PC3_out_11_port, B(10) => 
                           PC3_out_10_port, B(9) => PC3_out_9_port, B(8) => 
                           PC3_out_8_port, B(7) => PC3_out_7_port, B(6) => 
                           PC3_out_6_port, B(5) => PC3_out_5_port, B(4) => 
                           PC3_out_4_port, B(3) => PC3_out_3_port, B(2) => 
                           PC3_out_2_port, B(1) => PC3_out_1_port, B(0) => 
                           PC3_out_0_port, SEL => BPR_EN2, Y(31) => 
                           BHT_in_31_port, Y(30) => BHT_in_30_port, Y(29) => 
                           BHT_in_29_port, Y(28) => BHT_in_28_port, Y(27) => 
                           BHT_in_27_port, Y(26) => BHT_in_26_port, Y(25) => 
                           BHT_in_25_port, Y(24) => BHT_in_24_port, Y(23) => 
                           BHT_in_23_port, Y(22) => BHT_in_22_port, Y(21) => 
                           BHT_in_21_port, Y(20) => BHT_in_20_port, Y(19) => 
                           BHT_in_19_port, Y(18) => BHT_in_18_port, Y(17) => 
                           BHT_in_17_port, Y(16) => BHT_in_16_port, Y(15) => 
                           BHT_in_15_port, Y(14) => BHT_in_14_port, Y(13) => 
                           BHT_in_13_port, Y(12) => BHT_in_12_port, Y(11) => 
                           BHT_in_11_port, Y(10) => BHT_in_10_port, Y(9) => 
                           BHT_in_9_port, Y(8) => BHT_in_8_port, Y(7) => 
                           BHT_in_7_port, Y(6) => BHT_in_6_port, Y(5) => 
                           BHT_in_5_port, Y(4) => BHT_in_4_port, Y(3) => 
                           BHT_in_3_port, Y(2) => BHT_in_2_port, Y(1) => 
                           BHT_in_1_port, Y(0) => BHT_in_0_port);
   RegAMUX : MUX2to1_NBIT32_6 port map( A(31) => FWDA_OUT_31_port, A(30) => 
                           FWDA_OUT_30_port, A(29) => FWDA_OUT_29_port, A(28) 
                           => FWDA_OUT_28_port, A(27) => FWDA_OUT_27_port, 
                           A(26) => FWDA_OUT_26_port, A(25) => FWDA_OUT_25_port
                           , A(24) => FWDA_OUT_24_port, A(23) => 
                           FWDA_OUT_23_port, A(22) => FWDA_OUT_22_port, A(21) 
                           => FWDA_OUT_21_port, A(20) => FWDA_OUT_20_port, 
                           A(19) => FWDA_OUT_19_port, A(18) => FWDA_OUT_18_port
                           , A(17) => FWDA_OUT_17_port, A(16) => 
                           FWDA_OUT_16_port, A(15) => FWDA_OUT_15_port, A(14) 
                           => FWDA_OUT_14_port, A(13) => FWDA_OUT_13_port, 
                           A(12) => FWDA_OUT_12_port, A(11) => FWDA_OUT_11_port
                           , A(10) => FWDA_OUT_10_port, A(9) => FWDA_OUT_9_port
                           , A(8) => FWDA_OUT_8_port, A(7) => FWDA_OUT_7_port, 
                           A(6) => FWDA_OUT_6_port, A(5) => FWDA_OUT_5_port, 
                           A(4) => FWDA_OUT_4_port, A(3) => FWDA_OUT_3_port, 
                           A(2) => FWDA_OUT_2_port, A(1) => FWDA_OUT_1_port, 
                           A(0) => FWDA_OUT_0_port, B(31) => X_Logic0_port, 
                           B(30) => X_Logic0_port, B(29) => X_Logic0_port, 
                           B(28) => X_Logic0_port, B(27) => X_Logic0_port, 
                           B(26) => X_Logic0_port, B(25) => X_Logic0_port, 
                           B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
                           B(22) => X_Logic0_port, B(21) => X_Logic0_port, 
                           B(20) => X_Logic0_port, B(19) => X_Logic0_port, 
                           B(18) => X_Logic0_port, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => X_Logic0_port, 
                           B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
                           B(12) => X_Logic0_port, B(11) => X_Logic0_port, 
                           B(10) => X_Logic0_port, B(9) => X_Logic0_port, B(8) 
                           => X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => ALUA_SEL, Y(31) => 
                           A_in_31_port, Y(30) => A_in_30_port, Y(29) => 
                           A_in_29_port, Y(28) => A_in_28_port, Y(27) => 
                           A_in_27_port, Y(26) => A_in_26_port, Y(25) => 
                           A_in_25_port, Y(24) => A_in_24_port, Y(23) => 
                           A_in_23_port, Y(22) => A_in_22_port, Y(21) => 
                           A_in_21_port, Y(20) => A_in_20_port, Y(19) => 
                           A_in_19_port, Y(18) => A_in_18_port, Y(17) => 
                           A_in_17_port, Y(16) => A_in_16_port, Y(15) => 
                           A_in_15_port, Y(14) => A_in_14_port, Y(13) => 
                           A_in_13_port, Y(12) => A_in_12_port, Y(11) => 
                           A_in_11_port, Y(10) => A_in_10_port, Y(9) => 
                           A_in_9_port, Y(8) => A_in_8_port, Y(7) => 
                           A_in_7_port, Y(6) => A_in_6_port, Y(5) => 
                           A_in_5_port, Y(4) => A_in_4_port, Y(3) => 
                           A_in_3_port, Y(2) => A_in_2_port, Y(1) => 
                           A_in_1_port, Y(0) => A_in_0_port);
   RegBMUX : MUX2to1_NBIT32_5 port map( A(31) => FWDB_OUT_31_port, A(30) => 
                           FWDB_OUT_30_port, A(29) => FWDB_OUT_29_port, A(28) 
                           => FWDB_OUT_28_port, A(27) => FWDB_OUT_27_port, 
                           A(26) => FWDB_OUT_26_port, A(25) => FWDB_OUT_25_port
                           , A(24) => FWDB_OUT_24_port, A(23) => 
                           FWDB_OUT_23_port, A(22) => FWDB_OUT_22_port, A(21) 
                           => FWDB_OUT_21_port, A(20) => FWDB_OUT_20_port, 
                           A(19) => FWDB_OUT_19_port, A(18) => FWDB_OUT_18_port
                           , A(17) => FWDB_OUT_17_port, A(16) => 
                           FWDB_OUT_16_port, A(15) => FWDB_OUT_15_port, A(14) 
                           => FWDB_OUT_14_port, A(13) => FWDB_OUT_13_port, 
                           A(12) => FWDB_OUT_12_port, A(11) => FWDB_OUT_11_port
                           , A(10) => FWDB_OUT_10_port, A(9) => FWDB_OUT_9_port
                           , A(8) => FWDB_OUT_8_port, A(7) => FWDB_OUT_7_port, 
                           A(6) => FWDB_OUT_6_port, A(5) => FWDB_OUT_5_port, 
                           A(4) => FWDB_OUT_4_port, A(3) => FWDB_OUT_3_port, 
                           A(2) => FWDB_OUT_2_port, A(1) => FWDB_OUT_1_port, 
                           A(0) => FWDB_OUT_0_port, B(31) => RIMM_out_31_port, 
                           B(30) => RIMM_out_30_port, B(29) => RIMM_out_29_port
                           , B(28) => RIMM_out_28_port, B(27) => 
                           RIMM_out_27_port, B(26) => RIMM_out_26_port, B(25) 
                           => RIMM_out_25_port, B(24) => RIMM_out_24_port, 
                           B(23) => RIMM_out_23_port, B(22) => RIMM_out_22_port
                           , B(21) => RIMM_out_21_port, B(20) => 
                           RIMM_out_20_port, B(19) => RIMM_out_19_port, B(18) 
                           => RIMM_out_18_port, B(17) => RIMM_out_17_port, 
                           B(16) => RIMM_out_16_port, B(15) => RIMM_out_15_port
                           , B(14) => RIMM_out_14_port, B(13) => 
                           RIMM_out_13_port, B(12) => RIMM_out_12_port, B(11) 
                           => RIMM_out_11_port, B(10) => RIMM_out_10_port, B(9)
                           => RIMM_out_9_port, B(8) => RIMM_out_8_port, B(7) =>
                           RIMM_out_7_port, B(6) => RIMM_out_6_port, B(5) => 
                           RIMM_out_5_port, B(4) => RIMM_out_4_port, B(3) => 
                           RIMM_out_3_port, B(2) => RIMM_out_2_port, B(1) => 
                           RIMM_out_1_port, B(0) => RIMM_out_0_port, SEL => 
                           ALUB_SEL, Y(31) => B_in_31_port, Y(30) => 
                           B_in_30_port, Y(29) => B_in_29_port, Y(28) => 
                           B_in_28_port, Y(27) => B_in_27_port, Y(26) => 
                           B_in_26_port, Y(25) => B_in_25_port, Y(24) => 
                           B_in_24_port, Y(23) => B_in_23_port, Y(22) => 
                           B_in_22_port, Y(21) => B_in_21_port, Y(20) => 
                           B_in_20_port, Y(19) => B_in_19_port, Y(18) => 
                           B_in_18_port, Y(17) => B_in_17_port, Y(16) => 
                           B_in_16_port, Y(15) => B_in_15_port, Y(14) => 
                           B_in_14_port, Y(13) => B_in_13_port, Y(12) => 
                           B_in_12_port, Y(11) => B_in_11_port, Y(10) => 
                           B_in_10_port, Y(9) => B_in_9_port, Y(8) => 
                           B_in_8_port, Y(7) => B_in_7_port, Y(6) => 
                           B_in_6_port, Y(5) => B_in_5_port, Y(4) => 
                           B_in_4_port, Y(3) => B_in_3_port, Y(2) => 
                           B_in_2_port, Y(1) => B_in_1_port, Y(0) => 
                           B_in_0_port);
   FWDA_MUX : MUX3to1_NBIT32_3 port map( A(31) => RA_out_31_port, A(30) => 
                           RA_out_30_port, A(29) => RA_out_29_port, A(28) => 
                           RA_out_28_port, A(27) => RA_out_27_port, A(26) => 
                           RA_out_26_port, A(25) => RA_out_25_port, A(24) => 
                           RA_out_24_port, A(23) => RA_out_23_port, A(22) => 
                           RA_out_22_port, A(21) => RA_out_21_port, A(20) => 
                           RA_out_20_port, A(19) => RA_out_19_port, A(18) => 
                           RA_out_18_port, A(17) => RA_out_17_port, A(16) => 
                           RA_out_16_port, A(15) => RA_out_15_port, A(14) => 
                           RA_out_14_port, A(13) => RA_out_13_port, A(12) => 
                           RA_out_12_port, A(11) => RA_out_11_port, A(10) => 
                           RA_out_10_port, A(9) => RA_out_9_port, A(8) => 
                           RA_out_8_port, A(7) => RA_out_7_port, A(6) => 
                           RA_out_6_port, A(5) => RA_out_5_port, A(4) => 
                           RA_out_4_port, A(3) => RA_out_3_port, A(2) => 
                           RA_out_2_port, A(1) => RA_out_1_port, A(0) => 
                           RA_out_0_port, B(31) => DATA_ADDR_31_port, B(30) => 
                           DATA_ADDR_30_port, B(29) => DATA_ADDR_29_port, B(28)
                           => DATA_ADDR_28_port, B(27) => DATA_ADDR_27_port, 
                           B(26) => DATA_ADDR_26_port, B(25) => 
                           DATA_ADDR_25_port, B(24) => DATA_ADDR_24_port, B(23)
                           => DATA_ADDR_23_port, B(22) => DATA_ADDR_22_port, 
                           B(21) => DATA_ADDR_21_port, B(20) => 
                           DATA_ADDR_20_port, B(19) => DATA_ADDR_19_port, B(18)
                           => DATA_ADDR_18_port, B(17) => DATA_ADDR_17_port, 
                           B(16) => DATA_ADDR_16_port, B(15) => 
                           DATA_ADDR_15_port, B(14) => DATA_ADDR_14_port, B(13)
                           => DATA_ADDR_13_port, B(12) => DATA_ADDR_12_port, 
                           B(11) => DATA_ADDR_11_port, B(10) => 
                           DATA_ADDR_10_port, B(9) => DATA_ADDR_9_port, B(8) =>
                           DATA_ADDR_8_port, B(7) => DATA_ADDR_7_port, B(6) => 
                           DATA_ADDR_6_port, B(5) => DATA_ADDR_5_port, B(4) => 
                           DATA_ADDR_4_port, B(3) => DATA_ADDR_3_port, B(2) => 
                           DATA_ADDR_2_port, B(1) => DATA_ADDR_1_port, B(0) => 
                           DATA_ADDR_0_port, C(31) => WB_in_31_port, C(30) => 
                           WB_in_30_port, C(29) => WB_in_29_port, C(28) => 
                           WB_in_28_port, C(27) => WB_in_27_port, C(26) => 
                           WB_in_26_port, C(25) => WB_in_25_port, C(24) => 
                           WB_in_24_port, C(23) => WB_in_23_port, C(22) => 
                           WB_in_22_port, C(21) => WB_in_21_port, C(20) => 
                           WB_in_20_port, C(19) => WB_in_19_port, C(18) => 
                           WB_in_18_port, C(17) => WB_in_17_port, C(16) => 
                           WB_in_16_port, C(15) => WB_in_15_port, C(14) => 
                           WB_in_14_port, C(13) => WB_in_13_port, C(12) => 
                           WB_in_12_port, C(11) => WB_in_11_port, C(10) => 
                           WB_in_10_port, C(9) => WB_in_9_port, C(8) => 
                           WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => FWDA_SEL_1_port, SEL(0) => 
                           FWDA_SEL_0_port, Y(31) => FWDA_OUT_31_port, Y(30) =>
                           FWDA_OUT_30_port, Y(29) => FWDA_OUT_29_port, Y(28) 
                           => FWDA_OUT_28_port, Y(27) => FWDA_OUT_27_port, 
                           Y(26) => FWDA_OUT_26_port, Y(25) => FWDA_OUT_25_port
                           , Y(24) => FWDA_OUT_24_port, Y(23) => 
                           FWDA_OUT_23_port, Y(22) => FWDA_OUT_22_port, Y(21) 
                           => FWDA_OUT_21_port, Y(20) => FWDA_OUT_20_port, 
                           Y(19) => FWDA_OUT_19_port, Y(18) => FWDA_OUT_18_port
                           , Y(17) => FWDA_OUT_17_port, Y(16) => 
                           FWDA_OUT_16_port, Y(15) => FWDA_OUT_15_port, Y(14) 
                           => FWDA_OUT_14_port, Y(13) => FWDA_OUT_13_port, 
                           Y(12) => FWDA_OUT_12_port, Y(11) => FWDA_OUT_11_port
                           , Y(10) => FWDA_OUT_10_port, Y(9) => FWDA_OUT_9_port
                           , Y(8) => FWDA_OUT_8_port, Y(7) => FWDA_OUT_7_port, 
                           Y(6) => FWDA_OUT_6_port, Y(5) => FWDA_OUT_5_port, 
                           Y(4) => FWDA_OUT_4_port, Y(3) => FWDA_OUT_3_port, 
                           Y(2) => FWDA_OUT_2_port, Y(1) => FWDA_OUT_1_port, 
                           Y(0) => FWDA_OUT_0_port);
   FWDB_MUX : MUX3to1_NBIT32_2 port map( A(31) => RB_out_31_port, A(30) => 
                           RB_out_30_port, A(29) => RB_out_29_port, A(28) => 
                           RB_out_28_port, A(27) => RB_out_27_port, A(26) => 
                           RB_out_26_port, A(25) => RB_out_25_port, A(24) => 
                           RB_out_24_port, A(23) => RB_out_23_port, A(22) => 
                           RB_out_22_port, A(21) => RB_out_21_port, A(20) => 
                           RB_out_20_port, A(19) => RB_out_19_port, A(18) => 
                           RB_out_18_port, A(17) => RB_out_17_port, A(16) => 
                           RB_out_16_port, A(15) => RB_out_15_port, A(14) => 
                           RB_out_14_port, A(13) => RB_out_13_port, A(12) => 
                           RB_out_12_port, A(11) => RB_out_11_port, A(10) => 
                           RB_out_10_port, A(9) => RB_out_9_port, A(8) => 
                           RB_out_8_port, A(7) => RB_out_7_port, A(6) => 
                           RB_out_6_port, A(5) => RB_out_5_port, A(4) => 
                           RB_out_4_port, A(3) => RB_out_3_port, A(2) => 
                           RB_out_2_port, A(1) => RB_out_1_port, A(0) => 
                           RB_out_0_port, B(31) => DATA_ADDR_31_port, B(30) => 
                           DATA_ADDR_30_port, B(29) => DATA_ADDR_29_port, B(28)
                           => DATA_ADDR_28_port, B(27) => DATA_ADDR_27_port, 
                           B(26) => DATA_ADDR_26_port, B(25) => 
                           DATA_ADDR_25_port, B(24) => DATA_ADDR_24_port, B(23)
                           => DATA_ADDR_23_port, B(22) => DATA_ADDR_22_port, 
                           B(21) => DATA_ADDR_21_port, B(20) => 
                           DATA_ADDR_20_port, B(19) => DATA_ADDR_19_port, B(18)
                           => DATA_ADDR_18_port, B(17) => DATA_ADDR_17_port, 
                           B(16) => DATA_ADDR_16_port, B(15) => 
                           DATA_ADDR_15_port, B(14) => DATA_ADDR_14_port, B(13)
                           => DATA_ADDR_13_port, B(12) => DATA_ADDR_12_port, 
                           B(11) => DATA_ADDR_11_port, B(10) => 
                           DATA_ADDR_10_port, B(9) => DATA_ADDR_9_port, B(8) =>
                           DATA_ADDR_8_port, B(7) => DATA_ADDR_7_port, B(6) => 
                           DATA_ADDR_6_port, B(5) => DATA_ADDR_5_port, B(4) => 
                           DATA_ADDR_4_port, B(3) => DATA_ADDR_3_port, B(2) => 
                           DATA_ADDR_2_port, B(1) => DATA_ADDR_1_port, B(0) => 
                           DATA_ADDR_0_port, C(31) => WB_in_31_port, C(30) => 
                           WB_in_30_port, C(29) => WB_in_29_port, C(28) => 
                           WB_in_28_port, C(27) => WB_in_27_port, C(26) => 
                           WB_in_26_port, C(25) => WB_in_25_port, C(24) => 
                           WB_in_24_port, C(23) => WB_in_23_port, C(22) => 
                           WB_in_22_port, C(21) => WB_in_21_port, C(20) => 
                           WB_in_20_port, C(19) => WB_in_19_port, C(18) => 
                           WB_in_18_port, C(17) => WB_in_17_port, C(16) => 
                           WB_in_16_port, C(15) => WB_in_15_port, C(14) => 
                           WB_in_14_port, C(13) => WB_in_13_port, C(12) => 
                           WB_in_12_port, C(11) => WB_in_11_port, C(10) => 
                           WB_in_10_port, C(9) => WB_in_9_port, C(8) => 
                           WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => FWDB_SEL_1_port, SEL(0) => 
                           FWDB_SEL_0_port, Y(31) => FWDB_OUT_31_port, Y(30) =>
                           FWDB_OUT_30_port, Y(29) => FWDB_OUT_29_port, Y(28) 
                           => FWDB_OUT_28_port, Y(27) => FWDB_OUT_27_port, 
                           Y(26) => FWDB_OUT_26_port, Y(25) => FWDB_OUT_25_port
                           , Y(24) => FWDB_OUT_24_port, Y(23) => 
                           FWDB_OUT_23_port, Y(22) => FWDB_OUT_22_port, Y(21) 
                           => FWDB_OUT_21_port, Y(20) => FWDB_OUT_20_port, 
                           Y(19) => FWDB_OUT_19_port, Y(18) => FWDB_OUT_18_port
                           , Y(17) => FWDB_OUT_17_port, Y(16) => 
                           FWDB_OUT_16_port, Y(15) => FWDB_OUT_15_port, Y(14) 
                           => FWDB_OUT_14_port, Y(13) => FWDB_OUT_13_port, 
                           Y(12) => FWDB_OUT_12_port, Y(11) => FWDB_OUT_11_port
                           , Y(10) => FWDB_OUT_10_port, Y(9) => FWDB_OUT_9_port
                           , Y(8) => FWDB_OUT_8_port, Y(7) => FWDB_OUT_7_port, 
                           Y(6) => FWDB_OUT_6_port, Y(5) => FWDB_OUT_5_port, 
                           Y(4) => FWDB_OUT_4_port, Y(3) => FWDB_OUT_3_port, 
                           Y(2) => FWDB_OUT_2_port, Y(1) => FWDB_OUT_1_port, 
                           Y(0) => FWDB_OUT_0_port);
   ZDU_MUX : MUX3to1_NBIT32_1 port map( A(31) => RA_out_31_port, A(30) => 
                           RA_out_30_port, A(29) => RA_out_29_port, A(28) => 
                           RA_out_28_port, A(27) => RA_out_27_port, A(26) => 
                           RA_out_26_port, A(25) => RA_out_25_port, A(24) => 
                           RA_out_24_port, A(23) => RA_out_23_port, A(22) => 
                           RA_out_22_port, A(21) => RA_out_21_port, A(20) => 
                           RA_out_20_port, A(19) => RA_out_19_port, A(18) => 
                           RA_out_18_port, A(17) => RA_out_17_port, A(16) => 
                           RA_out_16_port, A(15) => RA_out_15_port, A(14) => 
                           RA_out_14_port, A(13) => RA_out_13_port, A(12) => 
                           RA_out_12_port, A(11) => RA_out_11_port, A(10) => 
                           RA_out_10_port, A(9) => RA_out_9_port, A(8) => 
                           RA_out_8_port, A(7) => RA_out_7_port, A(6) => 
                           RA_out_6_port, A(5) => RA_out_5_port, A(4) => 
                           RA_out_4_port, A(3) => RA_out_3_port, A(2) => 
                           RA_out_2_port, A(1) => RA_out_1_port, A(0) => 
                           RA_out_0_port, B(31) => CWB_MUX2_out_31_port, B(30) 
                           => CWB_MUX2_out_30_port, B(29) => 
                           CWB_MUX2_out_29_port, B(28) => CWB_MUX2_out_28_port,
                           B(27) => CWB_MUX2_out_27_port, B(26) => 
                           CWB_MUX2_out_26_port, B(25) => CWB_MUX2_out_25_port,
                           B(24) => CWB_MUX2_out_24_port, B(23) => 
                           CWB_MUX2_out_23_port, B(22) => CWB_MUX2_out_22_port,
                           B(21) => CWB_MUX2_out_21_port, B(20) => 
                           CWB_MUX2_out_20_port, B(19) => CWB_MUX2_out_19_port,
                           B(18) => CWB_MUX2_out_18_port, B(17) => 
                           CWB_MUX2_out_17_port, B(16) => CWB_MUX2_out_16_port,
                           B(15) => CWB_MUX2_out_15_port, B(14) => 
                           CWB_MUX2_out_14_port, B(13) => CWB_MUX2_out_13_port,
                           B(12) => CWB_MUX2_out_12_port, B(11) => 
                           CWB_MUX2_out_11_port, B(10) => CWB_MUX2_out_10_port,
                           B(9) => CWB_MUX2_out_9_port, B(8) => 
                           CWB_MUX2_out_8_port, B(7) => CWB_MUX2_out_7_port, 
                           B(6) => CWB_MUX2_out_6_port, B(5) => 
                           CWB_MUX2_out_5_port, B(4) => CWB_MUX2_out_4_port, 
                           B(3) => CWB_MUX2_out_3_port, B(2) => 
                           CWB_MUX2_out_2_port, B(1) => CWB_MUX2_out_1_port, 
                           B(0) => CWB_MUX2_out_0_port, C(31) => WB_in_31_port,
                           C(30) => WB_in_30_port, C(29) => WB_in_29_port, 
                           C(28) => WB_in_28_port, C(27) => WB_in_27_port, 
                           C(26) => WB_in_26_port, C(25) => WB_in_25_port, 
                           C(24) => WB_in_24_port, C(23) => WB_in_23_port, 
                           C(22) => WB_in_22_port, C(21) => WB_in_21_port, 
                           C(20) => WB_in_20_port, C(19) => WB_in_19_port, 
                           C(18) => WB_in_18_port, C(17) => WB_in_17_port, 
                           C(16) => WB_in_16_port, C(15) => WB_in_15_port, 
                           C(14) => WB_in_14_port, C(13) => WB_in_13_port, 
                           C(12) => WB_in_12_port, C(11) => WB_in_11_port, 
                           C(10) => WB_in_10_port, C(9) => WB_in_9_port, C(8) 
                           => WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => ZDU_SEL_1_port, SEL(0) => 
                           ZDU_SEL_0_port, Y(31) => n_1608, Y(30) => 
                           ZDU_MUX_out_30_port, Y(29) => ZDU_MUX_out_29_port, 
                           Y(28) => ZDU_MUX_out_28_port, Y(27) => 
                           ZDU_MUX_out_27_port, Y(26) => ZDU_MUX_out_26_port, 
                           Y(25) => ZDU_MUX_out_25_port, Y(24) => 
                           ZDU_MUX_out_24_port, Y(23) => ZDU_MUX_out_23_port, 
                           Y(22) => ZDU_MUX_out_22_port, Y(21) => 
                           ZDU_MUX_out_21_port, Y(20) => ZDU_MUX_out_20_port, 
                           Y(19) => ZDU_MUX_out_19_port, Y(18) => 
                           ZDU_MUX_out_18_port, Y(17) => ZDU_MUX_out_17_port, 
                           Y(16) => ZDU_MUX_out_16_port, Y(15) => 
                           ZDU_MUX_out_15_port, Y(14) => ZDU_MUX_out_14_port, 
                           Y(13) => ZDU_MUX_out_13_port, Y(12) => 
                           ZDU_MUX_out_12_port, Y(11) => ZDU_MUX_out_11_port, 
                           Y(10) => ZDU_MUX_out_10_port, Y(9) => 
                           ZDU_MUX_out_9_port, Y(8) => ZDU_MUX_out_8_port, Y(7)
                           => ZDU_MUX_out_7_port, Y(6) => ZDU_MUX_out_6_port, 
                           Y(5) => ZDU_MUX_out_5_port, Y(4) => 
                           ZDU_MUX_out_4_port, Y(3) => ZDU_MUX_out_3_port, Y(2)
                           => ZDU_MUX_out_2_port, Y(1) => ZDU_MUX_out_1_port, 
                           Y(0) => ZDU_MUX_out_0_port);
   MEMDATAMUX : MUX2to1_NBIT32_4 port map( A(31) => ALR2_out_31_port, A(30) => 
                           ALR2_out_30_port, A(29) => ALR2_out_29_port, A(28) 
                           => ALR2_out_28_port, A(27) => ALR2_out_27_port, 
                           A(26) => ALR2_out_26_port, A(25) => ALR2_out_25_port
                           , A(24) => ALR2_out_24_port, A(23) => 
                           ALR2_out_23_port, A(22) => ALR2_out_22_port, A(21) 
                           => ALR2_out_21_port, A(20) => ALR2_out_20_port, 
                           A(19) => ALR2_out_19_port, A(18) => ALR2_out_18_port
                           , A(17) => ALR2_out_17_port, A(16) => 
                           ALR2_out_16_port, A(15) => ALR2_out_15_port, A(14) 
                           => ALR2_out_14_port, A(13) => ALR2_out_13_port, 
                           A(12) => ALR2_out_12_port, A(11) => ALR2_out_11_port
                           , A(10) => ALR2_out_10_port, A(9) => ALR2_out_9_port
                           , A(8) => ALR2_out_8_port, A(7) => ALR2_out_7_port, 
                           A(6) => ALR2_out_6_port, A(5) => ALR2_out_5_port, 
                           A(4) => ALR2_out_4_port, A(3) => ALR2_out_3_port, 
                           A(2) => ALR2_out_2_port, A(1) => ALR2_out_1_port, 
                           A(0) => ALR2_out_0_port, B(31) => B2_MUX_out_31_port
                           , B(30) => B2_MUX_out_30_port, B(29) => 
                           B2_MUX_out_29_port, B(28) => B2_MUX_out_28_port, 
                           B(27) => B2_MUX_out_27_port, B(26) => 
                           B2_MUX_out_26_port, B(25) => B2_MUX_out_25_port, 
                           B(24) => B2_MUX_out_24_port, B(23) => 
                           B2_MUX_out_23_port, B(22) => B2_MUX_out_22_port, 
                           B(21) => B2_MUX_out_21_port, B(20) => 
                           B2_MUX_out_20_port, B(19) => B2_MUX_out_19_port, 
                           B(18) => B2_MUX_out_18_port, B(17) => 
                           B2_MUX_out_17_port, B(16) => B2_MUX_out_16_port, 
                           B(15) => B2_MUX_out_15_port, B(14) => 
                           B2_MUX_out_14_port, B(13) => B2_MUX_out_13_port, 
                           B(12) => B2_MUX_out_12_port, B(11) => 
                           B2_MUX_out_11_port, B(10) => B2_MUX_out_10_port, 
                           B(9) => B2_MUX_out_9_port, B(8) => B2_MUX_out_8_port
                           , B(7) => B2_MUX_out_7_port, B(6) => 
                           B2_MUX_out_6_port, B(5) => B2_MUX_out_5_port, B(4) 
                           => B2_MUX_out_4_port, B(3) => B2_MUX_out_3_port, 
                           B(2) => B2_MUX_out_2_port, B(1) => B2_MUX_out_1_port
                           , B(0) => B2_MUX_out_0_port, SEL => MEM_DATA_SEL, 
                           Y(31) => DATA_OUT(31), Y(30) => DATA_OUT(30), Y(29) 
                           => DATA_OUT(29), Y(28) => DATA_OUT(28), Y(27) => 
                           DATA_OUT(27), Y(26) => DATA_OUT(26), Y(25) => 
                           DATA_OUT(25), Y(24) => DATA_OUT(24), Y(23) => 
                           DATA_OUT(23), Y(22) => DATA_OUT(22), Y(21) => 
                           DATA_OUT(21), Y(20) => DATA_OUT(20), Y(19) => 
                           DATA_OUT(19), Y(18) => DATA_OUT(18), Y(17) => 
                           DATA_OUT(17), Y(16) => DATA_OUT(16), Y(15) => 
                           DATA_OUT(15), Y(14) => DATA_OUT(14), Y(13) => 
                           DATA_OUT(13), Y(12) => DATA_OUT(12), Y(11) => 
                           DATA_OUT(11), Y(10) => DATA_OUT(10), Y(9) => 
                           DATA_OUT(9), Y(8) => DATA_OUT(8), Y(7) => 
                           DATA_OUT(7), Y(6) => DATA_OUT(6), Y(5) => 
                           DATA_OUT(5), Y(4) => DATA_OUT(4), Y(3) => 
                           DATA_OUT(3), Y(2) => DATA_OUT(2), Y(1) => 
                           DATA_OUT(1), Y(0) => DATA_OUT(0));
   LMDMUX : MUX5to1_NBIT32_0 port map( A(31) => n43, A(30) => DATA_IN(6), A(29)
                           => DATA_IN(5), A(28) => DATA_IN(4), A(27) => 
                           DATA_IN(3), A(26) => DATA_IN(2), A(25) => DATA_IN(1)
                           , A(24) => DATA_IN(0), A(23) => DATA_IN(15), A(22) 
                           => DATA_IN(14), A(21) => DATA_IN(13), A(20) => 
                           DATA_IN(12), A(19) => DATA_IN(11), A(18) => 
                           DATA_IN(10), A(17) => DATA_IN(9), A(16) => 
                           DATA_IN(8), A(15) => DATA_IN(23), A(14) => 
                           DATA_IN(22), A(13) => DATA_IN(21), A(12) => 
                           DATA_IN(20), A(11) => DATA_IN(19), A(10) => 
                           DATA_IN(18), A(9) => DATA_IN(17), A(8) => 
                           DATA_IN(16), A(7) => DATA_IN(31), A(6) => 
                           DATA_IN(30), A(5) => DATA_IN(29), A(4) => 
                           DATA_IN(28), A(3) => DATA_IN(27), A(2) => 
                           DATA_IN(26), A(1) => DATA_IN(25), A(0) => 
                           DATA_IN(24), B(31) => n44, B(30) => n44, B(29) => 
                           n44, B(28) => n45, B(27) => n45, B(26) => n45, B(25)
                           => n45, B(24) => n45, B(23) => n45, B(22) => n45, 
                           B(21) => n45, B(20) => n45, B(19) => n45, B(18) => 
                           n45, B(17) => n45, B(16) => n45, B(15) => n46, B(14)
                           => n46, B(13) => n46, B(12) => n46, B(11) => n46, 
                           B(10) => n46, B(9) => n46, B(8) => n46, B(7) => n44,
                           B(6) => DATA_IN(6), B(5) => DATA_IN(5), B(4) => 
                           DATA_IN(4), B(3) => DATA_IN(3), B(2) => DATA_IN(2), 
                           B(1) => DATA_IN(1), B(0) => DATA_IN(0), C(31) => 
                           X_Logic0_port, C(30) => X_Logic0_port, C(29) => 
                           X_Logic0_port, C(28) => X_Logic0_port, C(27) => 
                           X_Logic0_port, C(26) => X_Logic0_port, C(25) => 
                           X_Logic0_port, C(24) => X_Logic0_port, C(23) => 
                           X_Logic0_port, C(22) => X_Logic0_port, C(21) => 
                           X_Logic0_port, C(20) => X_Logic0_port, C(19) => 
                           X_Logic0_port, C(18) => X_Logic0_port, C(17) => 
                           X_Logic0_port, C(16) => X_Logic0_port, C(15) => 
                           X_Logic0_port, C(14) => X_Logic0_port, C(13) => 
                           X_Logic0_port, C(12) => X_Logic0_port, C(11) => 
                           X_Logic0_port, C(10) => X_Logic0_port, C(9) => 
                           X_Logic0_port, C(8) => X_Logic0_port, C(7) => n44, 
                           C(6) => DATA_IN(6), C(5) => DATA_IN(5), C(4) => 
                           DATA_IN(4), C(3) => DATA_IN(3), C(2) => DATA_IN(2), 
                           C(1) => DATA_IN(1), C(0) => DATA_IN(0), D(31) => n44
                           , D(30) => n44, D(29) => n44, D(28) => n44, D(27) =>
                           n44, D(26) => n43, D(25) => n44, D(24) => n43, D(23)
                           => n43, D(22) => n43, D(21) => n43, D(20) => n43, 
                           D(19) => n43, D(18) => n43, D(17) => n43, D(16) => 
                           n43, D(15) => n43, D(14) => DATA_IN(6), D(13) => 
                           DATA_IN(5), D(12) => DATA_IN(4), D(11) => DATA_IN(3)
                           , D(10) => DATA_IN(2), D(9) => DATA_IN(1), D(8) => 
                           DATA_IN(0), D(7) => DATA_IN(15), D(6) => DATA_IN(14)
                           , D(5) => DATA_IN(13), D(4) => DATA_IN(12), D(3) => 
                           DATA_IN(11), D(2) => DATA_IN(10), D(1) => DATA_IN(9)
                           , D(0) => DATA_IN(8), E(31) => X_Logic0_port, E(30) 
                           => X_Logic0_port, E(29) => X_Logic0_port, E(28) => 
                           X_Logic0_port, E(27) => X_Logic0_port, E(26) => 
                           X_Logic0_port, E(25) => X_Logic0_port, E(24) => 
                           X_Logic0_port, E(23) => X_Logic0_port, E(22) => 
                           X_Logic0_port, E(21) => X_Logic0_port, E(20) => 
                           X_Logic0_port, E(19) => X_Logic0_port, E(18) => 
                           X_Logic0_port, E(17) => X_Logic0_port, E(16) => 
                           X_Logic0_port, E(15) => n44, E(14) => DATA_IN(6), 
                           E(13) => DATA_IN(5), E(12) => DATA_IN(4), E(11) => 
                           DATA_IN(3), E(10) => DATA_IN(2), E(9) => DATA_IN(1),
                           E(8) => DATA_IN(0), E(7) => DATA_IN(15), E(6) => 
                           DATA_IN(14), E(5) => DATA_IN(13), E(4) => 
                           DATA_IN(12), E(3) => DATA_IN(11), E(2) => 
                           DATA_IN(10), E(1) => DATA_IN(9), E(0) => DATA_IN(8),
                           SEL(2) => LD_SEL(2), SEL(1) => LD_SEL(1), SEL(0) => 
                           LD_SEL(0), Y(31) => LMD_out_31_port, Y(30) => 
                           LMD_out_30_port, Y(29) => LMD_out_29_port, Y(28) => 
                           LMD_out_28_port, Y(27) => LMD_out_27_port, Y(26) => 
                           LMD_out_26_port, Y(25) => LMD_out_25_port, Y(24) => 
                           LMD_out_24_port, Y(23) => LMD_out_23_port, Y(22) => 
                           LMD_out_22_port, Y(21) => LMD_out_21_port, Y(20) => 
                           LMD_out_20_port, Y(19) => LMD_out_19_port, Y(18) => 
                           LMD_out_18_port, Y(17) => LMD_out_17_port, Y(16) => 
                           LMD_out_16_port, Y(15) => LMD_out_15_port, Y(14) => 
                           LMD_out_14_port, Y(13) => LMD_out_13_port, Y(12) => 
                           LMD_out_12_port, Y(11) => LMD_out_11_port, Y(10) => 
                           LMD_out_10_port, Y(9) => LMD_out_9_port, Y(8) => 
                           LMD_out_8_port, Y(7) => LMD_out_7_port, Y(6) => 
                           LMD_out_6_port, Y(5) => LMD_out_5_port, Y(4) => 
                           LMD_out_4_port, Y(3) => LMD_out_3_port, Y(2) => 
                           LMD_out_2_port, Y(1) => LMD_out_1_port, Y(0) => 
                           LMD_out_0_port);
   ALR2_MUX : MUX2to1_NBIT32_3 port map( A(31) => CWB_MUX2_out_31_port, A(30) 
                           => CWB_MUX2_out_30_port, A(29) => 
                           CWB_MUX2_out_29_port, A(28) => CWB_MUX2_out_28_port,
                           A(27) => CWB_MUX2_out_27_port, A(26) => 
                           CWB_MUX2_out_26_port, A(25) => CWB_MUX2_out_25_port,
                           A(24) => CWB_MUX2_out_24_port, A(23) => 
                           CWB_MUX2_out_23_port, A(22) => CWB_MUX2_out_22_port,
                           A(21) => CWB_MUX2_out_21_port, A(20) => 
                           CWB_MUX2_out_20_port, A(19) => CWB_MUX2_out_19_port,
                           A(18) => CWB_MUX2_out_18_port, A(17) => 
                           CWB_MUX2_out_17_port, A(16) => CWB_MUX2_out_16_port,
                           A(15) => CWB_MUX2_out_15_port, A(14) => 
                           CWB_MUX2_out_14_port, A(13) => CWB_MUX2_out_13_port,
                           A(12) => CWB_MUX2_out_12_port, A(11) => 
                           CWB_MUX2_out_11_port, A(10) => CWB_MUX2_out_10_port,
                           A(9) => CWB_MUX2_out_9_port, A(8) => 
                           CWB_MUX2_out_8_port, A(7) => CWB_MUX2_out_7_port, 
                           A(6) => CWB_MUX2_out_6_port, A(5) => 
                           CWB_MUX2_out_5_port, A(4) => CWB_MUX2_out_4_port, 
                           A(3) => CWB_MUX2_out_3_port, A(2) => 
                           CWB_MUX2_out_2_port, A(1) => CWB_MUX2_out_1_port, 
                           A(0) => CWB_MUX2_out_0_port, B(31) => 
                           NPC3_out_31_port, B(30) => NPC3_out_30_port, B(29) 
                           => NPC3_out_29_port, B(28) => NPC3_out_28_port, 
                           B(27) => NPC3_out_27_port, B(26) => NPC3_out_26_port
                           , B(25) => NPC3_out_25_port, B(24) => 
                           NPC3_out_24_port, B(23) => NPC3_out_23_port, B(22) 
                           => NPC3_out_22_port, B(21) => NPC3_out_21_port, 
                           B(20) => NPC3_out_20_port, B(19) => NPC3_out_19_port
                           , B(18) => NPC3_out_18_port, B(17) => 
                           NPC3_out_17_port, B(16) => NPC3_out_16_port, B(15) 
                           => NPC3_out_15_port, B(14) => NPC3_out_14_port, 
                           B(13) => NPC3_out_13_port, B(12) => NPC3_out_12_port
                           , B(11) => NPC3_out_11_port, B(10) => 
                           NPC3_out_10_port, B(9) => NPC3_out_9_port, B(8) => 
                           NPC3_out_8_port, B(7) => NPC3_out_7_port, B(6) => 
                           NPC3_out_6_port, B(5) => NPC3_out_5_port, B(4) => 
                           NPC3_out_4_port, B(3) => NPC3_out_3_port, B(2) => 
                           NPC3_out_2_port, B(1) => NPC3_out_1_port, B(0) => 
                           NPC3_out_0_port, SEL => ALR2_SEL, Y(31) => 
                           ALR2_in_31_port, Y(30) => ALR2_in_30_port, Y(29) => 
                           ALR2_in_29_port, Y(28) => ALR2_in_28_port, Y(27) => 
                           ALR2_in_27_port, Y(26) => ALR2_in_26_port, Y(25) => 
                           ALR2_in_25_port, Y(24) => ALR2_in_24_port, Y(23) => 
                           ALR2_in_23_port, Y(22) => ALR2_in_22_port, Y(21) => 
                           ALR2_in_21_port, Y(20) => ALR2_in_20_port, Y(19) => 
                           ALR2_in_19_port, Y(18) => ALR2_in_18_port, Y(17) => 
                           ALR2_in_17_port, Y(16) => ALR2_in_16_port, Y(15) => 
                           ALR2_in_15_port, Y(14) => ALR2_in_14_port, Y(13) => 
                           ALR2_in_13_port, Y(12) => ALR2_in_12_port, Y(11) => 
                           ALR2_in_11_port, Y(10) => ALR2_in_10_port, Y(9) => 
                           ALR2_in_9_port, Y(8) => ALR2_in_8_port, Y(7) => 
                           ALR2_in_7_port, Y(6) => ALR2_in_6_port, Y(5) => 
                           ALR2_in_5_port, Y(4) => ALR2_in_4_port, Y(3) => 
                           ALR2_in_3_port, Y(2) => ALR2_in_2_port, Y(1) => 
                           ALR2_in_1_port, Y(0) => ALR2_in_0_port);
   CWB_MUX1 : MUX3to1_NBIT2 port map( A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, C(1) => CWB_out_1_port, C(0) => 
                           CWB_out_0_port, SEL(1) => CWB_MUX_SEL_1_port, SEL(0)
                           => CWB_MUX_SEL_0_port, Y(1) => CWB2_SEL_1_port, Y(0)
                           => CWB2_SEL_0_port);
   CWB_MUX2 : MUX4to1_NBIT32_0 port map( A(31) => DATA_ADDR_31_port, A(30) => 
                           DATA_ADDR_30_port, A(29) => DATA_ADDR_29_port, A(28)
                           => DATA_ADDR_28_port, A(27) => DATA_ADDR_27_port, 
                           A(26) => DATA_ADDR_26_port, A(25) => 
                           DATA_ADDR_25_port, A(24) => DATA_ADDR_24_port, A(23)
                           => DATA_ADDR_23_port, A(22) => DATA_ADDR_22_port, 
                           A(21) => DATA_ADDR_21_port, A(20) => 
                           DATA_ADDR_20_port, A(19) => DATA_ADDR_19_port, A(18)
                           => DATA_ADDR_18_port, A(17) => DATA_ADDR_17_port, 
                           A(16) => DATA_ADDR_16_port, A(15) => 
                           DATA_ADDR_15_port, A(14) => DATA_ADDR_14_port, A(13)
                           => DATA_ADDR_13_port, A(12) => DATA_ADDR_12_port, 
                           A(11) => DATA_ADDR_11_port, A(10) => 
                           DATA_ADDR_10_port, A(9) => DATA_ADDR_9_port, A(8) =>
                           DATA_ADDR_8_port, A(7) => DATA_ADDR_7_port, A(6) => 
                           DATA_ADDR_6_port, A(5) => DATA_ADDR_5_port, A(4) => 
                           DATA_ADDR_4_port, A(3) => DATA_ADDR_3_port, A(2) => 
                           DATA_ADDR_2_port, A(1) => DATA_ADDR_1_port, A(0) => 
                           DATA_ADDR_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, C(31) => X_Logic0_port, C(30) => 
                           X_Logic0_port, C(29) => X_Logic0_port, C(28) => 
                           X_Logic0_port, C(27) => X_Logic0_port, C(26) => 
                           X_Logic0_port, C(25) => X_Logic0_port, C(24) => 
                           X_Logic0_port, C(23) => X_Logic0_port, C(22) => 
                           X_Logic0_port, C(21) => X_Logic0_port, C(20) => 
                           X_Logic0_port, C(19) => X_Logic0_port, C(18) => 
                           X_Logic0_port, C(17) => X_Logic0_port, C(16) => 
                           X_Logic0_port, C(15) => X_Logic0_port, C(14) => 
                           X_Logic0_port, C(13) => X_Logic0_port, C(12) => 
                           X_Logic0_port, C(11) => X_Logic0_port, C(10) => 
                           X_Logic0_port, C(9) => X_Logic0_port, C(8) => 
                           X_Logic0_port, C(7) => X_Logic0_port, C(6) => 
                           X_Logic0_port, C(5) => X_Logic0_port, C(4) => 
                           X_Logic0_port, C(3) => X_Logic0_port, C(2) => 
                           X_Logic0_port, C(1) => X_Logic0_port, C(0) => 
                           X_Logic0_port, D(31) => DATA_ADDR_15_port, D(30) => 
                           DATA_ADDR_14_port, D(29) => DATA_ADDR_13_port, D(28)
                           => DATA_ADDR_12_port, D(27) => DATA_ADDR_11_port, 
                           D(26) => DATA_ADDR_10_port, D(25) => 
                           DATA_ADDR_9_port, D(24) => DATA_ADDR_8_port, D(23) 
                           => DATA_ADDR_7_port, D(22) => DATA_ADDR_6_port, 
                           D(21) => DATA_ADDR_5_port, D(20) => DATA_ADDR_4_port
                           , D(19) => DATA_ADDR_3_port, D(18) => 
                           DATA_ADDR_2_port, D(17) => DATA_ADDR_1_port, D(16) 
                           => DATA_ADDR_0_port, D(15) => X_Logic0_port, D(14) 
                           => X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, SEL(1) => CWB2_SEL_1_port, SEL(0) => 
                           CWB2_SEL_0_port, Y(31) => CWB_MUX2_out_31_port, 
                           Y(30) => CWB_MUX2_out_30_port, Y(29) => 
                           CWB_MUX2_out_29_port, Y(28) => CWB_MUX2_out_28_port,
                           Y(27) => CWB_MUX2_out_27_port, Y(26) => 
                           CWB_MUX2_out_26_port, Y(25) => CWB_MUX2_out_25_port,
                           Y(24) => CWB_MUX2_out_24_port, Y(23) => 
                           CWB_MUX2_out_23_port, Y(22) => CWB_MUX2_out_22_port,
                           Y(21) => CWB_MUX2_out_21_port, Y(20) => 
                           CWB_MUX2_out_20_port, Y(19) => CWB_MUX2_out_19_port,
                           Y(18) => CWB_MUX2_out_18_port, Y(17) => 
                           CWB_MUX2_out_17_port, Y(16) => CWB_MUX2_out_16_port,
                           Y(15) => CWB_MUX2_out_15_port, Y(14) => 
                           CWB_MUX2_out_14_port, Y(13) => CWB_MUX2_out_13_port,
                           Y(12) => CWB_MUX2_out_12_port, Y(11) => 
                           CWB_MUX2_out_11_port, Y(10) => CWB_MUX2_out_10_port,
                           Y(9) => CWB_MUX2_out_9_port, Y(8) => 
                           CWB_MUX2_out_8_port, Y(7) => CWB_MUX2_out_7_port, 
                           Y(6) => CWB_MUX2_out_6_port, Y(5) => 
                           CWB_MUX2_out_5_port, Y(4) => CWB_MUX2_out_4_port, 
                           Y(3) => CWB_MUX2_out_3_port, Y(2) => 
                           CWB_MUX2_out_2_port, Y(1) => CWB_MUX2_out_1_port, 
                           Y(0) => CWB_MUX2_out_0_port);
   B2_MUX : MUX2to1_NBIT32_2 port map( A(31) => B2_out_31_port, A(30) => 
                           B2_out_30_port, A(29) => B2_out_29_port, A(28) => 
                           B2_out_28_port, A(27) => B2_out_27_port, A(26) => 
                           B2_out_26_port, A(25) => B2_out_25_port, A(24) => 
                           B2_out_24_port, A(23) => B2_out_23_port, A(22) => 
                           B2_out_22_port, A(21) => B2_out_21_port, A(20) => 
                           B2_out_20_port, A(19) => B2_out_19_port, A(18) => 
                           B2_out_18_port, A(17) => B2_out_17_port, A(16) => 
                           B2_out_16_port, A(15) => B2_out_15_port, A(14) => 
                           B2_out_14_port, A(13) => B2_out_13_port, A(12) => 
                           B2_out_12_port, A(11) => B2_out_11_port, A(10) => 
                           B2_out_10_port, A(9) => B2_out_9_port, A(8) => 
                           B2_out_8_port, A(7) => B2_out_7_port, A(6) => 
                           B2_out_6_port, A(5) => B2_out_5_port, A(4) => 
                           B2_out_4_port, A(3) => B2_out_3_port, A(2) => 
                           B2_out_2_port, A(1) => B2_out_1_port, A(0) => 
                           B2_out_0_port, B(31) => WB_in_31_port, B(30) => 
                           WB_in_30_port, B(29) => WB_in_29_port, B(28) => 
                           WB_in_28_port, B(27) => WB_in_27_port, B(26) => 
                           WB_in_26_port, B(25) => WB_in_25_port, B(24) => 
                           WB_in_24_port, B(23) => WB_in_23_port, B(22) => 
                           WB_in_22_port, B(21) => WB_in_21_port, B(20) => 
                           WB_in_20_port, B(19) => WB_in_19_port, B(18) => 
                           WB_in_18_port, B(17) => WB_in_17_port, B(16) => 
                           WB_in_16_port, B(15) => WB_in_15_port, B(14) => 
                           WB_in_14_port, B(13) => WB_in_13_port, B(12) => 
                           WB_in_12_port, B(11) => WB_in_11_port, B(10) => 
                           WB_in_10_port, B(9) => WB_in_9_port, B(8) => 
                           WB_in_8_port, B(7) => WB_in_7_port, B(6) => 
                           WB_in_6_port, B(5) => WB_in_5_port, B(4) => 
                           WB_in_4_port, B(3) => WB_in_3_port, B(2) => 
                           WB_in_2_port, B(1) => WB_in_1_port, B(0) => 
                           WB_in_0_port, SEL => FWDB2_SEL, Y(31) => 
                           B2_MUX_out_31_port, Y(30) => B2_MUX_out_30_port, 
                           Y(29) => B2_MUX_out_29_port, Y(28) => 
                           B2_MUX_out_28_port, Y(27) => B2_MUX_out_27_port, 
                           Y(26) => B2_MUX_out_26_port, Y(25) => 
                           B2_MUX_out_25_port, Y(24) => B2_MUX_out_24_port, 
                           Y(23) => B2_MUX_out_23_port, Y(22) => 
                           B2_MUX_out_22_port, Y(21) => B2_MUX_out_21_port, 
                           Y(20) => B2_MUX_out_20_port, Y(19) => 
                           B2_MUX_out_19_port, Y(18) => B2_MUX_out_18_port, 
                           Y(17) => B2_MUX_out_17_port, Y(16) => 
                           B2_MUX_out_16_port, Y(15) => B2_MUX_out_15_port, 
                           Y(14) => B2_MUX_out_14_port, Y(13) => 
                           B2_MUX_out_13_port, Y(12) => B2_MUX_out_12_port, 
                           Y(11) => B2_MUX_out_11_port, Y(10) => 
                           B2_MUX_out_10_port, Y(9) => B2_MUX_out_9_port, Y(8) 
                           => B2_MUX_out_8_port, Y(7) => B2_MUX_out_7_port, 
                           Y(6) => B2_MUX_out_6_port, Y(5) => B2_MUX_out_5_port
                           , Y(4) => B2_MUX_out_4_port, Y(3) => 
                           B2_MUX_out_3_port, Y(2) => B2_MUX_out_2_port, Y(1) 
                           => B2_MUX_out_1_port, Y(0) => B2_MUX_out_0_port);
   WBMUX : MUX2to1_NBIT32_1 port map( A(31) => ALR2_out_31_port, A(30) => 
                           ALR2_out_30_port, A(29) => ALR2_out_29_port, A(28) 
                           => ALR2_out_28_port, A(27) => ALR2_out_27_port, 
                           A(26) => ALR2_out_26_port, A(25) => ALR2_out_25_port
                           , A(24) => ALR2_out_24_port, A(23) => 
                           ALR2_out_23_port, A(22) => ALR2_out_22_port, A(21) 
                           => ALR2_out_21_port, A(20) => ALR2_out_20_port, 
                           A(19) => ALR2_out_19_port, A(18) => ALR2_out_18_port
                           , A(17) => ALR2_out_17_port, A(16) => 
                           ALR2_out_16_port, A(15) => ALR2_out_15_port, A(14) 
                           => ALR2_out_14_port, A(13) => ALR2_out_13_port, 
                           A(12) => ALR2_out_12_port, A(11) => ALR2_out_11_port
                           , A(10) => ALR2_out_10_port, A(9) => ALR2_out_9_port
                           , A(8) => ALR2_out_8_port, A(7) => ALR2_out_7_port, 
                           A(6) => ALR2_out_6_port, A(5) => ALR2_out_5_port, 
                           A(4) => ALR2_out_4_port, A(3) => ALR2_out_3_port, 
                           A(2) => ALR2_out_2_port, A(1) => ALR2_out_1_port, 
                           A(0) => ALR2_out_0_port, B(31) => LMD_out_31_port, 
                           B(30) => LMD_out_30_port, B(29) => LMD_out_29_port, 
                           B(28) => LMD_out_28_port, B(27) => LMD_out_27_port, 
                           B(26) => LMD_out_26_port, B(25) => LMD_out_25_port, 
                           B(24) => LMD_out_24_port, B(23) => LMD_out_23_port, 
                           B(22) => LMD_out_22_port, B(21) => LMD_out_21_port, 
                           B(20) => LMD_out_20_port, B(19) => LMD_out_19_port, 
                           B(18) => LMD_out_18_port, B(17) => LMD_out_17_port, 
                           B(16) => LMD_out_16_port, B(15) => LMD_out_15_port, 
                           B(14) => LMD_out_14_port, B(13) => LMD_out_13_port, 
                           B(12) => LMD_out_12_port, B(11) => LMD_out_11_port, 
                           B(10) => LMD_out_10_port, B(9) => LMD_out_9_port, 
                           B(8) => LMD_out_8_port, B(7) => LMD_out_7_port, B(6)
                           => LMD_out_6_port, B(5) => LMD_out_5_port, B(4) => 
                           LMD_out_4_port, B(3) => LMD_out_3_port, B(2) => 
                           LMD_out_2_port, B(1) => LMD_out_1_port, B(0) => 
                           LMD_out_0_port, SEL => WB_SEL, Y(31) => 
                           WB_in_31_port, Y(30) => WB_in_30_port, Y(29) => 
                           WB_in_29_port, Y(28) => WB_in_28_port, Y(27) => 
                           WB_in_27_port, Y(26) => WB_in_26_port, Y(25) => 
                           WB_in_25_port, Y(24) => WB_in_24_port, Y(23) => 
                           WB_in_23_port, Y(22) => WB_in_22_port, Y(21) => 
                           WB_in_21_port, Y(20) => WB_in_20_port, Y(19) => 
                           WB_in_19_port, Y(18) => WB_in_18_port, Y(17) => 
                           WB_in_17_port, Y(16) => WB_in_16_port, Y(15) => 
                           WB_in_15_port, Y(14) => WB_in_14_port, Y(13) => 
                           WB_in_13_port, Y(12) => WB_in_12_port, Y(11) => 
                           WB_in_11_port, Y(10) => WB_in_10_port, Y(9) => 
                           WB_in_9_port, Y(8) => WB_in_8_port, Y(7) => 
                           WB_in_7_port, Y(6) => WB_in_6_port, Y(5) => 
                           WB_in_5_port, Y(4) => WB_in_4_port, Y(3) => 
                           WB_in_3_port, Y(2) => WB_in_2_port, Y(1) => 
                           WB_in_1_port, Y(0) => WB_in_0_port);
   RF_MUX_ADDR : MUX3to1_NBIT5 port map( A(4) => RWB3_out_15_port, A(3) => 
                           RWB3_out_14_port, A(2) => RWB3_out_13_port, A(1) => 
                           RWB3_out_12_port, A(0) => RWB3_out_11_port, B(4) => 
                           RWB3_out_20_port, B(3) => RWB3_out_19_port, B(2) => 
                           RWB3_out_18_port, B(1) => RWB3_out_17_port, B(0) => 
                           RWB3_out_16_port, C(4) => X_Logic1_port, C(3) => 
                           X_Logic1_port, C(2) => X_Logic1_port, C(1) => 
                           X_Logic1_port, C(0) => X_Logic1_port, SEL(1) => 
                           RF_MUX_SEL(1), SEL(0) => RF_MUX_SEL(0), Y(4) => 
                           RF_MUX_out_4_port, Y(3) => RF_MUX_out_3_port, Y(2) 
                           => RF_MUX_out_2_port, Y(1) => RF_MUX_out_1_port, 
                           Y(0) => RF_MUX_out_0_port);
   ALU1 : ALU_NBIT32 port map( CLOCK => CLK, AluOpcode(0) => ALU_OPCODE(0), 
                           AluOpcode(1) => ALU_OPCODE(1), AluOpcode(2) => 
                           ALU_OPCODE(2), AluOpcode(3) => ALU_OPCODE(3), 
                           AluOpcode(4) => ALU_OPCODE(4), A(31) => A_in_31_port
                           , A(30) => A_in_30_port, A(29) => A_in_29_port, 
                           A(28) => A_in_28_port, A(27) => A_in_27_port, A(26) 
                           => A_in_26_port, A(25) => A_in_25_port, A(24) => 
                           A_in_24_port, A(23) => A_in_23_port, A(22) => 
                           A_in_22_port, A(21) => A_in_21_port, A(20) => 
                           A_in_20_port, A(19) => A_in_19_port, A(18) => 
                           A_in_18_port, A(17) => A_in_17_port, A(16) => 
                           A_in_16_port, A(15) => A_in_15_port, A(14) => 
                           A_in_14_port, A(13) => A_in_13_port, A(12) => 
                           A_in_12_port, A(11) => A_in_11_port, A(10) => 
                           A_in_10_port, A(9) => A_in_9_port, A(8) => 
                           A_in_8_port, A(7) => A_in_7_port, A(6) => 
                           A_in_6_port, A(5) => A_in_5_port, A(4) => 
                           A_in_4_port, A(3) => A_in_3_port, A(2) => 
                           A_in_2_port, A(1) => A_in_1_port, A(0) => 
                           A_in_0_port, B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Cin => PSW_out_6_port, ALU_out(31) => 
                           ALR_in_31_port, ALU_out(30) => ALR_in_30_port, 
                           ALU_out(29) => ALR_in_29_port, ALU_out(28) => 
                           ALR_in_28_port, ALU_out(27) => ALR_in_27_port, 
                           ALU_out(26) => ALR_in_26_port, ALU_out(25) => 
                           ALR_in_25_port, ALU_out(24) => ALR_in_24_port, 
                           ALU_out(23) => ALR_in_23_port, ALU_out(22) => 
                           ALR_in_22_port, ALU_out(21) => ALR_in_21_port, 
                           ALU_out(20) => ALR_in_20_port, ALU_out(19) => 
                           ALR_in_19_port, ALU_out(18) => ALR_in_18_port, 
                           ALU_out(17) => ALR_in_17_port, ALU_out(16) => 
                           ALR_in_16_port, ALU_out(15) => ALR_in_15_port, 
                           ALU_out(14) => ALR_in_14_port, ALU_out(13) => 
                           ALR_in_13_port, ALU_out(12) => ALR_in_12_port, 
                           ALU_out(11) => ALR_in_11_port, ALU_out(10) => 
                           ALR_in_10_port, ALU_out(9) => ALR_in_9_port, 
                           ALU_out(8) => ALR_in_8_port, ALU_out(7) => 
                           ALR_in_7_port, ALU_out(6) => ALR_in_6_port, 
                           ALU_out(5) => ALR_in_5_port, ALU_out(4) => 
                           ALR_in_4_port, ALU_out(3) => ALR_in_3_port, 
                           ALU_out(2) => ALR_in_2_port, ALU_out(1) => 
                           ALR_in_1_port, ALU_out(0) => ALR_in_0_port, Cout => 
                           PSW_in_6_port, COND(5) => PSW_in_5_port, COND(4) => 
                           PSW_in_4_port, COND(3) => PSW_in_3_port, COND(2) => 
                           PSW_in_2_port, COND(1) => PSW_in_1_port, COND(0) => 
                           PSW_in_0_port);
   FWD1 : FWDU_IR_SIZE32 port map( CLOCK => CLK, RESET => n51, EN => n38, 
                           IR(31) => IR_out_31_port, IR(30) => IR_out_30_port, 
                           IR(29) => IR_out_29_port, IR(28) => IR_out_28_port, 
                           IR(27) => IR_out_27_port, IR(26) => IR_out_26_port, 
                           IR(25) => IR_out_25_port, IR(24) => IR_out_24_port, 
                           IR(23) => IR_out_23_port, IR(22) => IR_out_22_port, 
                           IR(21) => IR_out_21_port, IR(20) => IR_out_20_port, 
                           IR(19) => IR_out_19_port, IR(18) => n36, IR(17) => 
                           IR_out_17_port, IR(16) => IR_out_16_port, IR(15) => 
                           IR_out_15_port, IR(14) => IR_out_14_port, IR(13) => 
                           IR_out_13_port, IR(12) => IR_out_12_port, IR(11) => 
                           IR_out_11_port, IR(10) => IR_out_10_port, IR(9) => 
                           IR_out_9_port, IR(8) => IR_out_8_port, IR(7) => 
                           IR_out_7_port, IR(6) => IR_out_6_port, IR(5) => 
                           IR_out_5_port, IR(4) => IR_out_4_port, IR(3) => 
                           IR_out_3_port, IR(2) => IR_out_2_port, IR(1) => 
                           IR_out_1_port, IR(0) => IR_out_0_port, FWD_A(1) => 
                           FWDA_SEL_1_port, FWD_A(0) => FWDA_SEL_0_port, 
                           FWD_B(1) => FWDB_SEL_1_port, FWD_B(0) => 
                           FWDB_SEL_0_port, FWD_B2 => FWDB2_SEL, ZDU_SEL(1) => 
                           ZDU_SEL_1_port, ZDU_SEL(0) => ZDU_SEL_0_port);
   HDU1 : HDU_IR_SIZE32 port map( clk => CLK, rst => n51, IR(31) => 
                           IR_out_31_port, IR(30) => IR_out_30_port, IR(29) => 
                           IR_out_29_port, IR(28) => IR_out_28_port, IR(27) => 
                           IR_out_27_port, IR(26) => IR_out_26_port, IR(25) => 
                           IR_out_25_port, IR(24) => IR_out_24_port, IR(23) => 
                           IR_out_23_port, IR(22) => IR_out_22_port, IR(21) => 
                           IR_out_21_port, IR(20) => IR_out_20_port, IR(19) => 
                           IR_out_19_port, IR(18) => n36, IR(17) => 
                           IR_out_17_port, IR(16) => IR_out_16_port, IR(15) => 
                           IR_out_15_port, IR(14) => IR_out_14_port, IR(13) => 
                           IR_out_13_port, IR(12) => IR_out_12_port, IR(11) => 
                           IR_out_11_port, IR(10) => IR_out_10_port, IR(9) => 
                           IR_out_9_port, IR(8) => IR_out_8_port, IR(7) => 
                           IR_out_7_port, IR(6) => IR_out_6_port, IR(5) => 
                           IR_out_5_port, IR(4) => IR_out_4_port, IR(3) => 
                           IR_out_3_port, IR(2) => IR_out_2_port, IR(1) => 
                           IR_out_1_port, IR(0) => IR_out_0_port, STALL_CODE(1)
                           => STALL(1), STALL_CODE(0) => STALL(0), IF_STALL => 
                           IF_STALL, ID_STALL => n_1609, EX_STALL => EX_STALL, 
                           MEM_STALL => MEM_STALL, WB_STALL => n_1610);
   BHT1 : BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 port map( clock => CLK, rst => n51
                           , address(31) => BHT_in_31_port, address(30) => 
                           BHT_in_30_port, address(29) => BHT_in_29_port, 
                           address(28) => BHT_in_28_port, address(27) => 
                           BHT_in_27_port, address(26) => BHT_in_26_port, 
                           address(25) => BHT_in_25_port, address(24) => 
                           BHT_in_24_port, address(23) => BHT_in_23_port, 
                           address(22) => BHT_in_22_port, address(21) => 
                           BHT_in_21_port, address(20) => BHT_in_20_port, 
                           address(19) => BHT_in_19_port, address(18) => 
                           BHT_in_18_port, address(17) => BHT_in_17_port, 
                           address(16) => BHT_in_16_port, address(15) => 
                           BHT_in_15_port, address(14) => BHT_in_14_port, 
                           address(13) => BHT_in_13_port, address(12) => 
                           BHT_in_12_port, address(11) => BHT_in_11_port, 
                           address(10) => BHT_in_10_port, address(9) => 
                           BHT_in_9_port, address(8) => BHT_in_8_port, 
                           address(7) => BHT_in_7_port, address(6) => 
                           BHT_in_6_port, address(5) => BHT_in_5_port, 
                           address(4) => BHT_in_4_port, address(3) => 
                           BHT_in_3_port, address(2) => BHT_in_2_port, 
                           address(1) => BHT_in_1_port, address(0) => 
                           BHT_in_0_port, d_in => n19, w_en => n37, d_out => 
                           BHT_out);
   CWBU1 : CWBU port map( CLOCK => CLK, ALU_OP(0) => ALU_OPCODE(0), ALU_OP(1) 
                           => ALU_OPCODE(1), ALU_OP(2) => ALU_OPCODE(2), 
                           ALU_OP(3) => ALU_OPCODE(3), ALU_OP(4) => 
                           ALU_OPCODE(4), PSW(6) => PSW_out_6_port, PSW(5) => 
                           PSW_out_5_port, PSW(4) => PSW_out_4_port, PSW(3) => 
                           PSW_out_3_port, PSW(2) => PSW_out_2_port, PSW(1) => 
                           PSW_out_1_port, PSW(0) => PSW_out_0_port, 
                           COND_SEL(1) => CWB_out_1_port, COND_SEL(0) => 
                           CWB_out_0_port, CWB_SEL(1) => CWB_SEL(1), CWB_SEL(0)
                           => CWB_SEL(0), CWB_MUW_SEL(1) => CWB_MUX_SEL_1_port,
                           CWB_MUW_SEL(0) => CWB_MUX_SEL_0_port);
   RF1 : RF_NBIT32_NREG32 port map( CLK => CLK, RESET => n50, ENABLE => 
                           X_Logic1_port, RD1 => RF_RD_en, RD2 => RF_RD_en, WR 
                           => RF_WR, ADD_WR(4) => RF_MUX_out_4_port, ADD_WR(3) 
                           => RF_MUX_out_3_port, ADD_WR(2) => RF_MUX_out_2_port
                           , ADD_WR(1) => RF_MUX_out_1_port, ADD_WR(0) => 
                           RF_MUX_out_0_port, ADD_RD1(4) => IR_out_25_port, 
                           ADD_RD1(3) => IR_out_24_port, ADD_RD1(2) => 
                           IR_out_23_port, ADD_RD1(1) => IR_out_22_port, 
                           ADD_RD1(0) => IR_out_21_port, ADD_RD2(4) => 
                           IR_out_20_port, ADD_RD2(3) => IR_out_19_port, 
                           ADD_RD2(2) => n36, ADD_RD2(1) => IR_out_17_port, 
                           ADD_RD2(0) => IR_out_16_port, DATAIN(31) => 
                           WB_in_31_port, DATAIN(30) => WB_in_30_port, 
                           DATAIN(29) => WB_in_29_port, DATAIN(28) => 
                           WB_in_28_port, DATAIN(27) => WB_in_27_port, 
                           DATAIN(26) => WB_in_26_port, DATAIN(25) => 
                           WB_in_25_port, DATAIN(24) => WB_in_24_port, 
                           DATAIN(23) => WB_in_23_port, DATAIN(22) => 
                           WB_in_22_port, DATAIN(21) => WB_in_21_port, 
                           DATAIN(20) => WB_in_20_port, DATAIN(19) => 
                           WB_in_19_port, DATAIN(18) => WB_in_18_port, 
                           DATAIN(17) => WB_in_17_port, DATAIN(16) => 
                           WB_in_16_port, DATAIN(15) => WB_in_15_port, 
                           DATAIN(14) => WB_in_14_port, DATAIN(13) => 
                           WB_in_13_port, DATAIN(12) => WB_in_12_port, 
                           DATAIN(11) => WB_in_11_port, DATAIN(10) => 
                           WB_in_10_port, DATAIN(9) => WB_in_9_port, DATAIN(8) 
                           => WB_in_8_port, DATAIN(7) => WB_in_7_port, 
                           DATAIN(6) => WB_in_6_port, DATAIN(5) => WB_in_5_port
                           , DATAIN(4) => WB_in_4_port, DATAIN(3) => 
                           WB_in_3_port, DATAIN(2) => WB_in_2_port, DATAIN(1) 
                           => WB_in_1_port, DATAIN(0) => WB_in_0_port, OUT1(31)
                           => RA_out_31_port, OUT1(30) => RA_out_30_port, 
                           OUT1(29) => RA_out_29_port, OUT1(28) => 
                           RA_out_28_port, OUT1(27) => RA_out_27_port, OUT1(26)
                           => RA_out_26_port, OUT1(25) => RA_out_25_port, 
                           OUT1(24) => RA_out_24_port, OUT1(23) => 
                           RA_out_23_port, OUT1(22) => RA_out_22_port, OUT1(21)
                           => RA_out_21_port, OUT1(20) => RA_out_20_port, 
                           OUT1(19) => RA_out_19_port, OUT1(18) => 
                           RA_out_18_port, OUT1(17) => RA_out_17_port, OUT1(16)
                           => RA_out_16_port, OUT1(15) => RA_out_15_port, 
                           OUT1(14) => RA_out_14_port, OUT1(13) => 
                           RA_out_13_port, OUT1(12) => RA_out_12_port, OUT1(11)
                           => RA_out_11_port, OUT1(10) => RA_out_10_port, 
                           OUT1(9) => RA_out_9_port, OUT1(8) => RA_out_8_port, 
                           OUT1(7) => RA_out_7_port, OUT1(6) => RA_out_6_port, 
                           OUT1(5) => RA_out_5_port, OUT1(4) => RA_out_4_port, 
                           OUT1(3) => RA_out_3_port, OUT1(2) => RA_out_2_port, 
                           OUT1(1) => RA_out_1_port, OUT1(0) => RA_out_0_port, 
                           OUT2(31) => RB_out_31_port, OUT2(30) => 
                           RB_out_30_port, OUT2(29) => RB_out_29_port, OUT2(28)
                           => RB_out_28_port, OUT2(27) => RB_out_27_port, 
                           OUT2(26) => RB_out_26_port, OUT2(25) => 
                           RB_out_25_port, OUT2(24) => RB_out_24_port, OUT2(23)
                           => RB_out_23_port, OUT2(22) => RB_out_22_port, 
                           OUT2(21) => RB_out_21_port, OUT2(20) => 
                           RB_out_20_port, OUT2(19) => RB_out_19_port, OUT2(18)
                           => RB_out_18_port, OUT2(17) => RB_out_17_port, 
                           OUT2(16) => RB_out_16_port, OUT2(15) => 
                           RB_out_15_port, OUT2(14) => RB_out_14_port, OUT2(13)
                           => RB_out_13_port, OUT2(12) => RB_out_12_port, 
                           OUT2(11) => RB_out_11_port, OUT2(10) => 
                           RB_out_10_port, OUT2(9) => RB_out_9_port, OUT2(8) =>
                           RB_out_8_port, OUT2(7) => RB_out_7_port, OUT2(6) => 
                           RB_out_6_port, OUT2(5) => RB_out_5_port, OUT2(4) => 
                           RB_out_4_port, OUT2(3) => RB_out_3_port, OUT2(2) => 
                           RB_out_2_port, OUT2(1) => RB_out_1_port, OUT2(0) => 
                           RB_out_0_port);
   U3 : XNOR2_X1 port map( A => n7, B => RWB1_out_26_port, ZN => n19);
   U4 : BUF_X1 port map( A => n49, Z => n51);
   U5 : BUF_X1 port map( A => n49, Z => n50);
   U6 : BUF_X1 port map( A => n42, Z => n47);
   U7 : BUF_X1 port map( A => IR_out_18_port, Z => n36);
   U8 : BUF_X1 port map( A => EX_ENABLE, Z => n40);
   U9 : BUF_X1 port map( A => ID_ENABLE, Z => n41);
   U10 : BUF_X1 port map( A => n47, Z => n45);
   U11 : BUF_X1 port map( A => n47, Z => n44);
   U12 : BUF_X1 port map( A => n47, Z => n46);
   U13 : BUF_X1 port map( A => n48, Z => n43);
   U14 : BUF_X1 port map( A => n42, Z => n48);
   U15 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n7)
                           ;
   U16 : AND4_X1 port map( A1 => n12, A2 => n13, A3 => n14_port, A4 => n15, ZN 
                           => n11);
   U17 : NOR4_X1 port map( A1 => ZDU_MUX_out_19_port, A2 => ZDU_MUX_out_18_port
                           , A3 => ZDU_MUX_out_17_port, A4 => 
                           ZDU_MUX_out_16_port, ZN => n8);
   U18 : BUF_X1 port map( A => n53, Z => n38);
   U19 : INV_X1 port map( A => IF_STALL, ZN => n53);
   U20 : AND2_X1 port map( A1 => SIGND, A2 => IR_out_15_port, ZN => N14);
   U21 : NOR4_X1 port map( A1 => ZDU_MUX_out_9_port, A2 => ZDU_MUX_out_8_port, 
                           A3 => ZDU_MUX_out_7_port, A4 => ZDU_MUX_out_6_port, 
                           ZN => n15);
   U22 : NOR4_X1 port map( A1 => ZDU_MUX_out_5_port, A2 => ZDU_MUX_out_4_port, 
                           A3 => ZDU_MUX_out_3_port, A4 => ZDU_MUX_out_30_port,
                           ZN => n14_port);
   U23 : NOR4_X1 port map( A1 => n16, A2 => ZDU_MUX_out_0_port, A3 => 
                           ZDU_MUX_out_11_port, A4 => ZDU_MUX_out_10_port, ZN 
                           => n10);
   U24 : OR4_X1 port map( A1 => ZDU_MUX_out_13_port, A2 => ZDU_MUX_out_12_port,
                           A3 => ZDU_MUX_out_15_port, A4 => ZDU_MUX_out_14_port
                           , ZN => n16);
   U25 : NOR4_X1 port map( A1 => ZDU_MUX_out_22_port, A2 => ZDU_MUX_out_21_port
                           , A3 => ZDU_MUX_out_20_port, A4 => 
                           ZDU_MUX_out_1_port, ZN => n9);
   U26 : NOR4_X1 port map( A1 => ZDU_MUX_out_2_port, A2 => ZDU_MUX_out_29_port,
                           A3 => ZDU_MUX_out_28_port, A4 => ZDU_MUX_out_27_port
                           , ZN => n13);
   U27 : NOR4_X1 port map( A1 => ZDU_MUX_out_26_port, A2 => ZDU_MUX_out_25_port
                           , A3 => ZDU_MUX_out_24_port, A4 => 
                           ZDU_MUX_out_23_port, ZN => n12);
   U29 : NOR3_X1 port map( A1 => n17, A2 => PRD_OUT, A3 => n52, ZN => 
                           PC_SEL_1_port);
   U30 : INV_X1 port map( A => n18, ZN => n52);
   U31 : NOR2_X1 port map( A1 => EX_STALL, A2 => n55, ZN => EX_ENABLE);
   U32 : INV_X1 port map( A => EX_EN, ZN => n55);
   U33 : BUF_X1 port map( A => MEM_ENABLE, Z => n39);
   U34 : NOR2_X1 port map( A1 => MEM_STALL, A2 => n54, ZN => MEM_ENABLE);
   U35 : INV_X1 port map( A => MEM_EN, ZN => n54);
   U36 : BUF_X1 port map( A => DATA_IN(7), Z => n42);
   U37 : BUF_X1 port map( A => RST, Z => n49);
   U38 : AND2_X1 port map( A1 => n3, A2 => n37, ZN => BMP);
   U39 : INV_X1 port map( A => BMP, ZN => n17);
   U40 : AND2_X1 port map( A1 => PRD_OUT, A2 => BMP, ZN => IRAMMUX_SEL);
   U41 : CLKBUF_X1 port map( A => BPR_EN2, Z => n37);
   U42 : AND2_X1 port map( A1 => ID_EN, A2 => n38, ZN => ID_ENABLE);
   U43 : AND2_X1 port map( A1 => RF_RD, A2 => n38, ZN => RF_RD_en);
   U44 : AOI21_X1 port map( B1 => BPR_EN, B2 => BHT_out, A => UCB_EN, ZN => n18
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26 is

   port( Clk, Rst : in std_logic;  STALL : in std_logic_vector (1 downto 0);  
         IR_IN : in std_logic_vector (31 downto 0);  BMP : in std_logic;  ID_EN
         , RF_RD, SIGND, IMM_SEL, BPR_EN, UCB_EN : out std_logic;  ALU_OPCODE :
         out std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, ALUB_SEL, MEM_EN, 
         MEM_DATA_SEL, MEM_RD, MEM_WR, CS, MEM_BLC0, MEM_BLC1, LD_SEL0, LD_SEL1
         , LD_SEL2, ALR2_SEL, CWB_SEL0, CWB_SEL1, WB_SEL, RF_WR, RF_MUX_SEL0, 
         RF_MUX_SEL1 : out std_logic);

end CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26;

architecture SYN_dlx_cu_hw of 
   CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n48, n50, n51, n52, n189, n190, n191, n192, n3, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n49, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
      n91, n97, n98, n100, n102, n104, n105, n106, n107, n108, n109, n133, n135
      , n137, n139, n140, n141, n142, n143, n144, n145, n92, n93, n94, n95, n96
      , n99, n101, n103, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n_1611, n_1612, 
      n_1613, n_1614, n_1615 : std_logic;

begin
   
   cw5_reg_3_inst : DFFR_X1 port map( D => n133, CK => Clk, RN => n94, Q => 
                           WB_SEL, QN => n102);
   cw5_reg_2_inst : DFFR_X1 port map( D => n135, CK => Clk, RN => n96, Q => 
                           RF_WR, QN => n100);
   cw5_reg_1_inst : DFFR_X1 port map( D => n137, CK => Clk, RN => n94, Q => 
                           RF_MUX_SEL0, QN => n98);
   cw5_reg_0_inst : DFFR_X1 port map( D => n139, CK => Clk, RN => n94, Q => 
                           RF_MUX_SEL1, QN => n97);
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => n192, CK => Clk, RN => n94, Q
                           => n_1611, QN => n48);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => n141, CK => Clk, RN => n94, Q
                           => n_1612, QN => n108);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => n191, CK => Clk, RN => n94, Q
                           => n_1613, QN => n50);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => n190, CK => Clk, RN => n94, Q
                           => n_1614, QN => n51);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => n189, CK => Clk, RN => n94, Q
                           => n_1615, QN => n52);
   UCB_EN <= '0';
   BPR_EN <= '0';
   IMM_SEL <= '0';
   SIGND <= '0';
   RF_RD <= '0';
   ID_EN <= '0';
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => n140, CK => Clk, RN => n93, Q
                           => ALU_OPCODE(0), QN => n109);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => n143, CK => Clk, RN => n93, Q
                           => ALU_OPCODE(2), QN => n106);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => n142, CK => Clk, RN => n93, Q
                           => ALU_OPCODE(1), QN => n107);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => n145, CK => Clk, RN => n93, Q
                           => ALU_OPCODE(4), QN => n104);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => n144, CK => Clk, RN => n93, Q
                           => ALU_OPCODE(3), QN => n105);
   ALUB_SEL <= '0';
   ALUA_SEL <= '0';
   EX_EN <= '0';
   U123 : NAND3_X1 port map( A1 => n99, A2 => n125, A3 => n58, ZN => n57);
   U124 : NAND3_X1 port map( A1 => n64, A2 => n59, A3 => IR_IN(30), ZN => n61);
   U125 : NAND3_X1 port map( A1 => n113, A2 => n103, A3 => n64, ZN => n45);
   U126 : NAND3_X1 port map( A1 => n113, A2 => n103, A3 => n114, ZN => n88);
   U3 : NOR2_X2 port map( A1 => n100, A2 => n92, ZN => n135);
   U4 : NOR2_X2 port map( A1 => n97, A2 => n92, ZN => n139);
   U5 : NOR2_X2 port map( A1 => n98, A2 => n26, ZN => n137);
   U6 : NOR2_X2 port map( A1 => n102, A2 => n26, ZN => n133);
   U7 : OAI21_X1 port map( B1 => STALL(1), B2 => STALL(0), A => n25, ZN => n27)
                           ;
   U8 : BUF_X1 port map( A => n96, Z => n95);
   U9 : NAND2_X1 port map( A1 => n27, A2 => n25, ZN => n28);
   U10 : INV_X1 port map( A => n27, ZN => n3);
   U11 : INV_X1 port map( A => n67, ZN => n124);
   U12 : INV_X1 port map( A => n70, ZN => n120);
   U13 : NAND2_X1 port map( A1 => STALL(1), A2 => n25, ZN => n26);
   U14 : NAND2_X1 port map( A1 => STALL(1), A2 => n25, ZN => n92);
   U15 : OAI22_X1 port map( A1 => n119, A2 => n110, B1 => n43, B2 => n34, ZN =>
                           n31);
   U16 : AOI22_X1 port map( A1 => n36, A2 => n124, B1 => n120, B2 => n126, ZN 
                           => n43);
   U17 : OAI22_X1 port map( A1 => n117, A2 => n45, B1 => n62, B2 => n118, ZN =>
                           n42);
   U18 : NOR2_X1 port map( A1 => n115, A2 => n114, ZN => n64);
   U19 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => n34);
   U20 : NOR3_X1 port map( A1 => n67, A2 => n68, A3 => n123, ZN => n65);
   U21 : OAI21_X1 port map( B1 => n116, B2 => n56, A => n57, ZN => n41);
   U22 : INV_X1 port map( A => n59, ZN => n116);
   U23 : INV_X1 port map( A => n34, ZN => n99);
   U30 : AOI21_X1 port map( B1 => n36, B2 => n126, A => n37, ZN => n33);
   U31 : INV_X1 port map( A => n49, ZN => n126);
   U32 : NAND2_X1 port map( A1 => n127, A2 => n125, ZN => n67);
   U33 : INV_X1 port map( A => n53, ZN => n110);
   U34 : NAND2_X1 port map( A1 => n46, A2 => n119, ZN => n59);
   U35 : NAND2_X1 port map( A1 => n77, A2 => n113, ZN => n62);
   U36 : NAND2_X1 port map( A1 => n83, A2 => n123, ZN => n70);
   U37 : INV_X1 port map( A => n78, ZN => n119);
   U38 : INV_X1 port map( A => n71, ZN => n121);
   U39 : INV_X1 port map( A => n63, ZN => n117);
   U40 : BUF_X1 port map( A => n95, Z => n94);
   U41 : BUF_X1 port map( A => n95, Z => n93);
   U42 : OAI22_X1 port map( A1 => n105, A2 => n27, B1 => n51, B2 => n28, ZN => 
                           n144);
   U43 : OAI22_X1 port map( A1 => n104, A2 => n27, B1 => n52, B2 => n28, ZN => 
                           n145);
   U44 : OAI22_X1 port map( A1 => n107, A2 => n27, B1 => n108, B2 => n28, ZN =>
                           n142);
   U45 : OAI22_X1 port map( A1 => n106, A2 => n27, B1 => n50, B2 => n28, ZN => 
                           n143);
   U46 : OAI22_X1 port map( A1 => n109, A2 => n27, B1 => n48, B2 => n28, ZN => 
                           n140);
   U47 : OAI22_X1 port map( A1 => n48, A2 => n27, B1 => n3, B2 => n38, ZN => 
                           n192);
   U48 : OAI22_X1 port map( A1 => n52, A2 => n27, B1 => n3, B2 => n72, ZN => 
                           n189);
   U49 : AOI211_X1 port map( C1 => n53, C2 => n63, A => n73, B => n74, ZN => 
                           n72);
   U50 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n38, A4 => n45, ZN => 
                           n73);
   U51 : OAI22_X1 port map( A1 => n75, A2 => n34, B1 => n76, B2 => n46, ZN => 
                           n74);
   U52 : OAI22_X1 port map( A1 => n51, A2 => n27, B1 => n3, B2 => n54, ZN => 
                           n190);
   U53 : NOR3_X1 port map( A1 => n55, A2 => n32, A3 => n41, ZN => n54);
   U54 : OAI221_X1 port map( B1 => n69, B2 => n34, C1 => n45, C2 => n119, A => 
                           n38, ZN => n55);
   U55 : AOI22_X1 port map( A1 => n124, A2 => n121, B1 => n120, B2 => IR_IN(1),
                           ZN => n69);
   U56 : OAI22_X1 port map( A1 => n50, A2 => n27, B1 => n3, B2 => n39, ZN => 
                           n191);
   U57 : NOR4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n31, ZN => 
                           n39);
   U58 : OAI222_X1 port map( A1 => n118, A2 => n110, B1 => n44, B2 => n34, C1 
                           => n45, C2 => n46, ZN => n40);
   U59 : AOI22_X1 port map( A1 => n121, A2 => n47, B1 => n36, B2 => IR_IN(1), 
                           ZN => n44);
   U60 : OAI22_X1 port map( A1 => n108, A2 => n27, B1 => n3, B2 => n29, ZN => 
                           n141);
   U61 : NOR3_X1 port map( A1 => n30, A2 => n31, A3 => n32, ZN => n29);
   U62 : OAI221_X1 port map( B1 => n33, B2 => n34, C1 => n117, C2 => n110, A =>
                           n35, ZN => n30);
   U63 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(27), A3 => IR_IN(29), 
                           A4 => n115, ZN => n35);
   U64 : NOR4_X1 port map( A1 => IR_IN(28), A2 => IR_IN(9), A3 => n88, A4 => 
                           n89, ZN => n79);
   U65 : OR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), A3 => IR_IN(8), A4 
                           => IR_IN(7), ZN => n89);
   U66 : NOR4_X1 port map( A1 => n113, A2 => n115, A3 => IR_IN(29), A4 => 
                           IR_IN(31), ZN => n53);
   U67 : NOR3_X1 port map( A1 => IR_IN(28), A2 => IR_IN(31), A3 => n114, ZN => 
                           n77);
   U68 : NOR2_X1 port map( A1 => n84, A2 => IR_IN(3), ZN => n36);
   U69 : NOR3_X1 port map( A1 => n68, A2 => IR_IN(2), A3 => n125, ZN => n37);
   U70 : NOR3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(4), A3 => n122, ZN => 
                           n83);
   U71 : INV_X1 port map( A => IR_IN(5), ZN => n122);
   U72 : AOI211_X1 port map( C1 => n36, C2 => n126, A => n80, B => n66, ZN => 
                           n75);
   U73 : OAI221_X1 port map( B1 => n67, B2 => n70, C1 => IR_IN(1), C2 => n71, A
                           => n82, ZN => n80);
   U74 : OAI21_X1 port map( B1 => n37, B2 => n58, A => IR_IN(0), ZN => n82);
   U75 : NOR3_X1 port map( A1 => IR_IN(2), A2 => IR_IN(4), A3 => n68, ZN => n58
                           );
   U76 : NAND4_X1 port map( A1 => IR_IN(3), A2 => n79, A3 => n126, A4 => n87, 
                           ZN => n38);
   U77 : NOR2_X1 port map( A1 => n84, A2 => n46, ZN => n87);
   U78 : OAI211_X1 port map( C1 => n60, C2 => n34, A => n61, B => n101, ZN => 
                           n32);
   U79 : INV_X1 port map( A => n42, ZN => n101);
   U80 : NOR2_X1 port map( A1 => n65, A2 => n66, ZN => n60);
   U81 : OAI21_X1 port map( B1 => n71, B2 => n49, A => n81, ZN => n66);
   U82 : OR4_X1 port map( A1 => n123, A2 => n127, A3 => n68, A4 => IR_IN(1), ZN
                           => n81);
   U83 : NOR2_X1 port map( A1 => n118, A2 => IR_IN(26), ZN => n63);
   U84 : NOR2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n78);
   U85 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n118, ZN => n46);
   U86 : AOI21_X1 port map( B1 => IR_IN(30), B2 => n64, A => n112, ZN => n76);
   U87 : INV_X1 port map( A => n56, ZN => n112);
   U88 : NAND2_X1 port map( A1 => IR_IN(5), A2 => IR_IN(3), ZN => n68);
   U89 : INV_X1 port map( A => IR_IN(28), ZN => n115);
   U90 : INV_X1 port map( A => IR_IN(30), ZN => n113);
   U91 : INV_X1 port map( A => IR_IN(27), ZN => n118);
   U92 : OAI21_X1 port map( B1 => IR_IN(1), B2 => n127, A => n49, ZN => n47);
   U93 : NAND2_X1 port map( A1 => n83, A2 => IR_IN(2), ZN => n71);
   U94 : INV_X1 port map( A => IR_IN(2), ZN => n123);
   U95 : OAI21_X1 port map( B1 => n91, B2 => n111, A => n59, ZN => n85);
   U96 : INV_X1 port map( A => n62, ZN => n111);
   U97 : NOR3_X1 port map( A1 => n103, A2 => IR_IN(30), A3 => n64, ZN => n91);
   U98 : NAND2_X1 port map( A1 => IR_IN(1), A2 => n127, ZN => n49);
   U99 : NAND4_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), A3 => n90, A4 => 
                           n115, ZN => n86);
   U100 : OAI22_X1 port map( A1 => IR_IN(30), A2 => n103, B1 => n114, B2 => 
                           n113, ZN => n90);
   U101 : INV_X1 port map( A => IR_IN(29), ZN => n114);
   U102 : INV_X1 port map( A => IR_IN(0), ZN => n127);
   U103 : INV_X1 port map( A => IR_IN(31), ZN => n103);
   U104 : NAND2_X1 port map( A1 => IR_IN(30), A2 => n77, ZN => n56);
   U105 : INV_X1 port map( A => IR_IN(1), ZN => n125);
   U106 : OR3_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), A3 => n123, ZN => 
                           n84);
   U107 : INV_X1 port map( A => Rst, ZN => n96);
   MEM_DATA_SEL <= '0';
   MEM_WR <= '0';
   MEM_BLC0 <= '0';
   LD_SEL0 <= '0';
   LD_SEL2 <= '0';
   CWB_SEL0 <= '0';
   CWB_SEL1 <= '0';
   CS <= '0';
   MEM_RD <= '0';
   LD_SEL1 <= '0';
   MEM_BLC1 <= '0';
   ALR2_SEL <= '0';
   MEM_EN <= '0';
   U121 : INV_X1 port map( A => BMP, ZN => n25);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector (31 
         downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out std_logic_vector (31 
         downto 0);  BLC : out std_logic_vector (1 downto 0);  MEM_WR, MEM_RD :
         out std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component Datapath
      port( CLK, RST : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector 
            (31 downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out 
            std_logic_vector (31 downto 0);  BMP : inout std_logic;  STALL : 
            out std_logic_vector (1 downto 0);  ID_EN, RF_RD, SIGND, IMM_SEL, 
            BPR_EN : in std_logic;  ALU_OPCODE : in std_logic_vector (0 to 4); 
            EX_EN, ALUA_SEL, ALUB_SEL, UCB_EN, MEM_EN, MEM_DATA_SEL : in 
            std_logic;  LD_SEL : in std_logic_vector (2 downto 0);  ALR2_SEL : 
            in std_logic;  CWB_SEL : in std_logic_vector (1 downto 0);  WB_SEL,
            RF_WR : in std_logic;  RF_MUX_SEL : in std_logic_vector (1 downto 
            0));
   end component;
   
   component 
      CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26
      port( Clk, Rst : in std_logic;  STALL : in std_logic_vector (1 downto 0);
            IR_IN : in std_logic_vector (31 downto 0);  BMP : in std_logic;  
            ID_EN, RF_RD, SIGND, IMM_SEL, BPR_EN, UCB_EN : out std_logic;  
            ALU_OPCODE : out std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, 
            ALUB_SEL, MEM_EN, MEM_DATA_SEL, MEM_RD, MEM_WR, CS, MEM_BLC0, 
            MEM_BLC1, LD_SEL0, LD_SEL1, LD_SEL2, ALR2_SEL, CWB_SEL0, CWB_SEL1, 
            WB_SEL, RF_WR, RF_MUX_SEL0, RF_MUX_SEL1 : out std_logic);
   end component;
   
   signal STALL_CODE_1_port, STALL_CODE_0_port, BMP_i, ID_EN_i, RF_RD_i, 
      SIGND_i, IMM_SEL_i, BPR_EN_i, UCB_EN_i, ALU_OPCODE_i_0_port, 
      ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_4_port, WB_SEL_i, RF_WR_i, RF_MUX_SEL_i_1_port, 
      RF_MUX_SEL_i_0_port, n1, MEM_WR_port, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637 : 
      std_logic;

begin
   BLC <= ( MEM_WR_port, MEM_WR_port );
   MEM_WR <= MEM_WR_port;
   MEM_RD <= MEM_WR_port;
   
   n1 <= '0';
   UCB_EN_i <= '0';
   BPR_EN_i <= '0';
   IMM_SEL_i <= '0';
   SIGND_i <= '0';
   RF_RD_i <= '0';
   ID_EN_i <= '0';
   CU_I : CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26
                           port map( Clk => Clk, Rst => Rst, STALL(1) => 
                           STALL_CODE_1_port, STALL(0) => STALL_CODE_0_port, 
                           IR_IN(31) => IRAM_OUT(31), IR_IN(30) => IRAM_OUT(30)
                           , IR_IN(29) => IRAM_OUT(29), IR_IN(28) => 
                           IRAM_OUT(28), IR_IN(27) => IRAM_OUT(27), IR_IN(26) 
                           => IRAM_OUT(26), IR_IN(25) => IRAM_OUT(25), 
                           IR_IN(24) => IRAM_OUT(24), IR_IN(23) => IRAM_OUT(23)
                           , IR_IN(22) => IRAM_OUT(22), IR_IN(21) => 
                           IRAM_OUT(21), IR_IN(20) => IRAM_OUT(20), IR_IN(19) 
                           => IRAM_OUT(19), IR_IN(18) => IRAM_OUT(18), 
                           IR_IN(17) => IRAM_OUT(17), IR_IN(16) => IRAM_OUT(16)
                           , IR_IN(15) => IRAM_OUT(15), IR_IN(14) => 
                           IRAM_OUT(14), IR_IN(13) => IRAM_OUT(13), IR_IN(12) 
                           => IRAM_OUT(12), IR_IN(11) => IRAM_OUT(11), 
                           IR_IN(10) => IRAM_OUT(10), IR_IN(9) => IRAM_OUT(9), 
                           IR_IN(8) => IRAM_OUT(8), IR_IN(7) => IRAM_OUT(7), 
                           IR_IN(6) => IRAM_OUT(6), IR_IN(5) => IRAM_OUT(5), 
                           IR_IN(4) => IRAM_OUT(4), IR_IN(3) => IRAM_OUT(3), 
                           IR_IN(2) => IRAM_OUT(2), IR_IN(1) => IRAM_OUT(1), 
                           IR_IN(0) => IRAM_OUT(0), BMP => BMP_i, ID_EN => 
                           n_1616, RF_RD => n_1617, SIGND => n_1618, IMM_SEL =>
                           n_1619, BPR_EN => n_1620, UCB_EN => n_1621, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_0_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, EX_EN => n_1622, ALUA_SEL => 
                           n_1623, ALUB_SEL => n_1624, MEM_EN => n_1625, 
                           MEM_DATA_SEL => n_1626, MEM_RD => n_1627, MEM_WR => 
                           n_1628, CS => n_1629, MEM_BLC0 => n_1630, MEM_BLC1 
                           => n_1631, LD_SEL0 => n_1632, LD_SEL1 => n_1633, 
                           LD_SEL2 => n_1634, ALR2_SEL => n_1635, CWB_SEL0 => 
                           n_1636, CWB_SEL1 => n_1637, WB_SEL => WB_SEL_i, 
                           RF_WR => RF_WR_i, RF_MUX_SEL0 => RF_MUX_SEL_i_0_port
                           , RF_MUX_SEL1 => RF_MUX_SEL_i_1_port);
   DATAP : Datapath port map( CLK => Clk, RST => Rst, DATA_IN(31) => 
                           DATA_IN(31), DATA_IN(30) => DATA_IN(30), DATA_IN(29)
                           => DATA_IN(29), DATA_IN(28) => DATA_IN(28), 
                           DATA_IN(27) => DATA_IN(27), DATA_IN(26) => 
                           DATA_IN(26), DATA_IN(25) => DATA_IN(25), DATA_IN(24)
                           => DATA_IN(24), DATA_IN(23) => DATA_IN(23), 
                           DATA_IN(22) => DATA_IN(22), DATA_IN(21) => 
                           DATA_IN(21), DATA_IN(20) => DATA_IN(20), DATA_IN(19)
                           => DATA_IN(19), DATA_IN(18) => DATA_IN(18), 
                           DATA_IN(17) => DATA_IN(17), DATA_IN(16) => 
                           DATA_IN(16), DATA_IN(15) => DATA_IN(15), DATA_IN(14)
                           => DATA_IN(14), DATA_IN(13) => DATA_IN(13), 
                           DATA_IN(12) => DATA_IN(12), DATA_IN(11) => 
                           DATA_IN(11), DATA_IN(10) => DATA_IN(10), DATA_IN(9) 
                           => DATA_IN(9), DATA_IN(8) => DATA_IN(8), DATA_IN(7) 
                           => DATA_IN(7), DATA_IN(6) => DATA_IN(6), DATA_IN(5) 
                           => DATA_IN(5), DATA_IN(4) => DATA_IN(4), DATA_IN(3) 
                           => DATA_IN(3), DATA_IN(2) => DATA_IN(2), DATA_IN(1) 
                           => DATA_IN(1), DATA_IN(0) => DATA_IN(0), 
                           IRAM_OUT(31) => IRAM_OUT(31), IRAM_OUT(30) => 
                           IRAM_OUT(30), IRAM_OUT(29) => IRAM_OUT(29), 
                           IRAM_OUT(28) => IRAM_OUT(28), IRAM_OUT(27) => 
                           IRAM_OUT(27), IRAM_OUT(26) => IRAM_OUT(26), 
                           IRAM_OUT(25) => IRAM_OUT(25), IRAM_OUT(24) => 
                           IRAM_OUT(24), IRAM_OUT(23) => IRAM_OUT(23), 
                           IRAM_OUT(22) => IRAM_OUT(22), IRAM_OUT(21) => 
                           IRAM_OUT(21), IRAM_OUT(20) => IRAM_OUT(20), 
                           IRAM_OUT(19) => IRAM_OUT(19), IRAM_OUT(18) => 
                           IRAM_OUT(18), IRAM_OUT(17) => IRAM_OUT(17), 
                           IRAM_OUT(16) => IRAM_OUT(16), IRAM_OUT(15) => 
                           IRAM_OUT(15), IRAM_OUT(14) => IRAM_OUT(14), 
                           IRAM_OUT(13) => IRAM_OUT(13), IRAM_OUT(12) => 
                           IRAM_OUT(12), IRAM_OUT(11) => IRAM_OUT(11), 
                           IRAM_OUT(10) => IRAM_OUT(10), IRAM_OUT(9) => 
                           IRAM_OUT(9), IRAM_OUT(8) => IRAM_OUT(8), IRAM_OUT(7)
                           => IRAM_OUT(7), IRAM_OUT(6) => IRAM_OUT(6), 
                           IRAM_OUT(5) => IRAM_OUT(5), IRAM_OUT(4) => 
                           IRAM_OUT(4), IRAM_OUT(3) => IRAM_OUT(3), IRAM_OUT(2)
                           => IRAM_OUT(2), IRAM_OUT(1) => IRAM_OUT(1), 
                           IRAM_OUT(0) => IRAM_OUT(0), IRAM_ADDR(31) => 
                           IRAM_ADDR(31), IRAM_ADDR(30) => IRAM_ADDR(30), 
                           IRAM_ADDR(29) => IRAM_ADDR(29), IRAM_ADDR(28) => 
                           IRAM_ADDR(28), IRAM_ADDR(27) => IRAM_ADDR(27), 
                           IRAM_ADDR(26) => IRAM_ADDR(26), IRAM_ADDR(25) => 
                           IRAM_ADDR(25), IRAM_ADDR(24) => IRAM_ADDR(24), 
                           IRAM_ADDR(23) => IRAM_ADDR(23), IRAM_ADDR(22) => 
                           IRAM_ADDR(22), IRAM_ADDR(21) => IRAM_ADDR(21), 
                           IRAM_ADDR(20) => IRAM_ADDR(20), IRAM_ADDR(19) => 
                           IRAM_ADDR(19), IRAM_ADDR(18) => IRAM_ADDR(18), 
                           IRAM_ADDR(17) => IRAM_ADDR(17), IRAM_ADDR(16) => 
                           IRAM_ADDR(16), IRAM_ADDR(15) => IRAM_ADDR(15), 
                           IRAM_ADDR(14) => IRAM_ADDR(14), IRAM_ADDR(13) => 
                           IRAM_ADDR(13), IRAM_ADDR(12) => IRAM_ADDR(12), 
                           IRAM_ADDR(11) => IRAM_ADDR(11), IRAM_ADDR(10) => 
                           IRAM_ADDR(10), IRAM_ADDR(9) => IRAM_ADDR(9), 
                           IRAM_ADDR(8) => IRAM_ADDR(8), IRAM_ADDR(7) => 
                           IRAM_ADDR(7), IRAM_ADDR(6) => IRAM_ADDR(6), 
                           IRAM_ADDR(5) => IRAM_ADDR(5), IRAM_ADDR(4) => 
                           IRAM_ADDR(4), IRAM_ADDR(3) => IRAM_ADDR(3), 
                           IRAM_ADDR(2) => IRAM_ADDR(2), IRAM_ADDR(1) => 
                           IRAM_ADDR(1), IRAM_ADDR(0) => IRAM_ADDR(0), 
                           DATA_OUT(31) => DATA_OUT(31), DATA_OUT(30) => 
                           DATA_OUT(30), DATA_OUT(29) => DATA_OUT(29), 
                           DATA_OUT(28) => DATA_OUT(28), DATA_OUT(27) => 
                           DATA_OUT(27), DATA_OUT(26) => DATA_OUT(26), 
                           DATA_OUT(25) => DATA_OUT(25), DATA_OUT(24) => 
                           DATA_OUT(24), DATA_OUT(23) => DATA_OUT(23), 
                           DATA_OUT(22) => DATA_OUT(22), DATA_OUT(21) => 
                           DATA_OUT(21), DATA_OUT(20) => DATA_OUT(20), 
                           DATA_OUT(19) => DATA_OUT(19), DATA_OUT(18) => 
                           DATA_OUT(18), DATA_OUT(17) => DATA_OUT(17), 
                           DATA_OUT(16) => DATA_OUT(16), DATA_OUT(15) => 
                           DATA_OUT(15), DATA_OUT(14) => DATA_OUT(14), 
                           DATA_OUT(13) => DATA_OUT(13), DATA_OUT(12) => 
                           DATA_OUT(12), DATA_OUT(11) => DATA_OUT(11), 
                           DATA_OUT(10) => DATA_OUT(10), DATA_OUT(9) => 
                           DATA_OUT(9), DATA_OUT(8) => DATA_OUT(8), DATA_OUT(7)
                           => DATA_OUT(7), DATA_OUT(6) => DATA_OUT(6), 
                           DATA_OUT(5) => DATA_OUT(5), DATA_OUT(4) => 
                           DATA_OUT(4), DATA_OUT(3) => DATA_OUT(3), DATA_OUT(2)
                           => DATA_OUT(2), DATA_OUT(1) => DATA_OUT(1), 
                           DATA_OUT(0) => DATA_OUT(0), DATA_ADDR(31) => 
                           DATA_ADDR(31), DATA_ADDR(30) => DATA_ADDR(30), 
                           DATA_ADDR(29) => DATA_ADDR(29), DATA_ADDR(28) => 
                           DATA_ADDR(28), DATA_ADDR(27) => DATA_ADDR(27), 
                           DATA_ADDR(26) => DATA_ADDR(26), DATA_ADDR(25) => 
                           DATA_ADDR(25), DATA_ADDR(24) => DATA_ADDR(24), 
                           DATA_ADDR(23) => DATA_ADDR(23), DATA_ADDR(22) => 
                           DATA_ADDR(22), DATA_ADDR(21) => DATA_ADDR(21), 
                           DATA_ADDR(20) => DATA_ADDR(20), DATA_ADDR(19) => 
                           DATA_ADDR(19), DATA_ADDR(18) => DATA_ADDR(18), 
                           DATA_ADDR(17) => DATA_ADDR(17), DATA_ADDR(16) => 
                           DATA_ADDR(16), DATA_ADDR(15) => DATA_ADDR(15), 
                           DATA_ADDR(14) => DATA_ADDR(14), DATA_ADDR(13) => 
                           DATA_ADDR(13), DATA_ADDR(12) => DATA_ADDR(12), 
                           DATA_ADDR(11) => DATA_ADDR(11), DATA_ADDR(10) => 
                           DATA_ADDR(10), DATA_ADDR(9) => DATA_ADDR(9), 
                           DATA_ADDR(8) => DATA_ADDR(8), DATA_ADDR(7) => 
                           DATA_ADDR(7), DATA_ADDR(6) => DATA_ADDR(6), 
                           DATA_ADDR(5) => DATA_ADDR(5), DATA_ADDR(4) => 
                           DATA_ADDR(4), DATA_ADDR(3) => DATA_ADDR(3), 
                           DATA_ADDR(2) => DATA_ADDR(2), DATA_ADDR(1) => 
                           DATA_ADDR(1), DATA_ADDR(0) => DATA_ADDR(0), BMP => 
                           BMP_i, STALL(1) => STALL_CODE_1_port, STALL(0) => 
                           STALL_CODE_0_port, ID_EN => ID_EN_i, RF_RD => 
                           RF_RD_i, SIGND => SIGND_i, IMM_SEL => IMM_SEL_i, 
                           BPR_EN => BPR_EN_i, ALU_OPCODE(0) => 
                           ALU_OPCODE_i_0_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, EX_EN => n1, ALUA_SEL => n1, 
                           ALUB_SEL => n1, UCB_EN => UCB_EN_i, MEM_EN => 
                           MEM_WR_port, MEM_DATA_SEL => MEM_WR_port, LD_SEL(2) 
                           => MEM_WR_port, LD_SEL(1) => MEM_WR_port, LD_SEL(0) 
                           => MEM_WR_port, ALR2_SEL => MEM_WR_port, CWB_SEL(1) 
                           => MEM_WR_port, CWB_SEL(0) => MEM_WR_port, WB_SEL =>
                           WB_SEL_i, RF_WR => RF_WR_i, RF_MUX_SEL(1) => 
                           RF_MUX_SEL_i_1_port, RF_MUX_SEL(0) => 
                           RF_MUX_SEL_i_0_port);
   MEM_WR_port <= '0';

end SYN_dlx_rtl;
