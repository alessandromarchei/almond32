
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_NOP, OP_ADD, OP_ADC, OP_AND, OP_SRA, OP_OR, OP_SEQ, OP_SNE, 
   OP_SLT, OP_SGT, OP_SLE, OP_SGE, OP_SLL, OP_SRL, OP_SUB, OP_XOR, OP_NOR, 
   OP_XNOR, OP_NAND, OP_MUL);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011";

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HDU_IR_SIZE32_DW01_dec_1 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end HDU_IR_SIZE32_DW01_dec_1;

architecture SYN_cla of HDU_IR_SIZE32_DW01_dec_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n34, A2 => n27, ZN => n41);
   U3 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => n91);
   U4 : NOR2_X1 port map( A1 => n103, A2 => n104, ZN => n95);
   U5 : NOR2_X1 port map( A1 => n97, A2 => n98, ZN => n96);
   U6 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => n30);
   U7 : NOR2_X1 port map( A1 => n35, A2 => n36, ZN => n33);
   U8 : NAND2_X1 port map( A1 => n37, A2 => n32, ZN => n36);
   U9 : INV_X1 port map( A => n29, ZN => n28);
   U10 : NAND2_X1 port map( A1 => n60, A2 => n80, ZN => n76);
   U11 : NAND2_X1 port map( A1 => n70, A2 => n65, ZN => n74);
   U12 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => SUM(8));
   U13 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => SUM(9));
   U14 : INV_X1 port map( A => A(9), ZN => n2);
   U15 : NAND2_X1 port map( A1 => n123, A2 => n124, ZN => SUM(10));
   U16 : NAND2_X1 port map( A1 => A(10), A2 => n3, ZN => n124);
   U17 : INV_X1 port map( A => A(11), ZN => n119);
   U18 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => SUM(12));
   U19 : NAND2_X1 port map( A1 => A(12), A2 => n116, ZN => n115);
   U20 : OAI21_X1 port map( B1 => n110, B2 => n111, A => n109, ZN => SUM(13));
   U21 : INV_X1 port map( A => A(13), ZN => n111);
   U22 : XNOR2_X1 port map( A => A(14), B => n109, ZN => SUM(14));
   U23 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n91, ZN => SUM(15));
   U24 : INV_X1 port map( A => A(15), ZN => n94);
   U25 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => SUM(16));
   U26 : NAND2_X1 port map( A1 => A(16), A2 => n91, ZN => n90);
   U27 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n85, ZN => SUM(17));
   U28 : INV_X1 port map( A => A(17), ZN => n87);
   U29 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => SUM(18));
   U30 : NAND2_X1 port map( A1 => A(18), A2 => n85, ZN => n84);
   U31 : INV_X1 port map( A => A(19), ZN => n79);
   U32 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => SUM(20));
   U33 : NAND2_X1 port map( A1 => A(20), A2 => n76, ZN => n75);
   U34 : OAI21_X1 port map( B1 => n72, B2 => n64, A => n71, ZN => SUM(21));
   U35 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n66, ZN => SUM(22));
   U36 : INV_X1 port map( A => A(22), ZN => n68);
   U37 : INV_X1 port map( A => A(23), ZN => n58);
   U38 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => SUM(24));
   U39 : NAND2_X1 port map( A1 => A(24), A2 => n29, ZN => n55);
   U40 : INV_X1 port map( A => A(25), ZN => n52);
   U41 : INV_X1 port map( A => A(26), ZN => n48);
   U42 : INV_X1 port map( A => A(27), ZN => n43);
   U43 : XNOR2_X1 port map( A => A(30), B => n30, ZN => SUM(30));
   U44 : XNOR2_X1 port map( A => A(31), B => n25, ZN => SUM(31));
   U45 : NAND4_X1 port map( A1 => n26, A2 => n32, A3 => n27, A4 => n28, ZN => 
                           n25);
   U46 : XNOR2_X1 port map( A => A(2), B => n24, ZN => SUM(2));
   U47 : OAI21_X1 port map( B1 => n20, B2 => n21, A => n18, ZN => SUM(3));
   U48 : INV_X1 port map( A => A(3), ZN => n21);
   U49 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => SUM(4));
   U50 : NAND2_X1 port map( A1 => A(4), A2 => n18, ZN => n17);
   U51 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n11, ZN => SUM(5));
   U52 : INV_X1 port map( A => A(5), ZN => n13);
   U53 : XNOR2_X1 port map( A => A(6), B => n11, ZN => SUM(6));
   U54 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n6, ZN => SUM(7));
   U55 : INV_X1 port map( A => A(7), ZN => n10);
   U56 : NAND2_X1 port map( A1 => n24, A2 => n77, ZN => SUM(1));
   U57 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => n29);
   U58 : NOR2_X1 port map( A1 => n61, A2 => n62, ZN => n59);
   U59 : NOR2_X1 port map( A1 => A(23), A2 => A(22), ZN => n63);
   U60 : NOR2_X1 port map( A1 => A(3), A2 => A(2), ZN => n99);
   U61 : NOR2_X1 port map( A1 => A(5), A2 => A(4), ZN => n100);
   U62 : NOR2_X1 port map( A1 => A(12), A2 => A(11), ZN => n106);
   U63 : NOR2_X1 port map( A1 => A(10), A2 => A(0), ZN => n105);
   U64 : NOR2_X1 port map( A1 => A(7), A2 => A(6), ZN => n101);
   U65 : NOR2_X1 port map( A1 => A(9), A2 => A(8), ZN => n102);
   U66 : NAND2_X1 port map( A1 => n34, A2 => n56, ZN => n54);
   U67 : INV_X1 port map( A => A(24), ZN => n56);
   U68 : NOR2_X1 port map( A1 => A(1), A2 => A(15), ZN => n108);
   U69 : NAND2_X1 port map( A1 => n40, A2 => n34, ZN => n38);
   U70 : NOR2_X1 port map( A1 => A(28), A2 => n35, ZN => n40);
   U71 : NAND2_X1 port map( A1 => n53, A2 => n34, ZN => n50);
   U72 : NOR2_X1 port map( A1 => A(25), A2 => A(24), ZN => n53);
   U73 : NAND2_X1 port map( A1 => n49, A2 => n34, ZN => n46);
   U74 : NOR3_X1 port map( A1 => A(24), A2 => A(26), A3 => A(25), ZN => n49);
   U75 : NOR2_X1 port map( A1 => A(14), A2 => A(13), ZN => n107);
   U76 : NAND2_X1 port map( A1 => n73, A2 => n70, ZN => n71);
   U77 : NOR2_X1 port map( A1 => A(21), A2 => A(20), ZN => n73);
   U78 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => n66);
   U79 : NOR3_X1 port map( A1 => A(20), A2 => A(22), A3 => A(21), ZN => n69);
   U80 : NAND2_X1 port map( A1 => n88, A2 => n60, ZN => n85);
   U81 : NOR2_X1 port map( A1 => A(17), A2 => A(16), ZN => n88);
   U82 : OR2_X1 port map( A1 => n85, A2 => A(18), ZN => n83);
   U83 : NAND4_X1 port map( A1 => n126, A2 => n127, A3 => n128, A4 => n129, ZN 
                           => n6);
   U84 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n126);
   U85 : NOR2_X1 port map( A1 => A(7), A2 => A(6), ZN => n129);
   U86 : NOR2_X1 port map( A1 => A(3), A2 => A(2), ZN => n127);
   U87 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => n109);
   U88 : NOR2_X1 port map( A1 => A(13), A2 => A(12), ZN => n112);
   U89 : NOR2_X1 port map( A1 => A(5), A2 => A(4), ZN => n128);
   U90 : NOR2_X1 port map( A1 => A(14), A2 => n109, ZN => n93);
   U91 : NAND2_X1 port map( A1 => n120, A2 => n7, ZN => n116);
   U92 : AND2_X1 port map( A1 => n121, A2 => n122, ZN => n120);
   U93 : NOR2_X1 port map( A1 => A(9), A2 => A(11), ZN => n122);
   U94 : NOR2_X1 port map( A1 => A(8), A2 => A(10), ZN => n121);
   U95 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n61);
   U96 : NOR2_X1 port map( A1 => A(19), A2 => A(18), ZN => n82);
   U97 : NOR2_X1 port map( A1 => A(17), A2 => A(16), ZN => n81);
   U98 : INV_X1 port map( A => A(20), ZN => n65);
   U99 : NAND2_X1 port map( A1 => n113, A2 => n117, ZN => n114);
   U100 : INV_X1 port map( A => A(12), ZN => n117);
   U101 : INV_X1 port map( A => A(21), ZN => n64);
   U102 : NAND2_X1 port map( A1 => n60, A2 => n92, ZN => n89);
   U103 : INV_X1 port map( A => A(16), ZN => n92);
   U104 : NAND2_X1 port map( A1 => n125, A2 => n7, ZN => n3);
   U105 : NOR2_X1 port map( A1 => A(9), A2 => A(8), ZN => n125);
   U106 : OR2_X1 port map( A1 => n3, A2 => A(10), ZN => n123);
   U107 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n11);
   U108 : NOR2_X1 port map( A1 => A(5), A2 => A(4), ZN => n14);
   U109 : NOR2_X1 port map( A1 => A(6), A2 => n11, ZN => n9);
   U110 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n18);
   U111 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n22);
   U112 : NOR2_X1 port map( A1 => A(3), A2 => A(2), ZN => n23);
   U113 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => n4);
   U114 : INV_X1 port map( A => A(8), ZN => n8);
   U115 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n35);
   U116 : NOR2_X1 port map( A1 => A(27), A2 => A(26), ZN => n45);
   U117 : NOR2_X1 port map( A1 => A(25), A2 => A(24), ZN => n44);
   U118 : NAND2_X1 port map( A1 => n15, A2 => n19, ZN => n16);
   U119 : INV_X1 port map( A => A(4), ZN => n19);
   U120 : INV_X1 port map( A => A(28), ZN => n37);
   U121 : INV_X1 port map( A => A(29), ZN => n32);
   U122 : OR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n24);
   U123 : NOR2_X1 port map( A1 => A(2), A2 => n24, ZN => n20);
   U124 : NOR2_X1 port map( A1 => A(28), A2 => A(30), ZN => n26);
   U125 : INV_X1 port map( A => n4, ZN => n1);
   U126 : NAND2_X1 port map( A1 => A(8), A2 => n6, ZN => n5);
   U127 : INV_X1 port map( A => n16, ZN => n12);
   U128 : INV_X1 port map( A => n18, ZN => n15);
   U129 : OAI21_X1 port map( B1 => n31, B2 => n32, A => n30, ZN => SUM(29));
   U130 : INV_X1 port map( A => n38, ZN => n31);
   U131 : OAI21_X1 port map( B1 => n39, B2 => n37, A => n38, ZN => SUM(28));
   U132 : INV_X1 port map( A => n41, ZN => n39);
   U133 : OAI21_X1 port map( B1 => n42, B2 => n43, A => n41, ZN => SUM(27));
   U134 : INV_X1 port map( A => n35, ZN => n27);
   U135 : INV_X1 port map( A => n46, ZN => n42);
   U136 : OAI21_X1 port map( B1 => n47, B2 => n48, A => n46, ZN => SUM(26));
   U137 : INV_X1 port map( A => n50, ZN => n47);
   U138 : OAI21_X1 port map( B1 => n51, B2 => n52, A => n50, ZN => SUM(25));
   U139 : INV_X1 port map( A => n54, ZN => n51);
   U140 : INV_X1 port map( A => n29, ZN => n34);
   U141 : OAI21_X1 port map( B1 => n57, B2 => n58, A => n29, ZN => SUM(23));
   U142 : NAND3_X1 port map( A1 => n63, A2 => n64, A3 => n65, ZN => n62);
   U143 : INV_X1 port map( A => n66, ZN => n57);
   U144 : INV_X1 port map( A => n71, ZN => n67);
   U145 : INV_X1 port map( A => n74, ZN => n72);
   U146 : INV_X1 port map( A => n76, ZN => n70);
   U147 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n77);
   U148 : OAI21_X1 port map( B1 => n78, B2 => n79, A => n76, ZN => SUM(19));
   U149 : INV_X1 port map( A => n61, ZN => n80);
   U150 : INV_X1 port map( A => n83, ZN => n78);
   U151 : INV_X1 port map( A => n89, ZN => n86);
   U152 : INV_X1 port map( A => n91, ZN => n60);
   U153 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n98);
   U154 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => n97);
   U155 : NAND2_X1 port map( A1 => n105, A2 => n106, ZN => n104);
   U156 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => n103);
   U157 : INV_X1 port map( A => n114, ZN => n110);
   U158 : INV_X1 port map( A => n116, ZN => n113);
   U159 : OAI21_X1 port map( B1 => n118, B2 => n119, A => n116, ZN => SUM(11));
   U160 : INV_X1 port map( A => n123, ZN => n118);
   U161 : INV_X1 port map( A => n6, ZN => n7);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_0_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_adder_0_DW01_add_1;

architecture SYN_cla of PC_adder_0_DW01_add_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => n199, A2 => n200, ZN => n1);
   U3 : AND3_X1 port map( A1 => n51, A2 => n52, A3 => n53, ZN => n2);
   U4 : AND2_X1 port map( A1 => n153, A2 => n154, ZN => n3);
   U5 : AND2_X1 port map( A1 => n108, A2 => n109, ZN => n4);
   U6 : AND2_X1 port map( A1 => n210, A2 => n211, ZN => n5);
   U7 : INV_X1 port map( A => n1, ZN => n6);
   U8 : INV_X1 port map( A => n1, ZN => n7);
   U9 : OR2_X2 port map( A1 => B(8), A2 => A(8), ZN => n22);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => n26);
   U11 : NOR2_X1 port map( A1 => n49, A2 => n236, ZN => n8);
   U12 : OR2_X1 port map( A1 => n282, A2 => n283, ZN => n9);
   U13 : AND2_X1 port map( A1 => n184, A2 => n289, ZN => SUM(0));
   U14 : NOR2_X1 port map( A1 => n122, A2 => n123, ZN => n119);
   U15 : NOR2_X1 port map( A1 => n124, A2 => n125, ZN => n123);
   U16 : INV_X1 port map( A => n121, ZN => n126);
   U17 : NAND2_X1 port map( A1 => n140, A2 => n141, ZN => n132);
   U18 : AND2_X1 port map( A1 => n113, A2 => n127, ZN => n140);
   U19 : INV_X1 port map( A => n125, ZN => n142);
   U20 : AND2_X1 port map( A1 => n116, A2 => n13, ZN => n11);
   U21 : NAND2_X1 port map( A1 => n11, A2 => n14, ZN => n69);
   U22 : NAND2_X1 port map( A1 => n116, A2 => n13, ZN => n125);
   U23 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n21);
   U24 : NAND2_X1 port map( A1 => n143, A2 => n13, ZN => n127);
   U25 : NAND2_X1 port map( A1 => n14, A2 => n93, ZN => n72);
   U26 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n73);
   U27 : NOR2_X1 port map( A1 => n230, A2 => n231, ZN => n214);
   U28 : NAND2_X1 port map( A1 => n227, A2 => n228, ZN => n231);
   U29 : AOI21_X1 port map( B1 => n201, B2 => n202, A => n203, ZN => n200);
   U30 : NOR2_X1 port map( A1 => n214, A2 => n215, ZN => n199);
   U31 : AOI21_X1 port map( B1 => n193, B2 => n175, A => n194, ZN => n192);
   U32 : NAND2_X1 port map( A1 => n175, A2 => n182, ZN => n191);
   U33 : NAND2_X1 port map( A1 => n114, A2 => n180, ZN => n185);
   U34 : NOR2_X1 port map( A1 => n67, A2 => n68, ZN => n62);
   U35 : NOR2_X1 port map( A1 => n124, A2 => n69, ZN => n68);
   U36 : XNOR2_X1 port map( A => n117, B => n118, ZN => SUM(27));
   U37 : NAND2_X1 port map( A1 => n92, A2 => n102, ZN => n118);
   U38 : OAI21_X1 port map( B1 => n119, B2 => n120, A => n103, ZN => n117);
   U39 : OAI21_X1 port map( B1 => n121, B2 => n15, A => n105, ZN => n120);
   U40 : NAND2_X1 port map( A1 => n146, A2 => n152, ZN => n162);
   U41 : NAND2_X1 port map( A1 => n168, A2 => n169, ZN => n166);
   U42 : AND2_X1 port map( A1 => n154, A2 => n161, ZN => n168);
   U43 : XNOR2_X1 port map( A => n128, B => n129, ZN => SUM(26));
   U44 : NOR2_X1 port map( A1 => n130, A2 => n131, ZN => n129);
   U45 : AOI21_X1 port map( B1 => n15, B2 => n132, A => n121, ZN => n128);
   U46 : XNOR2_X1 port map( A => n134, B => n135, ZN => SUM(25));
   U47 : NOR2_X1 port map( A1 => n136, A2 => n137, ZN => n135);
   U48 : AOI21_X1 port map( B1 => n132, B2 => n110, A => n138, ZN => n134);
   U49 : NAND2_X1 port map( A1 => n147, A2 => n151, ZN => n156);
   U50 : AND3_X1 port map( A1 => n7, A2 => n116, A3 => n144, ZN => n12);
   U51 : XNOR2_X1 port map( A => n96, B => n97, ZN => SUM(28));
   U52 : NAND2_X1 port map( A1 => n87, A2 => n90, ZN => n96);
   U53 : OAI21_X1 port map( B1 => n98, B2 => n95, A => n99, ZN => n97);
   U54 : NAND2_X1 port map( A1 => n66, A2 => n71, ZN => n84);
   U55 : NAND2_X1 port map( A1 => n176, A2 => n181, ZN => n190);
   U56 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => n139);
   U57 : NAND4_X1 port map( A1 => n182, A2 => n175, A3 => n176, A4 => n114, ZN 
                           => n160);
   U58 : NAND2_X1 port map( A1 => n144, A2 => n154, ZN => n171);
   U59 : NAND2_X1 port map( A1 => n175, A2 => n178, ZN => n195);
   U60 : NAND2_X1 port map( A1 => n145, A2 => n153, ZN => n167);
   U61 : AND4_X1 port map( A1 => n144, A2 => n145, A3 => n146, A4 => n147, ZN 
                           => n13);
   U62 : NAND4_X1 port map( A1 => n110, A2 => n111, A3 => n105, A4 => n92, ZN 
                           => n95);
   U63 : AND2_X1 port map( A1 => n94, A2 => n87, ZN => n14);
   U64 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => n111);
   U65 : INV_X1 port map( A => A(25), ZN => n106);
   U66 : XNOR2_X1 port map( A => n237, B => n238, ZN => SUM(15));
   U67 : NAND2_X1 port map( A1 => n220, A2 => n226, ZN => n238);
   U68 : NAND2_X1 port map( A1 => n242, A2 => n225, ZN => n239);
   U69 : NAND2_X1 port map( A1 => n250, A2 => n251, ZN => n246);
   U70 : AOI21_X1 port map( B1 => n213, B2 => n252, A => n253, ZN => n250);
   U71 : NAND2_X1 port map( A1 => n246, A2 => n247, ZN => n241);
   U72 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n198);
   U73 : XNOR2_X1 port map( A => n268, B => n269, ZN => SUM(11));
   U74 : NAND2_X1 port map( A1 => n208, A2 => n266, ZN => n268);
   U75 : NAND2_X1 port map( A1 => n270, A2 => n267, ZN => n269);
   U76 : OAI21_X1 port map( B1 => n271, B2 => n272, A => n273, ZN => n270);
   U77 : NAND2_X1 port map( A1 => n281, A2 => n22, ZN => n276);
   U78 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n281);
   U79 : XNOR2_X1 port map( A => n277, B => n278, ZN => SUM(10));
   U80 : NAND2_X1 port map( A1 => n267, A2 => n274, ZN => n277);
   U81 : NAND2_X1 port map( A1 => n279, A2 => n20, ZN => n278);
   U82 : NAND2_X1 port map( A1 => n280, A2 => n275, ZN => n279);
   U83 : NAND2_X1 port map( A1 => n276, A2 => n24, ZN => n280);
   U84 : AND2_X1 port map( A1 => n50, A2 => n53, ZN => n235);
   U85 : NAND4_X1 port map( A1 => n47, A2 => n41, A3 => n33, A4 => n36, ZN => 
                           n236);
   U86 : NAND2_X1 port map( A1 => n290, A2 => n291, ZN => n33);
   U87 : INV_X1 port map( A => A(6), ZN => n291);
   U88 : NAND2_X1 port map( A1 => n225, A2 => n223, ZN => n243);
   U89 : OAI21_X1 port map( B1 => n245, B2 => n221, A => n224, ZN => n244);
   U90 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM(7));
   U91 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => n29);
   U92 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => n30);
   U93 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => n32);
   U94 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n42);
   U95 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => n44);
   U96 : OAI21_X1 port map( B1 => n38, B2 => n39, A => n40, ZN => n34);
   U97 : OAI21_X1 port map( B1 => n2, B2 => n49, A => n50, ZN => n46);
   U98 : NAND2_X1 port map( A1 => n292, A2 => n293, ZN => n41);
   U99 : INV_X1 port map( A => A(5), ZN => n293);
   U100 : XNOR2_X1 port map( A => n248, B => n249, ZN => SUM(13));
   U101 : NAND2_X1 port map( A1 => n233, A2 => n224, ZN => n248);
   U102 : NAND2_X1 port map( A1 => n246, A2 => n247, ZN => n249);
   U103 : AND2_X1 port map( A1 => n110, A2 => n111, ZN => n15);
   U104 : XNOR2_X1 port map( A => n37, B => n34, ZN => SUM(6));
   U105 : NAND2_X1 port map( A1 => n33, A2 => n31, ZN => n37);
   U106 : AOI21_X1 port map( B1 => n25, B2 => n26, A => n213, ZN => n258);
   U107 : XNOR2_X1 port map( A => n254, B => n255, ZN => SUM(12));
   U108 : NOR2_X1 port map( A1 => n253, A2 => n256, ZN => n255);
   U109 : NOR2_X1 port map( A1 => n257, A2 => n258, ZN => n254);
   U110 : XNOR2_X1 port map( A => n16, B => n17, ZN => SUM(9));
   U111 : NOR2_X1 port map( A1 => n18, A2 => n19, ZN => n17);
   U112 : AOI21_X1 port map( B1 => n21, B2 => n22, A => n23, ZN => n16);
   U113 : XNOR2_X1 port map( A => n27, B => n28, ZN => SUM(8));
   U114 : NAND2_X1 port map( A1 => n24, A2 => n22, ZN => n27);
   U115 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n28);
   U116 : AND2_X1 port map( A1 => n145, A2 => n146, ZN => n159);
   U117 : XNOR2_X1 port map( A => n43, B => n42, ZN => SUM(5));
   U118 : NAND2_X1 port map( A1 => n41, A2 => n40, ZN => n43);
   U119 : NAND2_X1 port map( A1 => n45, A2 => n47, ZN => n48);
   U120 : NAND2_X1 port map( A1 => n59, A2 => n50, ZN => n54);
   U121 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n58);
   U122 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n79);
   U123 : INV_X1 port map( A => n184, ZN => n82);
   U124 : XNOR2_X1 port map( A => n78, B => n58, ZN => SUM(2));
   U125 : NAND2_X1 port map( A1 => n83, A2 => n53, ZN => n78);
   U126 : XNOR2_X1 port map( A => n183, B => n82, ZN => SUM(1));
   U127 : NAND2_X1 port map( A1 => n81, A2 => n80, ZN => n183);
   U128 : OAI21_X1 port map( B1 => n265, B2 => n207, A => n208, ZN => n252);
   U129 : AOI21_X1 port map( B1 => n20, B2 => n24, A => n209, ZN => n265);
   U130 : AND2_X1 port map( A1 => n212, A2 => n36, ZN => n202);
   U131 : OAI21_X1 port map( B1 => n206, B2 => n207, A => n208, ZN => n205);
   U132 : NOR2_X1 port map( A1 => n5, A2 => n209, ZN => n206);
   U133 : NAND2_X1 port map( A1 => n36, A2 => n212, ZN => n25);
   U134 : AND2_X1 port map( A1 => n226, A2 => n225, ZN => n217);
   U135 : OAI21_X1 port map( B1 => n4, B2 => n100, A => n101, ZN => n91);
   U136 : AND2_X1 port map( A1 => n102, A2 => n103, ZN => n101);
   U137 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => n100);
   U138 : AND2_X1 port map( A1 => n133, A2 => n111, ZN => n121);
   U139 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => n133);
   U140 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => n113);
   U141 : OAI21_X1 port map( B1 => n3, B2 => n149, A => n150, ZN => n148);
   U142 : AND2_X1 port map( A1 => n151, A2 => n152, ZN => n150);
   U143 : NAND2_X1 port map( A1 => n266, A2 => n267, ZN => n207);
   U144 : NAND2_X1 port map( A1 => n294, A2 => n295, ZN => n212);
   U145 : NOR2_X1 port map( A1 => n299, A2 => n300, ZN => n294);
   U146 : NAND2_X1 port map( A1 => n35, A2 => n31, ZN => n299);
   U147 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => n93);
   U148 : NAND2_X1 port map( A1 => n173, A2 => n174, ZN => n115);
   U149 : AND2_X1 port map( A1 => n180, A2 => n181, ZN => n173);
   U150 : NAND2_X1 port map( A1 => n178, A2 => n179, ZN => n177);
   U151 : NAND2_X1 port map( A1 => n51, A2 => n288, ZN => n282);
   U152 : AND2_X1 port map( A1 => n50, A2 => n53, ZN => n288);
   U153 : NAND2_X1 port map( A1 => n143, A2 => n144, ZN => n161);
   U154 : NAND2_X1 port map( A1 => n20, A2 => n24, ZN => n272);
   U155 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => n170);
   U156 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => n70);
   U157 : NAND2_X1 port map( A1 => n145, A2 => n146, ZN => n149);
   U158 : INV_X1 port map( A => A(0), ZN => n304);
   U159 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => n104);
   U160 : NAND2_X1 port map( A1 => n290, A2 => n291, ZN => n297);
   U161 : NAND2_X1 port map( A1 => n292, A2 => n293, ZN => n296);
   U162 : INV_X1 port map( A => n216, ZN => n215);
   U163 : AOI21_X1 port map( B1 => n217, B2 => n218, A => n219, ZN => n216);
   U164 : OAI211_X1 port map( C1 => n221, C2 => n222, A => n223, B => n224, ZN 
                           => n218);
   U165 : OR2_X1 port map( A1 => B(14), A2 => A(14), ZN => n225);
   U166 : XNOR2_X1 port map( A => n60, B => n61, ZN => SUM(31));
   U167 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n61);
   U168 : OAI21_X1 port map( B1 => n62, B2 => n63, A => n64, ZN => n60);
   U169 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => n63);
   U170 : OR2_X1 port map( A1 => B(13), A2 => A(13), ZN => n233);
   U171 : OR2_X1 port map( A1 => B(15), A2 => A(15), ZN => n226);
   U172 : OR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n232);
   U173 : OR2_X1 port map( A1 => B(17), A2 => A(17), ZN => n175);
   U174 : OR2_X1 port map( A1 => B(19), A2 => A(19), ZN => n114);
   U175 : OR2_X1 port map( A1 => B(21), A2 => A(21), ZN => n145);
   U176 : OR2_X1 port map( A1 => B(22), A2 => A(22), ZN => n146);
   U177 : OR2_X1 port map( A1 => B(23), A2 => A(23), ZN => n147);
   U178 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n176);
   U179 : OR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n144);
   U180 : OR2_X1 port map( A1 => B(16), A2 => A(16), ZN => n182);
   U181 : OR2_X1 port map( A1 => B(27), A2 => A(27), ZN => n92);
   U182 : OR2_X1 port map( A1 => B(26), A2 => A(26), ZN => n105);
   U183 : OR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n110);
   U184 : NAND2_X1 port map( A1 => n259, A2 => n260, ZN => n213);
   U185 : NOR2_X1 port map( A1 => A(9), A2 => B(9), ZN => n264);
   U186 : OR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n274);
   U187 : OR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n208);
   U188 : NOR2_X1 port map( A1 => A(1), A2 => B(1), ZN => n287);
   U189 : NAND2_X1 port map( A1 => n284, A2 => n285, ZN => n52);
   U190 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n284);
   U191 : NOR2_X1 port map( A1 => n286, A2 => n287, ZN => n285);
   U192 : NOR2_X1 port map( A1 => A(2), A2 => B(2), ZN => n286);
   U193 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n36);
   U194 : OR2_X1 port map( A1 => B(28), A2 => A(28), ZN => n87);
   U195 : OR2_X1 port map( A1 => B(4), A2 => A(4), ZN => n47);
   U196 : OR2_X1 port map( A1 => B(3), A2 => A(3), ZN => n59);
   U197 : OR2_X1 port map( A1 => B(29), A2 => A(29), ZN => n66);
   U198 : OR2_X1 port map( A1 => B(30), A2 => A(30), ZN => n65);
   U199 : OR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n275);
   U200 : OR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n81);
   U201 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n184);
   U202 : OR2_X1 port map( A1 => B(2), A2 => A(2), ZN => n83);
   U203 : NAND2_X1 port map( A1 => n303, A2 => n304, ZN => n289);
   U204 : INV_X1 port map( A => B(0), ZN => n303);
   U205 : OAI22_X1 port map( A1 => A(10), A2 => B(10), B1 => A(9), B2 => B(9), 
                           ZN => n209);
   U206 : OAI211_X1 port map( C1 => A(2), C2 => B(2), A => A(1), B => B(1), ZN 
                           => n51);
   U207 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n24);
   U208 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n20);
   U209 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n109);
   U210 : NAND2_X1 port map( A1 => B(13), A2 => A(13), ZN => n224);
   U211 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n53);
   U212 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n179);
   U213 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n154);
   U214 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n50);
   U215 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n31);
   U216 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n267);
   U217 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n153);
   U218 : NAND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n247);
   U219 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n223);
   U220 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n178);
   U221 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n108);
   U222 : NOR2_X1 port map( A1 => n301, A2 => n302, ZN => n300);
   U223 : NOR2_X1 port map( A1 => A(6), A2 => B(6), ZN => n301);
   U224 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n80);
   U225 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n181);
   U226 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n152);
   U227 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n71);
   U228 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => n103);
   U229 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n40);
   U230 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n45);
   U231 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n266);
   U232 : NAND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n64);
   U233 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n35);
   U234 : NAND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n90);
   U235 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n180);
   U236 : NAND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n151);
   U237 : NAND2_X1 port map( A1 => B(27), A2 => A(27), ZN => n102);
   U238 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n220);
   U239 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n298);
   U240 : INV_X1 port map( A => B(25), ZN => n107);
   U241 : INV_X1 port map( A => B(6), ZN => n290);
   U242 : INV_X1 port map( A => B(5), ZN => n292);
   U243 : NOR2_X1 port map( A1 => n204, A2 => n213, ZN => n201);
   U244 : NOR2_X1 port map( A1 => n204, A2 => n205, ZN => n203);
   U245 : NAND4_X1 port map( A1 => n232, A2 => n233, A3 => n225, A4 => n226, ZN
                           => n204);
   U246 : XNOR2_X1 port map( A => n155, B => n156, ZN => SUM(23));
   U247 : NAND2_X1 port map( A1 => n152, A2 => n157, ZN => n155);
   U248 : OAI21_X1 port map( B1 => n158, B2 => n12, A => n159, ZN => n157);
   U249 : XNOR2_X1 port map( A => n7, B => n198, ZN => SUM(16));
   U250 : OAI21_X1 port map( B1 => n85, B2 => n191, A => n192, ZN => n189);
   U251 : AOI21_X1 port map( B1 => n7, B2 => n11, A => n93, ZN => n98);
   U252 : OAI211_X1 port map( C1 => n85, C2 => n69, A => n72, B => n70, ZN => 
                           n77);
   U253 : NAND2_X1 port map( A1 => n7, A2 => n142, ZN => n141);
   U254 : INV_X1 port map( A => n7, ZN => n124);
   U255 : INV_X1 port map( A => n20, ZN => n18);
   U256 : INV_X1 port map( A => n24, ZN => n23);
   U257 : INV_X1 port map( A => n41, ZN => n39);
   U258 : INV_X1 port map( A => n42, ZN => n38);
   U259 : XNOR2_X1 port map( A => n48, B => n46, ZN => SUM(4));
   U260 : XNOR2_X1 port map( A => n54, B => n55, ZN => SUM(3));
   U261 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n53, ZN => n55);
   U262 : INV_X1 port map( A => n58, ZN => n56);
   U263 : NAND3_X1 port map( A1 => n70, A2 => n71, A3 => n72, ZN => n67);
   U264 : XNOR2_X1 port map( A => n74, B => n73, ZN => SUM(30));
   U265 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n71, ZN => n74);
   U266 : INV_X1 port map( A => n66, ZN => n76);
   U267 : INV_X1 port map( A => n77, ZN => n75);
   U268 : XNOR2_X1 port map( A => n77, B => n84, ZN => SUM(29));
   U269 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n86);
   U270 : INV_X1 port map( A => n91, ZN => n89);
   U271 : INV_X1 port map( A => n92, ZN => n88);
   U272 : INV_X1 port map( A => n95, ZN => n94);
   U273 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => n99);
   U274 : NAND3_X1 port map( A1 => n13, A2 => n114, A3 => n115, ZN => n112);
   U275 : NAND3_X1 port map( A1 => n126, A2 => n113, A3 => n127, ZN => n122);
   U276 : INV_X1 port map( A => n105, ZN => n131);
   U277 : INV_X1 port map( A => n103, ZN => n130);
   U278 : INV_X1 port map( A => n111, ZN => n137);
   U279 : INV_X1 port map( A => n108, ZN => n136);
   U280 : INV_X1 port map( A => n109, ZN => n138);
   U281 : XNOR2_X1 port map( A => n139, B => n132, ZN => SUM(24));
   U282 : NAND3_X1 port map( A1 => n153, A2 => n154, A3 => n161, ZN => n158);
   U283 : XNOR2_X1 port map( A => n163, B => n162, ZN => SUM(22));
   U284 : OAI21_X1 port map( B1 => n164, B2 => n165, A => n153, ZN => n163);
   U285 : INV_X1 port map( A => n145, ZN => n165);
   U286 : INV_X1 port map( A => n166, ZN => n164);
   U287 : XNOR2_X1 port map( A => n167, B => n166, ZN => SUM(21));
   U288 : NAND3_X1 port map( A1 => n7, A2 => n116, A3 => n144, ZN => n169);
   U289 : INV_X1 port map( A => n160, ZN => n116);
   U290 : INV_X1 port map( A => n170, ZN => n143);
   U291 : XNOR2_X1 port map( A => n171, B => n172, ZN => SUM(20));
   U292 : OAI21_X1 port map( B1 => n85, B2 => n160, A => n170, ZN => n172);
   U293 : NAND3_X1 port map( A1 => n175, A2 => n176, A3 => n177, ZN => n174);
   U294 : XNOR2_X1 port map( A => n185, B => n186, ZN => SUM(19));
   U295 : OAI21_X1 port map( B1 => n187, B2 => n188, A => n181, ZN => n186);
   U296 : INV_X1 port map( A => n176, ZN => n188);
   U297 : INV_X1 port map( A => n189, ZN => n187);
   U298 : XNOR2_X1 port map( A => n190, B => n189, ZN => SUM(18));
   U299 : INV_X1 port map( A => n178, ZN => n194);
   U300 : INV_X1 port map( A => n179, ZN => n193);
   U301 : XNOR2_X1 port map( A => n195, B => n196, ZN => SUM(17));
   U302 : OAI21_X1 port map( B1 => n85, B2 => n197, A => n179, ZN => n196);
   U303 : INV_X1 port map( A => n182, ZN => n197);
   U304 : INV_X1 port map( A => n6, ZN => n85);
   U305 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n211);
   U306 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n210);
   U307 : INV_X1 port map( A => n220, ZN => n219);
   U308 : NAND2_X1 port map( A1 => A(12), A2 => B(12), ZN => n222);
   U309 : INV_X1 port map( A => n204, ZN => n228);
   U310 : INV_X1 port map( A => n213, ZN => n227);
   U311 : NAND3_X1 port map( A1 => n229, A2 => n59, A3 => n234, ZN => n230);
   U312 : NAND3_X1 port map( A1 => n51, A2 => n235, A3 => n52, ZN => n234);
   U313 : INV_X1 port map( A => n236, ZN => n229);
   U314 : NAND3_X1 port map( A1 => n223, A2 => n239, A3 => n240, ZN => n237);
   U315 : NAND3_X1 port map( A1 => n233, A2 => n225, A3 => n241, ZN => n240);
   U316 : INV_X1 port map( A => n224, ZN => n242);
   U317 : XNOR2_X1 port map( A => n243, B => n244, ZN => SUM(14));
   U318 : INV_X1 port map( A => n233, ZN => n221);
   U319 : INV_X1 port map( A => n241, ZN => n245);
   U320 : NAND3_X1 port map( A1 => n25, A2 => n252, A3 => n26, ZN => n251);
   U321 : INV_X1 port map( A => n247, ZN => n256);
   U322 : INV_X1 port map( A => n232, ZN => n253);
   U323 : NOR2_X1 port map( A1 => n261, A2 => n262, ZN => n260);
   U324 : INV_X1 port map( A => n22, ZN => n261);
   U325 : NOR2_X1 port map( A1 => n263, A2 => n264, ZN => n259);
   U326 : INV_X1 port map( A => n208, ZN => n263);
   U327 : INV_X1 port map( A => n252, ZN => n257);
   U328 : NOR2_X1 port map( A1 => n19, A2 => n262, ZN => n273);
   U329 : INV_X1 port map( A => n274, ZN => n262);
   U330 : INV_X1 port map( A => n275, ZN => n19);
   U331 : INV_X1 port map( A => n276, ZN => n271);
   U332 : INV_X1 port map( A => n52, ZN => n283);
   U333 : INV_X1 port map( A => n83, ZN => n57);
   U334 : INV_X1 port map( A => n59, ZN => n49);
   U335 : NAND3_X1 port map( A1 => n296, A2 => n297, A3 => n298, ZN => n295);
   U336 : NAND2_X1 port map( A1 => A(5), A2 => B(5), ZN => n302);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_1_DW01_add_0_DW01_add_128 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_adder_1_DW01_add_0_DW01_add_128;

architecture SYN_rpl of PC_adder_1_DW01_add_0_DW01_add_128 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1005 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1005, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_63;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_63 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_62;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : AOI22_X1 port map( A1 => B(3), A2 => SEL, B1 => A(3), B2 => n1, ZN => 
                           n2);
   U6 : INV_X1 port map( A => n2, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_61;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_61 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U5 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_60;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_60 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_59;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_59 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_58;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_58 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_57;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_57 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_56;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_55;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_54;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_53;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_52;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_51;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_50;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_49;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_48;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_48 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_47;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_47 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_46;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_46 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_45;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_45 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_44;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_44 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_43;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_43 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_42;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_42 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_41;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_41 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_40;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_40 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_39;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_39 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_38;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_38 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_37;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_37 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_36;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_36 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_35;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_35 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_34;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_34 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => A(3), ZN => n2);
   U2 : NAND2_X1 port map( A1 => B(3), A2 => SEL, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(3));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U6 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U7 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_33;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_33 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_32;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_31;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_30;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_29;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_28;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_27;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_26;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_25;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_24;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_23;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_22;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_21;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_20;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_19;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_18;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_17;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_16;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_15;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_14;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_13;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_12;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_11;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_10;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_9;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_8;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_7;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_6;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_5;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_4;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_3;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : AOI22_X1 port map( A1 => B(3), A2 => SEL, B1 => A(3), B2 => n1, ZN => 
                           n2);
   U6 : INV_X1 port map( A => n2, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_2;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : AOI22_X1 port map( A1 => B(3), A2 => SEL, B1 => A(3), B2 => n1, ZN => 
                           n2);
   U6 : INV_X1 port map( A => n2, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_1;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_127 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_127;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_127 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n17, B => n16, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n13);
   U4 : XNOR2_X1 port map( A => n14, B => n13, ZN => S(2));
   U5 : XNOR2_X1 port map( A => n12, B => n11, ZN => S(1));
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U9 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n14);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U12 : INV_X1 port map( A => A(3), ZN => n15);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : INV_X1 port map( A => A(2), ZN => n7);
   U15 : INV_X1 port map( A => B(2), ZN => n6);
   U16 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n5);
   U17 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n5, ZN => n16);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n15, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U21 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U22 : XOR2_X1 port map( A => n15, B => B(3), Z => n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_126 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_126;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_126 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n_1006 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A(3), ZN => n11);
   U2 : INV_X1 port map( A => B(3), ZN => n10);
   U3 : INV_X1 port map( A => A(2), ZN => n8);
   U4 : INV_X1 port map( A => B(2), ZN => n7);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n16);
   U6 : INV_X1 port map( A => n16, ZN => n5);
   U7 : INV_X1 port map( A => A(0), ZN => n3);
   U8 : INV_X1 port map( A => B(0), ZN => n2);
   U9 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n1);
   U10 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => n13);
   U11 : INV_X1 port map( A => A(1), ZN => n12);
   U12 : INV_X1 port map( A => B(1), ZN => n4);
   U13 : NAND2_X1 port map( A1 => n12, A2 => n4, ZN => n15);
   U14 : OAI221_X1 port map( B1 => B(2), B2 => A(2), C1 => n5, C2 => n13, A => 
                           n15, ZN => n6);
   U15 : OAI21_X1 port map( B1 => n8, B2 => n7, A => n6, ZN => n21);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n21, ZN => n9);
   U17 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => Co);
   U18 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1006, S => 
                           S(0));
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n13, ZN => n17);
   U21 : XOR2_X1 port map( A => n14, B => n17, Z => S(1));
   U22 : INV_X1 port map( A => n15, ZN => n18);
   U23 : OAI21_X1 port map( B1 => n18, B2 => n17, A => n16, ZN => n20);
   U24 : XOR2_X1 port map( A => B(2), B => A(2), Z => n19);
   U25 : XOR2_X1 port map( A => n20, B => n19, Z => S(2));
   U26 : XOR2_X1 port map( A => n21, B => A(3), Z => n22);
   U27 : XOR2_X1 port map( A => n22, B => B(3), Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_125 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_125;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_125 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n_1007 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n10);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : INV_X1 port map( A => A(3), ZN => n17);
   U5 : INV_X1 port map( A => B(3), ZN => n8);
   U6 : INV_X1 port map( A => A(2), ZN => n13);
   U7 : INV_X1 port map( A => B(2), ZN => n6);
   U8 : INV_X1 port map( A => A(1), ZN => n9);
   U9 : INV_X1 port map( A => B(1), ZN => n4);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n10, ZN => n3);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n4, A => n3, ZN => n14);
   U12 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n5);
   U13 : OAI21_X1 port map( B1 => n13, B2 => n6, A => n5, ZN => n18);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n17, B2 => n8, A => n7, ZN => Co);
   U16 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1007, S => 
                           S(0));
   U17 : XOR2_X1 port map( A => n9, B => B(1), Z => n12);
   U18 : INV_X1 port map( A => n10, ZN => n11);
   U19 : XOR2_X1 port map( A => n12, B => n11, Z => S(1));
   U20 : XOR2_X1 port map( A => n13, B => B(2), Z => n16);
   U21 : INV_X1 port map( A => n14, ZN => n15);
   U22 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));
   U23 : XOR2_X1 port map( A => n17, B => B(3), Z => n20);
   U24 : INV_X1 port map( A => n18, ZN => n19);
   U25 : XOR2_X1 port map( A => n20, B => n19, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_124 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_124;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_124 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U2 : INV_X1 port map( A => n22, ZN => n9);
   U3 : INV_X1 port map( A => n19, ZN => n3);
   U4 : OR2_X1 port map( A1 => A(2), A2 => B(2), ZN => n8);
   U5 : NAND4_X1 port map( A1 => n13, A2 => n12, A3 => n11, A4 => n10, ZN => 
                           n26);
   U6 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n13);
   U7 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n10);
   U8 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n27);
   U9 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n11);
   U10 : INV_X1 port map( A => n20, ZN => n6);
   U11 : NOR2_X1 port map( A1 => n23, A2 => n5, ZN => n7);
   U12 : AND2_X1 port map( A1 => n20, A2 => n19, ZN => n1);
   U13 : INV_X1 port map( A => A(3), ZN => n16);
   U14 : INV_X1 port map( A => B(3), ZN => n15);
   U15 : INV_X1 port map( A => A(1), ZN => n18);
   U16 : INV_X1 port map( A => B(1), ZN => n2);
   U17 : NAND2_X1 port map( A1 => n18, A2 => n2, ZN => n4);
   U18 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n19);
   U19 : NAND3_X1 port map( A1 => n4, A2 => n3, A3 => n8, ZN => n12);
   U20 : INV_X1 port map( A => n4, ZN => n23);
   U21 : INV_X1 port map( A => n8, ZN => n5);
   U22 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n20);
   U23 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n22);
   U24 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n26, ZN => n14);
   U25 : OAI21_X1 port map( B1 => n16, B2 => n15, A => n14, ZN => Co);
   U26 : XOR2_X1 port map( A => B(0), B => A(0), Z => n17);
   U27 : XOR2_X1 port map( A => Ci, B => n17, Z => S(0));
   U28 : XOR2_X1 port map( A => n18, B => B(1), Z => n21);
   U29 : XOR2_X1 port map( A => n21, B => n1, Z => S(1));
   U30 : OAI21_X1 port map( B1 => n23, B2 => n1, A => n22, ZN => n25);
   U31 : XOR2_X1 port map( A => B(2), B => A(2), Z => n24);
   U32 : XOR2_X1 port map( A => n25, B => n24, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_123 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_123;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_123 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n17, B => n16, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n16);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n6);
   U5 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U6 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n17);
   U7 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U8 : XNOR2_X1 port map( A => n12, B => n11, ZN => S(1));
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n13);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U12 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U15 : INV_X1 port map( A => A(3), ZN => n9);
   U16 : INV_X1 port map( A => B(3), ZN => n8);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n7);
   U18 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U20 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U21 : INV_X1 port map( A => n13, ZN => n14);
   U22 : XOR2_X1 port map( A => n15, B => n14, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_122 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_122;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_122 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n_1008 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n10);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : INV_X1 port map( A => A(3), ZN => n17);
   U5 : INV_X1 port map( A => B(3), ZN => n8);
   U6 : INV_X1 port map( A => A(2), ZN => n13);
   U7 : INV_X1 port map( A => B(2), ZN => n6);
   U8 : INV_X1 port map( A => A(1), ZN => n9);
   U9 : INV_X1 port map( A => B(1), ZN => n4);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n10, ZN => n3);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n4, A => n3, ZN => n14);
   U12 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n5);
   U13 : OAI21_X1 port map( B1 => n13, B2 => n6, A => n5, ZN => n18);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n17, B2 => n8, A => n7, ZN => Co);
   U16 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1008, S => 
                           S(0));
   U17 : XOR2_X1 port map( A => n9, B => B(1), Z => n12);
   U18 : INV_X1 port map( A => n10, ZN => n11);
   U19 : XOR2_X1 port map( A => n12, B => n11, Z => S(1));
   U20 : XOR2_X1 port map( A => n13, B => B(2), Z => n16);
   U21 : INV_X1 port map( A => n14, ZN => n15);
   U22 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));
   U23 : XOR2_X1 port map( A => n17, B => B(3), Z => n20);
   U24 : INV_X1 port map( A => n18, ZN => n19);
   U25 : XOR2_X1 port map( A => n20, B => n19, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_121 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_121;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_121 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n_1009 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n10);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : INV_X1 port map( A => A(3), ZN => n17);
   U5 : INV_X1 port map( A => B(3), ZN => n8);
   U6 : INV_X1 port map( A => A(2), ZN => n13);
   U7 : INV_X1 port map( A => B(2), ZN => n6);
   U8 : INV_X1 port map( A => A(1), ZN => n9);
   U9 : INV_X1 port map( A => B(1), ZN => n4);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n10, ZN => n3);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n4, A => n3, ZN => n14);
   U12 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n5);
   U13 : OAI21_X1 port map( B1 => n13, B2 => n6, A => n5, ZN => n18);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n17, B2 => n8, A => n7, ZN => Co);
   U16 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1009, S => 
                           S(0));
   U17 : XOR2_X1 port map( A => n9, B => B(1), Z => n12);
   U18 : INV_X1 port map( A => n10, ZN => n11);
   U19 : XOR2_X1 port map( A => n12, B => n11, Z => S(1));
   U20 : XOR2_X1 port map( A => n13, B => B(2), Z => n16);
   U21 : INV_X1 port map( A => n14, ZN => n15);
   U22 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));
   U23 : XOR2_X1 port map( A => n17, B => B(3), Z => n20);
   U24 : INV_X1 port map( A => n18, ZN => n19);
   U25 : XOR2_X1 port map( A => n20, B => n19, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_120 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_120;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_120 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U6 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_119 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_119;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_119 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U9 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_118 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_118;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_118 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U3 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U4 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n10, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n10);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : INV_X1 port map( A => A(3), ZN => n17);
   U9 : INV_X1 port map( A => B(3), ZN => n8);
   U10 : INV_X1 port map( A => A(2), ZN => n13);
   U11 : INV_X1 port map( A => B(2), ZN => n6);
   U12 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n5);
   U13 : OAI21_X1 port map( B1 => n13, B2 => n6, A => n5, ZN => n18);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n17, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n9);
   U17 : XOR2_X1 port map( A => Ci, B => n9, Z => S(0));
   U18 : INV_X1 port map( A => n10, ZN => n11);
   U19 : XOR2_X1 port map( A => n12, B => n11, Z => S(1));
   U20 : XOR2_X1 port map( A => n13, B => B(2), Z => n16);
   U21 : INV_X1 port map( A => n14, ZN => n15);
   U22 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));
   U23 : XOR2_X1 port map( A => n17, B => B(3), Z => n20);
   U24 : INV_X1 port map( A => n18, ZN => n19);
   U25 : XOR2_X1 port map( A => n20, B => n19, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_117 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_117;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_117 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n15);
   U2 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U3 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U5 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U6 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U7 : INV_X1 port map( A => A(3), ZN => n18);
   U8 : INV_X1 port map( A => B(3), ZN => n8);
   U9 : INV_X1 port map( A => A(2), ZN => n14);
   U10 : INV_X1 port map( A => B(2), ZN => n6);
   U11 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n15, ZN => n5);
   U12 : OAI21_X1 port map( B1 => n14, B2 => n6, A => n5, ZN => n19);
   U13 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U14 : OAI21_X1 port map( B1 => n18, B2 => n8, A => n7, ZN => Co);
   U15 : XOR2_X1 port map( A => B(0), B => A(0), Z => n9);
   U16 : XOR2_X1 port map( A => Ci, B => n9, Z => S(0));
   U17 : INV_X1 port map( A => A(1), ZN => n10);
   U18 : XOR2_X1 port map( A => n10, B => B(1), Z => n13);
   U19 : INV_X1 port map( A => n11, ZN => n12);
   U20 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U21 : XOR2_X1 port map( A => n14, B => B(2), Z => n17);
   U22 : INV_X1 port map( A => n15, ZN => n16);
   U23 : XOR2_X1 port map( A => n17, B => n16, Z => S(2));
   U24 : XOR2_X1 port map( A => n18, B => B(3), Z => n21);
   U25 : INV_X1 port map( A => n19, ZN => n20);
   U26 : XOR2_X1 port map( A => n21, B => n20, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_116 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_116;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_116 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U6 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_115 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_115;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_115 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U6 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U7 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U8 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U9 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U10 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U11 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_114 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_114;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_114 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U2 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n15);
   U3 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U8 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U9 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U10 : INV_X1 port map( A => A(3), ZN => n16);
   U11 : INV_X1 port map( A => B(3), ZN => n9);
   U12 : INV_X1 port map( A => A(2), ZN => n7);
   U13 : INV_X1 port map( A => B(2), ZN => n6);
   U14 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n5);
   U15 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n5, ZN => n17);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n8);
   U17 : OAI21_X1 port map( B1 => n16, B2 => n9, A => n8, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : XOR2_X1 port map( A => n16, B => B(3), Z => n19);
   U23 : INV_X1 port map( A => n17, ZN => n18);
   U24 : XOR2_X1 port map( A => n19, B => n18, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_113 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_113;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_113 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n16, B => n15, ZN => S(2));
   U2 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n16);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n15);
   U4 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U5 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : INV_X1 port map( A => A(3), ZN => n17);
   U10 : INV_X1 port map( A => B(3), ZN => n9);
   U11 : INV_X1 port map( A => A(2), ZN => n7);
   U12 : INV_X1 port map( A => B(2), ZN => n6);
   U13 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n15, ZN => n5);
   U14 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n5, ZN => n18);
   U15 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n8);
   U16 : OAI21_X1 port map( B1 => n17, B2 => n9, A => n8, ZN => Co);
   U17 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U18 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U19 : INV_X1 port map( A => A(1), ZN => n11);
   U20 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U21 : INV_X1 port map( A => n12, ZN => n13);
   U22 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U23 : XOR2_X1 port map( A => n17, B => B(3), Z => n20);
   U24 : INV_X1 port map( A => n18, ZN => n19);
   U25 : XOR2_X1 port map( A => n20, B => n19, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_112 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_112;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_112 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_111 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_111;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_111 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_110 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_110;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_110 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_109 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_109;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_109 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_108 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_108;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_108 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_107 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_107;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_107 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_106 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_106;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_106 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_105 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_105;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_105 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_104 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_104;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_104 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_103 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_103;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_103 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_102 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_102;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_102 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_101 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_101;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_101 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_100 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_100;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_100 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_99 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_99;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_99 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_98 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_98;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_98 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_97 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_97;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_97 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_96 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_96;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_96 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_95 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_95;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n17, ZN => S(2));
   U2 : XOR2_X1 port map( A => n16, B => B(2), Z => n1);
   U3 : XNOR2_X1 port map( A => n2, B => n18, ZN => S(3));
   U4 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n2);
   U5 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(1));
   U6 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n18);
   U7 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n7);
   U8 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n8);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n4);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U12 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U13 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n5);
   U14 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n14, ZN => n6);
   U15 : INV_X1 port map( A => A(3), ZN => n11);
   U16 : INV_X1 port map( A => B(3), ZN => n10);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n9);
   U18 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n12);
   U20 : XOR2_X1 port map( A => Ci, B => n12, Z => S(0));
   U21 : INV_X1 port map( A => A(1), ZN => n13);
   U22 : XOR2_X1 port map( A => n13, B => B(1), Z => n15);
   U23 : INV_X1 port map( A => A(2), ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_94 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_94;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_94 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_93 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_93;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_93 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_92 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_92;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_92 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_91 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_91;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_91 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_90 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_90;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_90 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_89 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_89;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_89 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_88 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_88;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_88 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_87 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_87;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_87 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_86 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_86;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_86 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_85 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_85;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_85 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_84 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_84;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_84 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_83 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_83;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_83 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_82 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_82;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1010, 
      n_1011, n_1012 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n9);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n10);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n9, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n10, ZN => n6);
   U10 : INV_X1 port map( A => A(3), ZN => n11);
   U11 : INV_X1 port map( A => B(3), ZN => n8);
   U12 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n12, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n11, B2 => n8, A => n7, ZN => Co);
   U14 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1010, S => 
                           S(0));
   U15 : FA_X1 port map( A => A(1), B => B(1), CI => n9, CO => n_1011, S => 
                           S(1));
   U16 : FA_X1 port map( A => A(2), B => B(2), CI => n10, CO => n_1012, S => 
                           S(2));
   U17 : XOR2_X1 port map( A => n11, B => B(3), Z => n14);
   U18 : INV_X1 port map( A => n12, ZN => n13);
   U19 : XOR2_X1 port map( A => n14, B => n13, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_81 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_81;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1013, 
      n_1014, n_1015 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n9);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n10);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n9, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n10, ZN => n6);
   U10 : INV_X1 port map( A => A(3), ZN => n11);
   U11 : INV_X1 port map( A => B(3), ZN => n8);
   U12 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n12, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n11, B2 => n8, A => n7, ZN => Co);
   U14 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1013, S => 
                           S(0));
   U15 : FA_X1 port map( A => A(1), B => B(1), CI => n9, CO => n_1014, S => 
                           S(1));
   U16 : FA_X1 port map( A => A(2), B => B(2), CI => n10, CO => n_1015, S => 
                           S(2));
   U17 : XOR2_X1 port map( A => n11, B => B(3), Z => n14);
   U18 : INV_X1 port map( A => n12, ZN => n13);
   U19 : XOR2_X1 port map( A => n14, B => n13, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_80 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_80;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_80 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_79 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_79;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_79 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n16);
   U2 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U3 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U4 : XOR2_X1 port map( A => n1, B => n19, Z => S(3));
   U5 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U6 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n14);
   U7 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U8 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U9 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U10 : INV_X1 port map( A => A(3), ZN => n10);
   U11 : INV_X1 port map( A => B(3), ZN => n9);
   U12 : INV_X1 port map( A => A(2), ZN => n15);
   U13 : INV_X1 port map( A => B(2), ZN => n7);
   U14 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U15 : OAI21_X1 port map( B1 => n15, B2 => n7, A => n6, ZN => n19);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n8);
   U17 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U19 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U23 : INV_X1 port map( A => n16, ZN => n17);
   U24 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_78 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_78;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_78 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_77 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_77;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_77 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U8 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U9 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_76 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_76;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_76 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_75 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_75;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_74 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_74;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_73 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_73;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_73 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_72 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_72;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_72 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_71 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_71;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_71 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_70 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_70;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_70 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_69 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_69;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_69 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_68 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_68;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_68 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_67 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_67;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_66 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_66;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n12, Z => S(1));
   U2 : XOR2_X1 port map( A => A(1), B => B(1), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n7);
   U6 : XNOR2_X1 port map( A => n17, B => n16, ZN => S(3));
   U7 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n17);
   U8 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n13);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U11 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U12 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U14 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U15 : INV_X1 port map( A => A(3), ZN => n10);
   U16 : INV_X1 port map( A => B(3), ZN => n9);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U18 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U20 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U21 : INV_X1 port map( A => n13, ZN => n14);
   U22 : XOR2_X1 port map( A => n15, B => n14, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_65 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_65;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_65 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U8 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_64 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_64;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_64 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_63;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n17, ZN => S(2));
   U2 : XOR2_X1 port map( A => n16, B => B(2), Z => n1);
   U3 : XNOR2_X1 port map( A => n2, B => n18, ZN => S(3));
   U4 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n2);
   U5 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(1));
   U6 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n18);
   U7 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n7);
   U8 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n8);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n4);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U12 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U13 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n5);
   U14 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n14, ZN => n6);
   U15 : INV_X1 port map( A => A(3), ZN => n11);
   U16 : INV_X1 port map( A => B(3), ZN => n10);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n9);
   U18 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n12);
   U20 : XOR2_X1 port map( A => Ci, B => n12, Z => S(0));
   U21 : INV_X1 port map( A => A(1), ZN => n13);
   U22 : XOR2_X1 port map( A => n13, B => B(1), Z => n15);
   U23 : INV_X1 port map( A => A(2), ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_62;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_61;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_60;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_59;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_58;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_57;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_56;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_55;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_54;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_53;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_52;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_51;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n20, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n20);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U9 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n17);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n8);
   U15 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U17 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n12);
   U19 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U20 : INV_X1 port map( A => n13, ZN => n14);
   U21 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n16);
   U23 : XOR2_X1 port map( A => n16, B => B(2), Z => n19);
   U24 : INV_X1 port map( A => n17, ZN => n18);
   U25 : XOR2_X1 port map( A => n19, B => n18, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_50;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1016, 
      n_1017, n_1018 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n9);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n10);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n9, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n10, ZN => n6);
   U10 : INV_X1 port map( A => A(3), ZN => n11);
   U11 : INV_X1 port map( A => B(3), ZN => n8);
   U12 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n12, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n11, B2 => n8, A => n7, ZN => Co);
   U14 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1016, S => 
                           S(0));
   U15 : FA_X1 port map( A => A(1), B => B(1), CI => n9, CO => n_1017, S => 
                           S(1));
   U16 : FA_X1 port map( A => A(2), B => B(2), CI => n10, CO => n_1018, S => 
                           S(2));
   U17 : XOR2_X1 port map( A => n11, B => B(3), Z => n14);
   U18 : INV_X1 port map( A => n12, ZN => n13);
   U19 : XOR2_X1 port map( A => n14, B => n13, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_49;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1019, 
      n_1020, n_1021 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n9);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n10);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n9, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n10, ZN => n6);
   U10 : INV_X1 port map( A => A(3), ZN => n11);
   U11 : INV_X1 port map( A => B(3), ZN => n8);
   U12 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n12, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n11, B2 => n8, A => n7, ZN => Co);
   U14 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1019, S => 
                           S(0));
   U15 : FA_X1 port map( A => A(1), B => B(1), CI => n9, CO => n_1020, S => 
                           S(1));
   U16 : FA_X1 port map( A => A(2), B => B(2), CI => n10, CO => n_1021, S => 
                           S(2));
   U17 : XOR2_X1 port map( A => n11, B => B(3), Z => n14);
   U18 : INV_X1 port map( A => n12, ZN => n13);
   U19 : XOR2_X1 port map( A => n14, B => n13, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_48;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_48 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_47;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S(0));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => n1);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n6);
   U6 : XOR2_X1 port map( A => n2, B => n19, Z => S(3));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => n2);
   U8 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n14);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n12);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n4);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U12 : INV_X1 port map( A => A(3), ZN => n11);
   U13 : INV_X1 port map( A => B(3), ZN => n10);
   U14 : INV_X1 port map( A => A(2), ZN => n15);
   U15 : INV_X1 port map( A => B(2), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n15, B2 => n8, A => n7, ZN => n19);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n9);
   U19 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => Co);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U23 : INV_X1 port map( A => n16, ZN => n17);
   U24 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_46;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_45;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U8 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U9 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_44;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_43;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_42;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_41;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_40;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_39;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_38;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_37;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_36;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n16, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n15, B => n14, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U11 : XNOR2_X1 port map( A => n13, B => n12, ZN => S(1));
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U16 : INV_X1 port map( A => A(3), ZN => n10);
   U17 : INV_X1 port map( A => B(3), ZN => n9);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U19 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U21 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_35;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U8 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_34;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n12, Z => S(1));
   U2 : XOR2_X1 port map( A => A(1), B => B(1), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n16);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n7);
   U6 : XNOR2_X1 port map( A => n17, B => n16, ZN => S(3));
   U7 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n17);
   U8 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n13);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U11 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U12 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U14 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U15 : INV_X1 port map( A => A(3), ZN => n10);
   U16 : INV_X1 port map( A => B(3), ZN => n9);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n8);
   U18 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U20 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U21 : INV_X1 port map( A => n13, ZN => n14);
   U22 : XOR2_X1 port map( A => n15, B => n14, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_33;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U8 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U9 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_32;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_32 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_31;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n17, B => n16, ZN => S(2));
   U2 : XOR2_X1 port map( A => n1, B => n14, Z => S(1));
   U3 : XNOR2_X1 port map( A => n13, B => B(1), ZN => n1);
   U4 : XOR2_X1 port map( A => n2, B => n18, Z => S(3));
   U5 : XOR2_X1 port map( A => B(3), B => A(3), Z => n2);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n18);
   U7 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n7);
   U8 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n8);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n4);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U12 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n16);
   U13 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n5);
   U14 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n14, ZN => n6);
   U15 : INV_X1 port map( A => A(3), ZN => n11);
   U16 : INV_X1 port map( A => B(3), ZN => n10);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n9);
   U18 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n12);
   U20 : XOR2_X1 port map( A => Ci, B => n12, Z => S(0));
   U21 : INV_X1 port map( A => A(1), ZN => n13);
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_30;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n12, B => n11, ZN => S(1));
   U2 : XNOR2_X1 port map( A => n17, B => n16, ZN => S(3));
   U3 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n17);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n13);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n6);
   U10 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U11 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U14 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n15);
   U15 : INV_X1 port map( A => A(3), ZN => n9);
   U16 : INV_X1 port map( A => B(3), ZN => n8);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n16, ZN => n7);
   U18 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U20 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U21 : INV_X1 port map( A => n13, ZN => n14);
   U22 : XOR2_X1 port map( A => n15, B => n14, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_29;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n19, B => n18, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n15);
   U3 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U4 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n18);
   U6 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U7 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n15, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U9 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U10 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n19);
   U13 : INV_X1 port map( A => A(3), ZN => n9);
   U14 : INV_X1 port map( A => B(3), ZN => n8);
   U15 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n7);
   U16 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U17 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U18 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U19 : INV_X1 port map( A => n11, ZN => n12);
   U20 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U21 : INV_X1 port map( A => A(2), ZN => n14);
   U22 : XOR2_X1 port map( A => n14, B => B(2), Z => n17);
   U23 : INV_X1 port map( A => n15, ZN => n16);
   U24 : XOR2_X1 port map( A => n17, B => n16, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_28;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_27;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_26;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_25;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_24;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_23;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_22;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_21;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_20;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U6 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U8 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U9 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U10 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U11 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U12 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U13 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_19;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U10 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U11 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_18;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1022, 
      n_1023, n_1024 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n9);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n10);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n9, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n10, ZN => n6);
   U10 : INV_X1 port map( A => A(3), ZN => n11);
   U11 : INV_X1 port map( A => B(3), ZN => n8);
   U12 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n12, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n11, B2 => n8, A => n7, ZN => Co);
   U14 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1022, S => 
                           S(0));
   U15 : FA_X1 port map( A => A(1), B => B(1), CI => n9, CO => n_1023, S => 
                           S(1));
   U16 : FA_X1 port map( A => A(2), B => B(2), CI => n10, CO => n_1024, S => 
                           S(2));
   U17 : XOR2_X1 port map( A => n11, B => B(3), Z => n14);
   U18 : INV_X1 port map( A => n12, ZN => n13);
   U19 : XOR2_X1 port map( A => n14, B => n13, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_17;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1025, 
      n_1026, n_1027 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n9);
   U2 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n10);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U6 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n9, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n10, ZN => n6);
   U10 : INV_X1 port map( A => A(3), ZN => n11);
   U11 : INV_X1 port map( A => B(3), ZN => n8);
   U12 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n12, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n11, B2 => n8, A => n7, ZN => Co);
   U14 : FA_X1 port map( A => B(0), B => A(0), CI => Ci, CO => n_1025, S => 
                           S(0));
   U15 : FA_X1 port map( A => A(1), B => B(1), CI => n9, CO => n_1026, S => 
                           S(1));
   U16 : FA_X1 port map( A => A(2), B => B(2), CI => n10, CO => n_1027, S => 
                           S(2));
   U17 : XOR2_X1 port map( A => n11, B => B(3), Z => n14);
   U18 : INV_X1 port map( A => n12, ZN => n13);
   U19 : XOR2_X1 port map( A => n14, B => n13, Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_16;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_16 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_15;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n17);
   U2 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n6);
   U3 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n15, ZN => n7);
   U4 : XOR2_X1 port map( A => n1, B => n15, Z => S(1));
   U5 : XNOR2_X1 port map( A => n14, B => B(1), ZN => n1);
   U6 : XOR2_X1 port map( A => n2, B => n17, Z => S(2));
   U7 : XNOR2_X1 port map( A => n16, B => B(2), ZN => n2);
   U8 : XOR2_X1 port map( A => n3, B => n18, Z => S(3));
   U9 : XOR2_X1 port map( A => B(3), B => A(3), Z => n3);
   U10 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n15);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n4);
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n5);
   U13 : INV_X1 port map( A => A(3), ZN => n12);
   U14 : INV_X1 port map( A => B(3), ZN => n11);
   U15 : INV_X1 port map( A => A(2), ZN => n16);
   U16 : INV_X1 port map( A => B(2), ZN => n9);
   U17 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n17, ZN => n8);
   U18 : OAI21_X1 port map( B1 => n16, B2 => n9, A => n8, ZN => n18);
   U19 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n18, ZN => n10);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n11, A => n10, ZN => Co);
   U21 : XOR2_X1 port map( A => B(0), B => A(0), Z => n13);
   U22 : XOR2_X1 port map( A => Ci, B => n13, Z => S(0));
   U23 : INV_X1 port map( A => A(1), ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_14;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n14, B => n13, ZN => S(2));
   U2 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U3 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n14);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n15);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n13);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n12, B => n11, ZN => S(1));
   U11 : XNOR2_X1 port map( A => n16, B => n15, ZN => S(3));
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n16);
   U13 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U16 : INV_X1 port map( A => A(3), ZN => n9);
   U17 : INV_X1 port map( A => B(3), ZN => n8);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n15, ZN => n7);
   U19 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U21 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_13;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U2 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U3 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_12;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n14, B => n13, ZN => S(2));
   U2 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U3 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n14);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n15);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n13);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n12, B => n11, ZN => S(1));
   U11 : XNOR2_X1 port map( A => n16, B => n15, ZN => S(3));
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n16);
   U13 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U16 : INV_X1 port map( A => A(3), ZN => n9);
   U17 : INV_X1 port map( A => B(3), ZN => n8);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n15, ZN => n7);
   U19 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U21 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_11;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U2 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U3 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_10;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U2 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U9 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U10 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_9;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U2 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U3 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_8;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n14, B => n13, ZN => S(2));
   U2 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n12);
   U3 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n14);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n15);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n13, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n13);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n12, B => n11, ZN => S(1));
   U11 : XNOR2_X1 port map( A => n16, B => n15, ZN => S(3));
   U12 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n16);
   U13 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U15 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U16 : INV_X1 port map( A => A(3), ZN => n9);
   U17 : INV_X1 port map( A => B(3), ZN => n8);
   U18 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n15, ZN => n7);
   U19 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U20 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U21 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_7;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U2 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U3 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U5 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U6 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U8 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U9 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U10 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_6;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U2 : NAND2_X1 port map( A1 => n18, A2 => n17, ZN => n19);
   U3 : XOR2_X1 port map( A => n1, B => n21, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n1);
   U5 : OAI22_X1 port map( A1 => n2, A2 => n7, B1 => n6, B2 => n5, ZN => n22);
   U6 : INV_X1 port map( A => B(2), ZN => n6);
   U7 : INV_X1 port map( A => A(2), ZN => n5);
   U8 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n18, ZN => n7);
   U9 : AND3_X1 port map( A1 => n13, A2 => n14, A3 => n20, ZN => n2);
   U10 : XOR2_X1 port map( A => n3, B => n22, Z => S(3));
   U11 : XOR2_X1 port map( A => B(3), B => A(3), Z => n3);
   U12 : INV_X1 port map( A => A(3), ZN => n10);
   U13 : INV_X1 port map( A => B(3), ZN => n9);
   U14 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n13);
   U15 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n14);
   U16 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n20);
   U17 : INV_X1 port map( A => A(1), ZN => n12);
   U18 : INV_X1 port map( A => B(1), ZN => n4);
   U19 : NAND2_X1 port map( A1 => n12, A2 => n4, ZN => n18);
   U20 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n22, ZN => n8);
   U21 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U22 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U23 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U24 : XOR2_X1 port map( A => n12, B => B(1), Z => n16);
   U25 : NAND2_X1 port map( A1 => n14, A2 => n13, ZN => n17);
   U26 : INV_X1 port map( A => n17, ZN => n15);
   U27 : XOR2_X1 port map( A => n16, B => n15, Z => S(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_5;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n19, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n16);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n13, ZN => n5);
   U9 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n18);
   U10 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n13);
   U11 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U13 : INV_X1 port map( A => A(3), ZN => n10);
   U14 : INV_X1 port map( A => B(3), ZN => n9);
   U15 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n8);
   U16 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U17 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U18 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U19 : INV_X1 port map( A => A(1), ZN => n12);
   U20 : XOR2_X1 port map( A => n12, B => B(1), Z => n15);
   U21 : INV_X1 port map( A => n13, ZN => n14);
   U22 : XOR2_X1 port map( A => n15, B => n14, Z => S(1));
   U23 : INV_X1 port map( A => n16, ZN => n17);
   U24 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_4;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n10, A2 => n11, A3 => n16, ZN => n1);
   U2 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(2));
   U3 : NAND2_X1 port map( A1 => n16, A2 => n15, ZN => n17);
   U4 : NAND2_X1 port map( A1 => n14, A2 => n13, ZN => n15);
   U5 : OAI22_X1 port map( A1 => n1, A2 => n5, B1 => n4, B2 => n3, ZN => n20);
   U6 : INV_X1 port map( A => B(2), ZN => n4);
   U7 : INV_X1 port map( A => A(2), ZN => n3);
   U8 : XNOR2_X1 port map( A => n21, B => n20, ZN => S(3));
   U9 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n5);
   U10 : XNOR2_X1 port map( A => n12, B => n13, ZN => S(1));
   U11 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n18);
   U12 : INV_X1 port map( A => A(3), ZN => n19);
   U13 : INV_X1 port map( A => B(3), ZN => n7);
   U14 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n10);
   U15 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n11);
   U16 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n16);
   U17 : INV_X1 port map( A => A(1), ZN => n9);
   U18 : INV_X1 port map( A => B(1), ZN => n2);
   U19 : NAND2_X1 port map( A1 => n9, A2 => n2, ZN => n14);
   U20 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n20, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n19, B2 => n7, A => n6, ZN => Co);
   U22 : XOR2_X1 port map( A => B(0), B => A(0), Z => n8);
   U23 : XOR2_X1 port map( A => Ci, B => n8, Z => S(0));
   U24 : XOR2_X1 port map( A => n9, B => B(1), Z => n12);
   U25 : NAND2_X1 port map( A1 => n11, A2 => n10, ZN => n13);
   U26 : XOR2_X1 port map( A => n19, B => B(3), Z => n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_3;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => n17, Z => S(3));
   U2 : XOR2_X1 port map( A => B(3), B => A(3), Z => n1);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n17);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n6);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n15, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n15);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n4);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n5);
   U9 : XNOR2_X1 port map( A => n16, B => n15, ZN => S(2));
   U10 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U11 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n14);
   U12 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n12);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n3);
   U14 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n2);
   U15 : INV_X1 port map( A => A(3), ZN => n10);
   U16 : INV_X1 port map( A => B(3), ZN => n9);
   U17 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n8);
   U18 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U19 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U20 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U21 : INV_X1 port map( A => n12, ZN => n13);
   U22 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_2;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n18, B => n17, ZN => S(3));
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n17);
   U3 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n14, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n14);
   U6 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U7 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n11, ZN => n4);
   U8 : XNOR2_X1 port map( A => A(1), B => B(1), ZN => n13);
   U9 : XNOR2_X1 port map( A => A(2), B => B(2), ZN => n16);
   U10 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n18);
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n11);
   U12 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U13 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U14 : INV_X1 port map( A => A(3), ZN => n9);
   U15 : INV_X1 port map( A => B(3), ZN => n8);
   U16 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n17, ZN => n7);
   U17 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U18 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U19 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U20 : INV_X1 port map( A => n11, ZN => n12);
   U21 : XOR2_X1 port map( A => n13, B => n12, Z => S(1));
   U22 : INV_X1 port map( A => n14, ZN => n15);
   U23 : XOR2_X1 port map( A => n16, B => n15, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_1;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(3));
   U2 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n20);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n19);
   U4 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => A(2), A => n16, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n16);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U8 : OAI21_X1 port map( B1 => B(1), B2 => A(1), A => n12, ZN => n4);
   U9 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n12);
   U10 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U11 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U12 : INV_X1 port map( A => A(3), ZN => n9);
   U13 : INV_X1 port map( A => B(3), ZN => n8);
   U14 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n19, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => Co);
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U17 : XOR2_X1 port map( A => Ci, B => n10, Z => S(0));
   U18 : INV_X1 port map( A => A(1), ZN => n11);
   U19 : XOR2_X1 port map( A => n11, B => B(1), Z => n14);
   U20 : INV_X1 port map( A => n12, ZN => n13);
   U21 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U22 : INV_X1 port map( A => A(2), ZN => n15);
   U23 : XOR2_X1 port map( A => n15, B => B(2), Z => n18);
   U24 : INV_X1 port map( A => n16, ZN => n17);
   U25 : XOR2_X1 port map( A => n18, B => n17, Z => S(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_63;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_63 is

   component MUX2to1_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_125
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_126
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1028, n_1029 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_126 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1028);
   RCA0 : RCAN_NBIT4_125 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1029);
   MUX21 : MUX2to1_NBIT4_63 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_62;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_62 is

   component MUX2to1_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_123
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_124
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1030, n_1031 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_124 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1030);
   RCA0 : RCAN_NBIT4_123 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1031);
   MUX21 : MUX2to1_NBIT4_62 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_61;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_61 is

   component MUX2to1_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_121
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_122
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1032, n_1033 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_122 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1032);
   RCA0 : RCAN_NBIT4_121 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1033);
   MUX21 : MUX2to1_NBIT4_61 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_60;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_60 is

   component MUX2to1_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_119
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_120
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1034, n_1035 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_120 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1034);
   RCA0 : RCAN_NBIT4_119 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1035);
   MUX21 : MUX2to1_NBIT4_60 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_59;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_59 is

   component MUX2to1_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_117
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_118
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1036, n_1037 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_118 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1036);
   RCA0 : RCAN_NBIT4_117 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1037);
   MUX21 : MUX2to1_NBIT4_59 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_58;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_58 is

   component MUX2to1_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_115
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_116
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1038, n_1039 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_116 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1038);
   RCA0 : RCAN_NBIT4_115 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1039);
   MUX21 : MUX2to1_NBIT4_58 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_57;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_57 is

   component MUX2to1_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_113
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_114
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1040, n_1041 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_114 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1040);
   RCA0 : RCAN_NBIT4_113 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1041);
   MUX21 : MUX2to1_NBIT4_57 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_56;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_56 is

   component MUX2to1_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_111
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_112
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1042, n_1043 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_112 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1042);
   RCA0 : RCAN_NBIT4_111 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1043);
   MUX21 : MUX2to1_NBIT4_56 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_55;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_55 is

   component MUX2to1_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_109
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_110
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1044, n_1045 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_110 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1044);
   RCA0 : RCAN_NBIT4_109 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1045);
   MUX21 : MUX2to1_NBIT4_55 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_54;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_54 is

   component MUX2to1_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_107
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_108
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1046, n_1047 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_108 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1046);
   RCA0 : RCAN_NBIT4_107 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1047);
   MUX21 : MUX2to1_NBIT4_54 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_53;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_53 is

   component MUX2to1_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_105
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_106
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1048, n_1049 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_106 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1048);
   RCA0 : RCAN_NBIT4_105 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1049);
   MUX21 : MUX2to1_NBIT4_53 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_52;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_52 is

   component MUX2to1_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_103
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_104
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1050, n_1051 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_104 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1050);
   RCA0 : RCAN_NBIT4_103 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1051);
   MUX21 : MUX2to1_NBIT4_52 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_51;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_51 is

   component MUX2to1_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_101
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_102
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1052, n_1053 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_102 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1052);
   RCA0 : RCAN_NBIT4_101 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1053);
   MUX21 : MUX2to1_NBIT4_51 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_50;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_50 is

   component MUX2to1_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_99
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_100
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1054, n_1055 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_100 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1054);
   RCA0 : RCAN_NBIT4_99 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1055);
   MUX21 : MUX2to1_NBIT4_50 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_49;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_49 is

   component MUX2to1_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_97
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_98
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1056, n_1057 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_98 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1056);
   RCA0 : RCAN_NBIT4_97 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1057);
   MUX21 : MUX2to1_NBIT4_49 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_48;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_48 is

   component MUX2to1_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_95
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_96
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1058, n_1059 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_96 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1058);
   RCA0 : RCAN_NBIT4_95 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1059);
   MUX21 : MUX2to1_NBIT4_48 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_47;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_47 is

   component MUX2to1_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_93
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_94
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1060, n_1061 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_94 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1060);
   RCA0 : RCAN_NBIT4_93 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1061);
   MUX21 : MUX2to1_NBIT4_47 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_46;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_46 is

   component MUX2to1_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_91
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_92
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1062, n_1063 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_92 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1062);
   RCA0 : RCAN_NBIT4_91 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1063);
   MUX21 : MUX2to1_NBIT4_46 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_45;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_45 is

   component MUX2to1_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_89
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_90
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1064, n_1065 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_90 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1064);
   RCA0 : RCAN_NBIT4_89 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1065);
   MUX21 : MUX2to1_NBIT4_45 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_44;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_44 is

   component MUX2to1_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_87
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_88
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1066, n_1067 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_88 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1066);
   RCA0 : RCAN_NBIT4_87 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1067);
   MUX21 : MUX2to1_NBIT4_44 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_43;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_43 is

   component MUX2to1_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_85
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_86
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1068, n_1069 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_86 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1068);
   RCA0 : RCAN_NBIT4_85 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1069);
   MUX21 : MUX2to1_NBIT4_43 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_42;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_42 is

   component MUX2to1_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_83
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_84
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1070, n_1071 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_84 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1070);
   RCA0 : RCAN_NBIT4_83 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1071);
   MUX21 : MUX2to1_NBIT4_42 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_41;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_41 is

   component MUX2to1_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_81
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_82
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1072, n_1073 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_82 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1072);
   RCA0 : RCAN_NBIT4_81 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1073);
   MUX21 : MUX2to1_NBIT4_41 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_40;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_40 is

   component MUX2to1_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_79
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_80
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1074, n_1075 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_80 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1074);
   RCA0 : RCAN_NBIT4_79 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1075);
   MUX21 : MUX2to1_NBIT4_40 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_39;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_39 is

   component MUX2to1_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_77
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_78
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1076, n_1077 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_78 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1076);
   RCA0 : RCAN_NBIT4_77 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1077);
   MUX21 : MUX2to1_NBIT4_39 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_38;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_38 is

   component MUX2to1_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_75
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_76
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1078, n_1079 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_76 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1078);
   RCA0 : RCAN_NBIT4_75 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1079);
   MUX21 : MUX2to1_NBIT4_38 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_37;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_37 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2to1_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_73
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_74
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n1, n_1080, n_1081
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_74 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1080);
   RCA0 : RCAN_NBIT4_73 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => n1, B(3) => B(3), B(2) => B(2), B(1) => B(1)
                           , B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1081);
   MUX21 : MUX2to1_NBIT4_37 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : BUF_X1 port map( A => A(0), Z => n1);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_36;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_36 is

   component MUX2to1_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_71
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_72
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1082, n_1083 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_72 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1082);
   RCA0 : RCAN_NBIT4_71 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1083);
   MUX21 : MUX2to1_NBIT4_36 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_35;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_35 is

   component MUX2to1_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_69
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_70
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1084, n_1085 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_70 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1084);
   RCA0 : RCAN_NBIT4_69 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1085);
   MUX21 : MUX2to1_NBIT4_35 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_34;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_34 is

   component MUX2to1_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_67
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_68
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1086, n_1087 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_68 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1086);
   RCA0 : RCAN_NBIT4_67 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1087);
   MUX21 : MUX2to1_NBIT4_34 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_33;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_33 is

   component MUX2to1_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_65
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_66
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1088, n_1089 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_66 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1088);
   RCA0 : RCAN_NBIT4_65 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1089);
   MUX21 : MUX2to1_NBIT4_33 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_32;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_32 is

   component MUX2to1_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_64
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1090, n_1091 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_64 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1090);
   RCA0 : RCAN_NBIT4_63 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1091);
   MUX21 : MUX2to1_NBIT4_32 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_31;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_31 is

   component MUX2to1_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1092, n_1093 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_62 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1092);
   RCA0 : RCAN_NBIT4_61 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1093);
   MUX21 : MUX2to1_NBIT4_31 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_30;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_30 is

   component MUX2to1_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1094, n_1095 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_60 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1094);
   RCA0 : RCAN_NBIT4_59 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1095);
   MUX21 : MUX2to1_NBIT4_30 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_29;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_29 is

   component MUX2to1_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1096, n_1097 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_58 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1096);
   RCA0 : RCAN_NBIT4_57 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1097);
   MUX21 : MUX2to1_NBIT4_29 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_28;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_28 is

   component MUX2to1_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1098, n_1099 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1098);
   RCA0 : RCAN_NBIT4_55 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1099);
   MUX21 : MUX2to1_NBIT4_28 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_27;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_27 is

   component MUX2to1_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1100, n_1101 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_54 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1100);
   RCA0 : RCAN_NBIT4_53 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1101);
   MUX21 : MUX2to1_NBIT4_27 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_26;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_26 is

   component MUX2to1_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1102, n_1103 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_52 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1102);
   RCA0 : RCAN_NBIT4_51 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1103);
   MUX21 : MUX2to1_NBIT4_26 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_25;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_25 is

   component MUX2to1_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1104, n_1105 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_50 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1104);
   RCA0 : RCAN_NBIT4_49 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1105);
   MUX21 : MUX2to1_NBIT4_25 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_24;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_24 is

   component MUX2to1_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1106, n_1107 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1106);
   RCA0 : RCAN_NBIT4_47 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1107);
   MUX21 : MUX2to1_NBIT4_24 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_23;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_23 is

   component MUX2to1_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1108, n_1109 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_46 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1108);
   RCA0 : RCAN_NBIT4_45 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1109);
   MUX21 : MUX2to1_NBIT4_23 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_22;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_22 is

   component MUX2to1_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1110, n_1111 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_44 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1110);
   RCA0 : RCAN_NBIT4_43 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1111);
   MUX21 : MUX2to1_NBIT4_22 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_21;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_21 is

   component MUX2to1_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1112, n_1113 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_42 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1112);
   RCA0 : RCAN_NBIT4_41 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1113);
   MUX21 : MUX2to1_NBIT4_21 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_20;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_20 is

   component MUX2to1_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1114, n_1115 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1114);
   RCA0 : RCAN_NBIT4_39 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1115);
   MUX21 : MUX2to1_NBIT4_20 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_19;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_19 is

   component MUX2to1_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1116, n_1117 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_38 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1116);
   RCA0 : RCAN_NBIT4_37 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1117);
   MUX21 : MUX2to1_NBIT4_19 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_18;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_18 is

   component MUX2to1_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1118, n_1119 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_36 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1118);
   RCA0 : RCAN_NBIT4_35 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1119);
   MUX21 : MUX2to1_NBIT4_18 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_17;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_17 is

   component MUX2to1_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1120, n_1121 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_34 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1120);
   RCA0 : RCAN_NBIT4_33 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1121);
   MUX21 : MUX2to1_NBIT4_17 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_16;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_16 is

   component MUX2to1_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1122, n_1123 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1122);
   RCA0 : RCAN_NBIT4_31 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1123);
   MUX21 : MUX2to1_NBIT4_16 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_15;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_15 is

   component MUX2to1_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1124, n_1125 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1124);
   RCA0 : RCAN_NBIT4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1125);
   MUX21 : MUX2to1_NBIT4_15 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_14;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_14 is

   component MUX2to1_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1126, n_1127 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1126);
   RCA0 : RCAN_NBIT4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1127);
   MUX21 : MUX2to1_NBIT4_14 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_13;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_13 is

   component MUX2to1_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1128, n_1129 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1128);
   RCA0 : RCAN_NBIT4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1129);
   MUX21 : MUX2to1_NBIT4_13 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_12;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_12 is

   component MUX2to1_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1130, n_1131 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1130);
   RCA0 : RCAN_NBIT4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1131);
   MUX21 : MUX2to1_NBIT4_12 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_11;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_11 is

   component MUX2to1_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1132, n_1133 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1132);
   RCA0 : RCAN_NBIT4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1133);
   MUX21 : MUX2to1_NBIT4_11 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_10;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_10 is

   component MUX2to1_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1134, n_1135 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1134);
   RCA0 : RCAN_NBIT4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1135);
   MUX21 : MUX2to1_NBIT4_10 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_9;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_9 is

   component MUX2to1_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1136, n_1137 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1136);
   RCA0 : RCAN_NBIT4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1137);
   MUX21 : MUX2to1_NBIT4_9 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_8;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_8 is

   component MUX2to1_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1138, n_1139 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1138);
   RCA0 : RCAN_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1139);
   MUX21 : MUX2to1_NBIT4_8 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_7;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_7 is

   component MUX2to1_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1140, n_1141 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1140);
   RCA0 : RCAN_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1141);
   MUX21 : MUX2to1_NBIT4_7 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_6;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_6 is

   component MUX2to1_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1142, n_1143 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1142);
   RCA0 : RCAN_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1143);
   MUX21 : MUX2to1_NBIT4_6 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_5;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_5 is

   component MUX2to1_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1144, n_1145 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1144);
   RCA0 : RCAN_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1145);
   MUX21 : MUX2to1_NBIT4_5 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_4;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_4 is

   component MUX2to1_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1146, n_1147 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1146);
   RCA0 : RCAN_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1147);
   MUX21 : MUX2to1_NBIT4_4 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_3;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_3 is

   component MUX2to1_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1148, n_1149 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1148);
   RCA0 : RCAN_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1149);
   MUX21 : MUX2to1_NBIT4_3 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_2;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_2 is

   component MUX2to1_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1150, n_1151 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1150);
   RCA0 : RCAN_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1151);
   MUX21 : MUX2to1_NBIT4_2 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_1;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_1 is

   component MUX2to1_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1152, n_1153 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1152);
   RCA0 : RCAN_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1153);
   MUX21 : MUX2to1_NBIT4_1 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_215 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_215;

architecture SYN_BEHAVIORAL of PG_block_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_214 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_214;

architecture SYN_BEHAVIORAL of PG_block_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_213 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_213;

architecture SYN_BEHAVIORAL of PG_block_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_212 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_212;

architecture SYN_BEHAVIORAL of PG_block_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_211 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_211;

architecture SYN_BEHAVIORAL of PG_block_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_210 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_210;

architecture SYN_BEHAVIORAL of PG_block_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_209 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_209;

architecture SYN_BEHAVIORAL of PG_block_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_208 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_208;

architecture SYN_BEHAVIORAL of PG_block_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_207 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_207;

architecture SYN_BEHAVIORAL of PG_block_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_206 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_206;

architecture SYN_BEHAVIORAL of PG_block_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_205 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_205;

architecture SYN_BEHAVIORAL of PG_block_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_204 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_204;

architecture SYN_BEHAVIORAL of PG_block_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_203 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_203;

architecture SYN_BEHAVIORAL of PG_block_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_202 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_202;

architecture SYN_BEHAVIORAL of PG_block_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_201 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_201;

architecture SYN_BEHAVIORAL of PG_block_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_200 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_200;

architecture SYN_BEHAVIORAL of PG_block_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_199 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_199;

architecture SYN_BEHAVIORAL of PG_block_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_198 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_198;

architecture SYN_BEHAVIORAL of PG_block_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_197 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_197;

architecture SYN_BEHAVIORAL of PG_block_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_196 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_196;

architecture SYN_BEHAVIORAL of PG_block_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n2, A2 => A(0), ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(1), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_195 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_195;

architecture SYN_BEHAVIORAL of PG_block_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_194 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_194;

architecture SYN_BEHAVIORAL of PG_block_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_193 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_193;

architecture SYN_BEHAVIORAL of PG_block_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_192 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_192;

architecture SYN_BEHAVIORAL of PG_block_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_191 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_191;

architecture SYN_BEHAVIORAL of PG_block_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n2, A2 => A(0), ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(1), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_190 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_190;

architecture SYN_BEHAVIORAL of PG_block_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_189 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_189;

architecture SYN_BEHAVIORAL of PG_block_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_188 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_188;

architecture SYN_BEHAVIORAL of PG_block_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_187 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_187;

architecture SYN_BEHAVIORAL of PG_block_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_186 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_186;

architecture SYN_BEHAVIORAL of PG_block_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_185 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_185;

architecture SYN_BEHAVIORAL of PG_block_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_184 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_184;

architecture SYN_BEHAVIORAL of PG_block_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_183 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_183;

architecture SYN_BEHAVIORAL of PG_block_183 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_182 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_182;

architecture SYN_BEHAVIORAL of PG_block_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_181 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_181;

architecture SYN_BEHAVIORAL of PG_block_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_180 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_180;

architecture SYN_BEHAVIORAL of PG_block_180 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_179 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_179;

architecture SYN_BEHAVIORAL of PG_block_179 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_178 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_178;

architecture SYN_BEHAVIORAL of PG_block_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_177 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_177;

architecture SYN_BEHAVIORAL of PG_block_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_176 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_176;

architecture SYN_BEHAVIORAL of PG_block_176 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_175 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_175;

architecture SYN_BEHAVIORAL of PG_block_175 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_174 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_174;

architecture SYN_BEHAVIORAL of PG_block_174 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_173 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_173;

architecture SYN_BEHAVIORAL of PG_block_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_172 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_172;

architecture SYN_BEHAVIORAL of PG_block_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_171 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_171;

architecture SYN_BEHAVIORAL of PG_block_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_170 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_170;

architecture SYN_BEHAVIORAL of PG_block_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_169 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_169;

architecture SYN_BEHAVIORAL of PG_block_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_168 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_168;

architecture SYN_BEHAVIORAL of PG_block_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_167 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_167;

architecture SYN_BEHAVIORAL of PG_block_167 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_166 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_166;

architecture SYN_BEHAVIORAL of PG_block_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_165 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_165;

architecture SYN_BEHAVIORAL of PG_block_165 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_164 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_164;

architecture SYN_BEHAVIORAL of PG_block_164 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_163 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_163;

architecture SYN_BEHAVIORAL of PG_block_163 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_162 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_162;

architecture SYN_BEHAVIORAL of PG_block_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_161 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_161;

architecture SYN_BEHAVIORAL of PG_block_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_160 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_160;

architecture SYN_BEHAVIORAL of PG_block_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_159 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_159;

architecture SYN_BEHAVIORAL of PG_block_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_158 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_158;

architecture SYN_BEHAVIORAL of PG_block_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_157 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_157;

architecture SYN_BEHAVIORAL of PG_block_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_156 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_156;

architecture SYN_BEHAVIORAL of PG_block_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_155 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_155;

architecture SYN_BEHAVIORAL of PG_block_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_154 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_154;

architecture SYN_BEHAVIORAL of PG_block_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_153 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_153;

architecture SYN_BEHAVIORAL of PG_block_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_152 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_152;

architecture SYN_BEHAVIORAL of PG_block_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_151 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_151;

architecture SYN_BEHAVIORAL of PG_block_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_150 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_150;

architecture SYN_BEHAVIORAL of PG_block_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_149 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_149;

architecture SYN_BEHAVIORAL of PG_block_149 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_148 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_148;

architecture SYN_BEHAVIORAL of PG_block_148 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_147 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_147;

architecture SYN_BEHAVIORAL of PG_block_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_146 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_146;

architecture SYN_BEHAVIORAL of PG_block_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_145 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_145;

architecture SYN_BEHAVIORAL of PG_block_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_144 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_144;

architecture SYN_BEHAVIORAL of PG_block_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_143 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_143;

architecture SYN_BEHAVIORAL of PG_block_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_142 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_142;

architecture SYN_BEHAVIORAL of PG_block_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_141 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_141;

architecture SYN_BEHAVIORAL of PG_block_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_140 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_140;

architecture SYN_BEHAVIORAL of PG_block_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_139 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_139;

architecture SYN_BEHAVIORAL of PG_block_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_138 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_138;

architecture SYN_BEHAVIORAL of PG_block_138 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_137 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_137;

architecture SYN_BEHAVIORAL of PG_block_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_136 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_136;

architecture SYN_BEHAVIORAL of PG_block_136 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_135 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_135;

architecture SYN_BEHAVIORAL of PG_block_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_134 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_134;

architecture SYN_BEHAVIORAL of PG_block_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_133 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_133;

architecture SYN_BEHAVIORAL of PG_block_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_132 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_132;

architecture SYN_BEHAVIORAL of PG_block_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_131 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_131;

architecture SYN_BEHAVIORAL of PG_block_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_130 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_130;

architecture SYN_BEHAVIORAL of PG_block_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PGout(0));
   U2 : INV_X1 port map( A => A(1), ZN => n1);
   U3 : INV_X1 port map( A => B(0), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_129 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_129;

architecture SYN_BEHAVIORAL of PG_block_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_128 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_128;

architecture SYN_BEHAVIORAL of PG_block_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_127 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_127;

architecture SYN_BEHAVIORAL of PG_block_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_126 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_126;

architecture SYN_BEHAVIORAL of PG_block_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_125 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_125;

architecture SYN_BEHAVIORAL of PG_block_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_124 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_124;

architecture SYN_BEHAVIORAL of PG_block_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_123 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_123;

architecture SYN_BEHAVIORAL of PG_block_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_122 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_122;

architecture SYN_BEHAVIORAL of PG_block_122 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_121 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_121;

architecture SYN_BEHAVIORAL of PG_block_121 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_120 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_120;

architecture SYN_BEHAVIORAL of PG_block_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_119 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_119;

architecture SYN_BEHAVIORAL of PG_block_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_118 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_118;

architecture SYN_BEHAVIORAL of PG_block_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_117 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_117;

architecture SYN_BEHAVIORAL of PG_block_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_116 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_116;

architecture SYN_BEHAVIORAL of PG_block_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_115 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_115;

architecture SYN_BEHAVIORAL of PG_block_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PGout(0));
   U2 : INV_X1 port map( A => B(0), ZN => n1);
   U3 : INV_X1 port map( A => A(1), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_114 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_114;

architecture SYN_BEHAVIORAL of PG_block_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_113 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_113;

architecture SYN_BEHAVIORAL of PG_block_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : INV_X2 port map( A => A(1), ZN => n2);
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PGout(0));
   U3 : INV_X1 port map( A => B(0), ZN => n1);
   U4 : INV_X1 port map( A => A(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_112 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_112;

architecture SYN_BEHAVIORAL of PG_block_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PGout(0));
   U2 : INV_X1 port map( A => B(0), ZN => n1);
   U3 : INV_X1 port map( A => A(1), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_111 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_111;

architecture SYN_BEHAVIORAL of PG_block_111 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_110 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_110;

architecture SYN_BEHAVIORAL of PG_block_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_109 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_109;

architecture SYN_BEHAVIORAL of PG_block_109 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_108 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_108;

architecture SYN_BEHAVIORAL of PG_block_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_107 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_107;

architecture SYN_BEHAVIORAL of PG_block_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_106 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_106;

architecture SYN_BEHAVIORAL of PG_block_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_105 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_105;

architecture SYN_BEHAVIORAL of PG_block_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_104 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_104;

architecture SYN_BEHAVIORAL of PG_block_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_103 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_103;

architecture SYN_BEHAVIORAL of PG_block_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_102 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_102;

architecture SYN_BEHAVIORAL of PG_block_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_101 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_101;

architecture SYN_BEHAVIORAL of PG_block_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_100 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_100;

architecture SYN_BEHAVIORAL of PG_block_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_99 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_99;

architecture SYN_BEHAVIORAL of PG_block_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_98 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_98;

architecture SYN_BEHAVIORAL of PG_block_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_97 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_97;

architecture SYN_BEHAVIORAL of PG_block_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_96 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_96;

architecture SYN_BEHAVIORAL of PG_block_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_95 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_95;

architecture SYN_BEHAVIORAL of PG_block_95 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_94 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_94;

architecture SYN_BEHAVIORAL of PG_block_94 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_93 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_93;

architecture SYN_BEHAVIORAL of PG_block_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_92 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_92;

architecture SYN_BEHAVIORAL of PG_block_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_91 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_91;

architecture SYN_BEHAVIORAL of PG_block_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_90 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_90;

architecture SYN_BEHAVIORAL of PG_block_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_89 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_89;

architecture SYN_BEHAVIORAL of PG_block_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_88 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_88;

architecture SYN_BEHAVIORAL of PG_block_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_87 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_87;

architecture SYN_BEHAVIORAL of PG_block_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_86 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_86;

architecture SYN_BEHAVIORAL of PG_block_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_85 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_85;

architecture SYN_BEHAVIORAL of PG_block_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_84 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_84;

architecture SYN_BEHAVIORAL of PG_block_84 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_83 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_83;

architecture SYN_BEHAVIORAL of PG_block_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_82 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_82;

architecture SYN_BEHAVIORAL of PG_block_82 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_81 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_81;

architecture SYN_BEHAVIORAL of PG_block_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_80 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_80;

architecture SYN_BEHAVIORAL of PG_block_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_79 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_79;

architecture SYN_BEHAVIORAL of PG_block_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_78 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_78;

architecture SYN_BEHAVIORAL of PG_block_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_77 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_77;

architecture SYN_BEHAVIORAL of PG_block_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_76 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_76;

architecture SYN_BEHAVIORAL of PG_block_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_75 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_75;

architecture SYN_BEHAVIORAL of PG_block_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_74 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_74;

architecture SYN_BEHAVIORAL of PG_block_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_73 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_73;

architecture SYN_BEHAVIORAL of PG_block_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_72 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_72;

architecture SYN_BEHAVIORAL of PG_block_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_71 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_71;

architecture SYN_BEHAVIORAL of PG_block_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_70 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_70;

architecture SYN_BEHAVIORAL of PG_block_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_69 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_69;

architecture SYN_BEHAVIORAL of PG_block_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => A(1), A2 => B(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_68 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_68;

architecture SYN_BEHAVIORAL of PG_block_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_67 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_67;

architecture SYN_BEHAVIORAL of PG_block_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_66 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_66;

architecture SYN_BEHAVIORAL of PG_block_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_65 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_65;

architecture SYN_BEHAVIORAL of PG_block_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_64 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_64;

architecture SYN_BEHAVIORAL of PG_block_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_63 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_63;

architecture SYN_BEHAVIORAL of PG_block_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_62 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_62;

architecture SYN_BEHAVIORAL of PG_block_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_61 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_61;

architecture SYN_BEHAVIORAL of PG_block_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_60 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_60;

architecture SYN_BEHAVIORAL of PG_block_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_59 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_59;

architecture SYN_BEHAVIORAL of PG_block_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PGout(0));
   U2 : INV_X1 port map( A => B(0), ZN => n1);
   U3 : INV_X1 port map( A => A(1), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_58 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_58;

architecture SYN_BEHAVIORAL of PG_block_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PGout(0));
   U2 : INV_X1 port map( A => B(0), ZN => n1);
   U3 : INV_X1 port map( A => A(1), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_57 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_57;

architecture SYN_BEHAVIORAL of PG_block_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_56 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_56;

architecture SYN_BEHAVIORAL of PG_block_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_55 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_55;

architecture SYN_BEHAVIORAL of PG_block_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_54 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_54;

architecture SYN_BEHAVIORAL of PG_block_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_53 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_53;

architecture SYN_BEHAVIORAL of PG_block_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_52 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_52;

architecture SYN_BEHAVIORAL of PG_block_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_51 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_51;

architecture SYN_BEHAVIORAL of PG_block_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_50 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_50;

architecture SYN_BEHAVIORAL of PG_block_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_49 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_49;

architecture SYN_BEHAVIORAL of PG_block_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_48 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_48;

architecture SYN_BEHAVIORAL of PG_block_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_47 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_47;

architecture SYN_BEHAVIORAL of PG_block_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_46 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_46;

architecture SYN_BEHAVIORAL of PG_block_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_45 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_45;

architecture SYN_BEHAVIORAL of PG_block_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_44 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_44;

architecture SYN_BEHAVIORAL of PG_block_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_43 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_43;

architecture SYN_BEHAVIORAL of PG_block_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_42 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_42;

architecture SYN_BEHAVIORAL of PG_block_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_41 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_41;

architecture SYN_BEHAVIORAL of PG_block_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_40 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_40;

architecture SYN_BEHAVIORAL of PG_block_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_39 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_39;

architecture SYN_BEHAVIORAL of PG_block_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_38 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_38;

architecture SYN_BEHAVIORAL of PG_block_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_37 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_37;

architecture SYN_BEHAVIORAL of PG_block_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_36 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_36;

architecture SYN_BEHAVIORAL of PG_block_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_35 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_35;

architecture SYN_BEHAVIORAL of PG_block_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_34 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_34;

architecture SYN_BEHAVIORAL of PG_block_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_33 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_33;

architecture SYN_BEHAVIORAL of PG_block_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_32 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_32;

architecture SYN_BEHAVIORAL of PG_block_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_31 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_31;

architecture SYN_BEHAVIORAL of PG_block_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_30 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_30;

architecture SYN_BEHAVIORAL of PG_block_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_29 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_29;

architecture SYN_BEHAVIORAL of PG_block_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_28 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_28;

architecture SYN_BEHAVIORAL of PG_block_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_27 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_27;

architecture SYN_BEHAVIORAL of PG_block_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_26 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_26;

architecture SYN_BEHAVIORAL of PG_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_25 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_25;

architecture SYN_BEHAVIORAL of PG_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_24 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_24;

architecture SYN_BEHAVIORAL of PG_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_23 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_23;

architecture SYN_BEHAVIORAL of PG_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_22 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_22;

architecture SYN_BEHAVIORAL of PG_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_21 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_21;

architecture SYN_BEHAVIORAL of PG_block_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_20 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_20;

architecture SYN_BEHAVIORAL of PG_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_19 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_19;

architecture SYN_BEHAVIORAL of PG_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_18 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_18;

architecture SYN_BEHAVIORAL of PG_block_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_17 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_17;

architecture SYN_BEHAVIORAL of PG_block_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_16 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_16;

architecture SYN_BEHAVIORAL of PG_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_15 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_15;

architecture SYN_BEHAVIORAL of PG_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_14 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_14;

architecture SYN_BEHAVIORAL of PG_block_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_13 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_13;

architecture SYN_BEHAVIORAL of PG_block_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_12 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_12;

architecture SYN_BEHAVIORAL of PG_block_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_11 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_11;

architecture SYN_BEHAVIORAL of PG_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_10 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_10;

architecture SYN_BEHAVIORAL of PG_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_9 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_9;

architecture SYN_BEHAVIORAL of PG_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_8 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_8;

architecture SYN_BEHAVIORAL of PG_block_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_7 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_7;

architecture SYN_BEHAVIORAL of PG_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_6 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_6;

architecture SYN_BEHAVIORAL of PG_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_5 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_5;

architecture SYN_BEHAVIORAL of PG_block_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_4 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_4;

architecture SYN_BEHAVIORAL of PG_block_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_3 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_3;

architecture SYN_BEHAVIORAL of PG_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_2 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_2;

architecture SYN_BEHAVIORAL of PG_block_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => B(0), A2 => A(0), B1 => A(0), B2 => A(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_1 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_1;

architecture SYN_BEHAVIORAL of PG_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_71 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_71;

architecture SYN_BEHAVIORAL of G_block_71 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_70 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_70;

architecture SYN_BEHAVIORAL of G_block_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => A(1), A2 => A(0), B1 => B, B2 => A(0), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_69 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_69;

architecture SYN_BEHAVIORAL of G_block_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_68 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_68;

architecture SYN_BEHAVIORAL of G_block_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_67 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_67;

architecture SYN_BEHAVIORAL of G_block_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_66 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_66;

architecture SYN_BEHAVIORAL of G_block_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_65 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_65;

architecture SYN_BEHAVIORAL of G_block_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_64 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_64;

architecture SYN_BEHAVIORAL of G_block_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_63 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_63;

architecture SYN_BEHAVIORAL of G_block_63 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_62 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_62;

architecture SYN_BEHAVIORAL of G_block_62 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_61 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_61;

architecture SYN_BEHAVIORAL of G_block_61 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_60 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_60;

architecture SYN_BEHAVIORAL of G_block_60 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_59 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_59;

architecture SYN_BEHAVIORAL of G_block_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_58 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_58;

architecture SYN_BEHAVIORAL of G_block_58 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_57 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_57;

architecture SYN_BEHAVIORAL of G_block_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_56 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_56;

architecture SYN_BEHAVIORAL of G_block_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_55 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_55;

architecture SYN_BEHAVIORAL of G_block_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_54 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_54;

architecture SYN_BEHAVIORAL of G_block_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_53 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_53;

architecture SYN_BEHAVIORAL of G_block_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_52 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_52;

architecture SYN_BEHAVIORAL of G_block_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_51 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_51;

architecture SYN_BEHAVIORAL of G_block_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_50 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_50;

architecture SYN_BEHAVIORAL of G_block_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_49 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_49;

architecture SYN_BEHAVIORAL of G_block_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_48 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_48;

architecture SYN_BEHAVIORAL of G_block_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_47 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_47;

architecture SYN_BEHAVIORAL of G_block_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_46 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_46;

architecture SYN_BEHAVIORAL of G_block_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_45 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_45;

architecture SYN_BEHAVIORAL of G_block_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_44 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_44;

architecture SYN_BEHAVIORAL of G_block_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_43 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_43;

architecture SYN_BEHAVIORAL of G_block_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_42 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_42;

architecture SYN_BEHAVIORAL of G_block_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_41 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_41;

architecture SYN_BEHAVIORAL of G_block_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X2 port map( A1 => n2, A2 => A(0), ZN => Gout);
   U2 : AND2_X1 port map( A1 => B, A2 => A(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_40 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_40;

architecture SYN_BEHAVIORAL of G_block_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_39 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_39;

architecture SYN_BEHAVIORAL of G_block_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_38 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_38;

architecture SYN_BEHAVIORAL of G_block_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_37 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_37;

architecture SYN_BEHAVIORAL of G_block_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_36 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_36;

architecture SYN_BEHAVIORAL of G_block_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_35 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_35;

architecture SYN_BEHAVIORAL of G_block_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_34 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_34;

architecture SYN_BEHAVIORAL of G_block_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_33 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_33;

architecture SYN_BEHAVIORAL of G_block_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_32 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_32;

architecture SYN_BEHAVIORAL of G_block_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_31 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_31;

architecture SYN_BEHAVIORAL of G_block_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_30 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_30;

architecture SYN_BEHAVIORAL of G_block_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_29 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_29;

architecture SYN_BEHAVIORAL of G_block_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_28 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_28;

architecture SYN_BEHAVIORAL of G_block_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_27 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_27;

architecture SYN_BEHAVIORAL of G_block_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_26 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_26;

architecture SYN_BEHAVIORAL of G_block_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_25 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_25;

architecture SYN_BEHAVIORAL of G_block_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_24 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_24;

architecture SYN_BEHAVIORAL of G_block_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_23 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_23;

architecture SYN_BEHAVIORAL of G_block_23 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X2 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_22 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_22;

architecture SYN_BEHAVIORAL of G_block_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_21 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_21;

architecture SYN_BEHAVIORAL of G_block_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_20 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_20;

architecture SYN_BEHAVIORAL of G_block_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X2 port map( B1 => n1, B2 => n2, A => n3, ZN => Gout);
   U2 : INV_X1 port map( A => B, ZN => n1);
   U3 : INV_X1 port map( A => A(1), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_19 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_19;

architecture SYN_BEHAVIORAL of G_block_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_18 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_18;

architecture SYN_BEHAVIORAL of G_block_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_17 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_17;

architecture SYN_BEHAVIORAL of G_block_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => B, A2 => A(0), B1 => A(0), B2 => A(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_16 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_16;

architecture SYN_BEHAVIORAL of G_block_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => B, A2 => A(0), B1 => A(0), B2 => A(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_15 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_15;

architecture SYN_BEHAVIORAL of G_block_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_14 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_14;

architecture SYN_BEHAVIORAL of G_block_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => B, A2 => A(0), B1 => A(0), B2 => A(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_13 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_13;

architecture SYN_BEHAVIORAL of G_block_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_12 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_12;

architecture SYN_BEHAVIORAL of G_block_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_11 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_11;

architecture SYN_BEHAVIORAL of G_block_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_10 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_10;

architecture SYN_BEHAVIORAL of G_block_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_9 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_9;

architecture SYN_BEHAVIORAL of G_block_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_8 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_8;

architecture SYN_BEHAVIORAL of G_block_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_7 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_7;

architecture SYN_BEHAVIORAL of G_block_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_6 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_6;

architecture SYN_BEHAVIORAL of G_block_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_5 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_5;

architecture SYN_BEHAVIORAL of G_block_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_4 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_4;

architecture SYN_BEHAVIORAL of G_block_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_3 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_3;

architecture SYN_BEHAVIORAL of G_block_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_2 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_2;

architecture SYN_BEHAVIORAL of G_block_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_1 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_1;

architecture SYN_BEHAVIORAL of G_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_7;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U2 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U3 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U4 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U5 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U6 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U7 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U8 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U9 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U10 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U11 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U14 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U18 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U20 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U21 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U22 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U23 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U24 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U25 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U26 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U27 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U28 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U29 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U30 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_6;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U64 : XOR2_X1 port map( A => n1, B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U2 : AND2_X1 port map( A1 => A(14), A2 => B(14), ZN => Gout(14));
   U3 : CLKBUF_X1 port map( A => B(0), Z => n1);
   U4 : AND2_X1 port map( A1 => A(4), A2 => B(4), ZN => Gout(4));
   U5 : AND2_X1 port map( A1 => A(5), A2 => B(5), ZN => Gout(5));
   U6 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U7 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U8 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U9 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U10 : INV_X1 port map( A => A(1), ZN => n3);
   U11 : INV_X1 port map( A => B(1), ZN => n2);
   U12 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Gout(1));
   U13 : INV_X1 port map( A => A(2), ZN => n5);
   U14 : INV_X1 port map( A => B(2), ZN => n4);
   U15 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Gout(2));
   U16 : INV_X1 port map( A => A(3), ZN => n7);
   U17 : INV_X1 port map( A => B(3), ZN => n6);
   U18 : NOR2_X1 port map( A1 => n7, A2 => n6, ZN => Gout(3));
   U19 : INV_X1 port map( A => A(6), ZN => n9);
   U20 : INV_X1 port map( A => B(6), ZN => n8);
   U21 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => Gout(6));
   U22 : INV_X1 port map( A => A(7), ZN => n11);
   U23 : INV_X1 port map( A => B(7), ZN => n10);
   U24 : NOR2_X1 port map( A1 => n11, A2 => n10, ZN => Gout(7));
   U25 : INV_X1 port map( A => A(8), ZN => n13);
   U26 : INV_X1 port map( A => B(8), ZN => n12);
   U27 : NOR2_X1 port map( A1 => n13, A2 => n12, ZN => Gout(8));
   U28 : INV_X1 port map( A => A(9), ZN => n15);
   U29 : INV_X1 port map( A => B(9), ZN => n14);
   U30 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => Gout(9));
   U31 : INV_X1 port map( A => A(10), ZN => n17);
   U32 : INV_X1 port map( A => B(10), ZN => n16);
   U33 : NOR2_X1 port map( A1 => n17, A2 => n16, ZN => Gout(10));
   U34 : INV_X1 port map( A => A(11), ZN => n19);
   U35 : INV_X1 port map( A => B(11), ZN => n18);
   U36 : NOR2_X1 port map( A1 => n19, A2 => n18, ZN => Gout(11));
   U37 : INV_X1 port map( A => A(12), ZN => n21);
   U38 : INV_X1 port map( A => B(12), ZN => n20);
   U39 : NOR2_X1 port map( A1 => n21, A2 => n20, ZN => Gout(12));
   U42 : INV_X1 port map( A => A(13), ZN => n23);
   U45 : INV_X1 port map( A => B(13), ZN => n22);
   U46 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => Gout(13));
   U47 : INV_X1 port map( A => A(15), ZN => n25);
   U48 : INV_X1 port map( A => B(15), ZN => n24);
   U49 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => Gout(15));
   U50 : INV_X1 port map( A => A(16), ZN => n27);
   U51 : INV_X1 port map( A => B(16), ZN => n26);
   U52 : NOR2_X1 port map( A1 => n27, A2 => n26, ZN => Gout(16));
   U53 : INV_X1 port map( A => A(17), ZN => n29);
   U54 : INV_X1 port map( A => B(17), ZN => n28);
   U55 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => Gout(17));
   U56 : INV_X1 port map( A => A(18), ZN => n31);
   U57 : INV_X1 port map( A => B(18), ZN => n30);
   U58 : NOR2_X1 port map( A1 => n31, A2 => n30, ZN => Gout(18));
   U59 : INV_X1 port map( A => A(19), ZN => n33);
   U60 : INV_X1 port map( A => B(19), ZN => n32);
   U61 : NOR2_X1 port map( A1 => n33, A2 => n32, ZN => Gout(19));
   U62 : INV_X1 port map( A => A(20), ZN => n35);
   U63 : INV_X1 port map( A => B(20), ZN => n34);
   U65 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => Gout(20));
   U66 : INV_X1 port map( A => A(21), ZN => n37);
   U67 : INV_X1 port map( A => B(21), ZN => n36);
   U68 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => Gout(21));
   U69 : INV_X1 port map( A => A(22), ZN => n39);
   U70 : INV_X1 port map( A => B(22), ZN => n38);
   U71 : NOR2_X1 port map( A1 => n39, A2 => n38, ZN => Gout(22));
   U72 : INV_X1 port map( A => A(23), ZN => n41);
   U73 : INV_X1 port map( A => B(23), ZN => n40);
   U74 : NOR2_X1 port map( A1 => n41, A2 => n40, ZN => Gout(23));
   U75 : INV_X1 port map( A => A(24), ZN => n43);
   U76 : INV_X1 port map( A => B(24), ZN => n42);
   U77 : NOR2_X1 port map( A1 => n43, A2 => n42, ZN => Gout(24));
   U78 : INV_X1 port map( A => A(25), ZN => n45);
   U79 : INV_X1 port map( A => B(25), ZN => n44);
   U80 : NOR2_X1 port map( A1 => n45, A2 => n44, ZN => Gout(25));
   U81 : INV_X1 port map( A => A(26), ZN => n47);
   U82 : INV_X1 port map( A => B(26), ZN => n46);
   U83 : NOR2_X1 port map( A1 => n47, A2 => n46, ZN => Gout(26));
   U84 : INV_X1 port map( A => A(27), ZN => n49);
   U85 : INV_X1 port map( A => B(27), ZN => n48);
   U86 : NOR2_X1 port map( A1 => n49, A2 => n48, ZN => Gout(27));
   U87 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U88 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U89 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U90 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U91 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U92 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U93 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U94 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U95 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U96 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U97 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U98 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U99 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U100 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U101 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U102 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U103 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U104 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U105 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U106 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U107 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U108 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U109 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U110 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U111 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U112 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U113 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_5;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : XNOR2_X1 port map( A => A(15), B => n32, ZN => Pout(15));
   U2 : XNOR2_X1 port map( A => n40, B => A(19), ZN => Pout(19));
   U3 : AND2_X1 port map( A1 => A(14), A2 => B(14), ZN => Gout(14));
   U4 : AND2_X1 port map( A1 => A(24), A2 => B(24), ZN => Gout(24));
   U5 : XOR2_X1 port map( A => A(24), B => B(24), Z => Pout(24));
   U6 : AND2_X1 port map( A1 => A(20), A2 => B(20), ZN => Gout(20));
   U7 : OAI21_X1 port map( B1 => n4, B2 => A(21), A => n5, ZN => Pout(21));
   U8 : XNOR2_X1 port map( A => n45, B => A(25), ZN => Pout(25));
   U9 : XNOR2_X1 port map( A => A(13), B => n30, ZN => Pout(13));
   U10 : OR2_X1 port map( A1 => A(23), A2 => n6, ZN => n8);
   U11 : OR2_X1 port map( A1 => A(27), A2 => n49, ZN => n2);
   U12 : NAND2_X1 port map( A1 => A(27), A2 => n1, ZN => n3);
   U13 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Pout(27));
   U14 : INV_X1 port map( A => B(27), ZN => n1);
   U15 : NAND2_X1 port map( A1 => A(21), A2 => n4, ZN => n5);
   U16 : INV_X1 port map( A => B(21), ZN => n4);
   U17 : NAND2_X1 port map( A1 => A(23), A2 => n6, ZN => n9);
   U18 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Pout(23));
   U19 : INV_X1 port map( A => B(23), ZN => n6);
   U20 : INV_X1 port map( A => A(23), ZN => n7);
   U21 : AND2_X1 port map( A1 => A(5), A2 => B(5), ZN => Gout(5));
   U22 : AND2_X1 port map( A1 => A(4), A2 => B(4), ZN => Gout(4));
   U23 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => Gout(0));
   U24 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U25 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U26 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U27 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U28 : INV_X1 port map( A => A(1), ZN => n11);
   U29 : INV_X1 port map( A => B(1), ZN => n10);
   U30 : NOR2_X1 port map( A1 => n11, A2 => n10, ZN => Gout(1));
   U31 : INV_X1 port map( A => A(2), ZN => n13);
   U32 : INV_X1 port map( A => B(2), ZN => n12);
   U33 : NOR2_X1 port map( A1 => n13, A2 => n12, ZN => Gout(2));
   U34 : INV_X1 port map( A => A(3), ZN => n15);
   U35 : INV_X1 port map( A => B(3), ZN => n14);
   U36 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => Gout(3));
   U37 : INV_X1 port map( A => A(6), ZN => n17);
   U38 : INV_X1 port map( A => B(6), ZN => n16);
   U39 : NOR2_X1 port map( A1 => n17, A2 => n16, ZN => Gout(6));
   U42 : INV_X1 port map( A => A(7), ZN => n19);
   U45 : INV_X1 port map( A => B(7), ZN => n18);
   U46 : NOR2_X1 port map( A1 => n19, A2 => n18, ZN => Gout(7));
   U47 : INV_X1 port map( A => A(8), ZN => n21);
   U48 : INV_X1 port map( A => B(8), ZN => n20);
   U49 : NOR2_X1 port map( A1 => n21, A2 => n20, ZN => Gout(8));
   U50 : INV_X1 port map( A => A(9), ZN => n23);
   U51 : INV_X1 port map( A => B(9), ZN => n22);
   U52 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => Gout(9));
   U53 : INV_X1 port map( A => A(10), ZN => n25);
   U54 : INV_X1 port map( A => B(10), ZN => n24);
   U55 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => Gout(10));
   U56 : INV_X1 port map( A => A(11), ZN => n27);
   U57 : INV_X1 port map( A => B(11), ZN => n26);
   U58 : NOR2_X1 port map( A1 => n27, A2 => n26, ZN => Gout(11));
   U59 : INV_X1 port map( A => A(12), ZN => n29);
   U60 : INV_X1 port map( A => B(12), ZN => n28);
   U61 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => Gout(12));
   U62 : INV_X1 port map( A => A(13), ZN => n31);
   U63 : INV_X1 port map( A => B(13), ZN => n30);
   U65 : NOR2_X1 port map( A1 => n31, A2 => n30, ZN => Gout(13));
   U66 : INV_X1 port map( A => A(15), ZN => n33);
   U67 : INV_X1 port map( A => B(15), ZN => n32);
   U68 : NOR2_X1 port map( A1 => n33, A2 => n32, ZN => Gout(15));
   U69 : INV_X1 port map( A => A(16), ZN => n35);
   U70 : INV_X1 port map( A => B(16), ZN => n34);
   U71 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => Gout(16));
   U72 : INV_X1 port map( A => A(17), ZN => n37);
   U73 : INV_X1 port map( A => B(17), ZN => n36);
   U74 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => Gout(17));
   U75 : INV_X1 port map( A => A(18), ZN => n39);
   U76 : INV_X1 port map( A => B(18), ZN => n38);
   U77 : NOR2_X1 port map( A1 => n39, A2 => n38, ZN => Gout(18));
   U78 : INV_X1 port map( A => A(19), ZN => n41);
   U79 : INV_X1 port map( A => B(19), ZN => n40);
   U80 : NOR2_X1 port map( A1 => n41, A2 => n40, ZN => Gout(19));
   U81 : INV_X1 port map( A => A(21), ZN => n42);
   U82 : NOR2_X1 port map( A1 => n42, A2 => n4, ZN => Gout(21));
   U83 : INV_X1 port map( A => A(22), ZN => n44);
   U84 : INV_X1 port map( A => B(22), ZN => n43);
   U85 : NOR2_X1 port map( A1 => n44, A2 => n43, ZN => Gout(22));
   U86 : NOR2_X1 port map( A1 => n7, A2 => n6, ZN => Gout(23));
   U87 : INV_X1 port map( A => A(25), ZN => n46);
   U88 : INV_X1 port map( A => B(25), ZN => n45);
   U89 : NOR2_X1 port map( A1 => n46, A2 => n45, ZN => Gout(25));
   U90 : INV_X1 port map( A => A(26), ZN => n48);
   U91 : INV_X1 port map( A => B(26), ZN => n47);
   U92 : NOR2_X1 port map( A1 => n48, A2 => n47, ZN => Gout(26));
   U93 : INV_X1 port map( A => A(27), ZN => n50);
   U94 : INV_X1 port map( A => B(27), ZN => n49);
   U95 : NOR2_X1 port map( A1 => n50, A2 => n49, ZN => Gout(27));
   U96 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U97 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U98 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U99 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U100 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U101 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U102 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U103 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U104 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U105 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U106 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U107 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U108 : XOR2_X1 port map( A => A(14), B => B(14), Z => Pout(14));
   U109 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U110 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U111 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U112 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U113 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U114 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_4;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U64 : XOR2_X1 port map( A => n1, B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => A(14), A2 => B(14), ZN => Gout(14));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U3 : XNOR2_X1 port map( A => B(3), B => n7, ZN => Pout(3));
   U4 : CLKBUF_X1 port map( A => B(0), Z => n1);
   U5 : AND2_X1 port map( A1 => A(4), A2 => B(4), ZN => Gout(4));
   U6 : AND2_X1 port map( A1 => A(5), A2 => B(5), ZN => Gout(5));
   U7 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U8 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U9 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U10 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U11 : INV_X1 port map( A => A(1), ZN => n3);
   U12 : INV_X1 port map( A => B(1), ZN => n2);
   U13 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Gout(1));
   U14 : INV_X1 port map( A => A(2), ZN => n5);
   U15 : INV_X1 port map( A => B(2), ZN => n4);
   U16 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Gout(2));
   U17 : INV_X1 port map( A => A(3), ZN => n7);
   U18 : INV_X1 port map( A => B(3), ZN => n6);
   U19 : NOR2_X1 port map( A1 => n7, A2 => n6, ZN => Gout(3));
   U20 : INV_X1 port map( A => A(6), ZN => n9);
   U21 : INV_X1 port map( A => B(6), ZN => n8);
   U22 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => Gout(6));
   U23 : INV_X1 port map( A => A(7), ZN => n11);
   U24 : INV_X1 port map( A => B(7), ZN => n10);
   U25 : NOR2_X1 port map( A1 => n11, A2 => n10, ZN => Gout(7));
   U26 : INV_X1 port map( A => A(8), ZN => n13);
   U27 : INV_X1 port map( A => B(8), ZN => n12);
   U28 : NOR2_X1 port map( A1 => n13, A2 => n12, ZN => Gout(8));
   U29 : INV_X1 port map( A => A(9), ZN => n15);
   U30 : INV_X1 port map( A => B(9), ZN => n14);
   U31 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => Gout(9));
   U32 : INV_X1 port map( A => A(10), ZN => n17);
   U33 : INV_X1 port map( A => B(10), ZN => n16);
   U34 : NOR2_X1 port map( A1 => n17, A2 => n16, ZN => Gout(10));
   U35 : INV_X1 port map( A => A(11), ZN => n19);
   U36 : INV_X1 port map( A => B(11), ZN => n18);
   U37 : NOR2_X1 port map( A1 => n19, A2 => n18, ZN => Gout(11));
   U38 : INV_X1 port map( A => A(12), ZN => n21);
   U39 : INV_X1 port map( A => B(12), ZN => n20);
   U42 : NOR2_X1 port map( A1 => n21, A2 => n20, ZN => Gout(12));
   U45 : INV_X1 port map( A => A(13), ZN => n23);
   U46 : INV_X1 port map( A => B(13), ZN => n22);
   U47 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => Gout(13));
   U48 : INV_X1 port map( A => A(15), ZN => n25);
   U49 : INV_X1 port map( A => B(15), ZN => n24);
   U50 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => Gout(15));
   U51 : INV_X1 port map( A => A(16), ZN => n27);
   U52 : INV_X1 port map( A => B(16), ZN => n26);
   U53 : NOR2_X1 port map( A1 => n27, A2 => n26, ZN => Gout(16));
   U54 : INV_X1 port map( A => A(17), ZN => n29);
   U55 : INV_X1 port map( A => B(17), ZN => n28);
   U56 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => Gout(17));
   U57 : INV_X1 port map( A => A(18), ZN => n31);
   U58 : INV_X1 port map( A => B(18), ZN => n30);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n30, ZN => Gout(18));
   U60 : INV_X1 port map( A => A(19), ZN => n33);
   U61 : INV_X1 port map( A => B(19), ZN => n32);
   U62 : NOR2_X1 port map( A1 => n33, A2 => n32, ZN => Gout(19));
   U63 : INV_X1 port map( A => A(20), ZN => n35);
   U65 : INV_X1 port map( A => B(20), ZN => n34);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => Gout(20));
   U67 : INV_X1 port map( A => A(21), ZN => n37);
   U68 : INV_X1 port map( A => B(21), ZN => n36);
   U69 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => Gout(21));
   U70 : INV_X1 port map( A => A(22), ZN => n39);
   U71 : INV_X1 port map( A => B(22), ZN => n38);
   U72 : NOR2_X1 port map( A1 => n39, A2 => n38, ZN => Gout(22));
   U73 : INV_X1 port map( A => A(23), ZN => n41);
   U74 : INV_X1 port map( A => B(23), ZN => n40);
   U75 : NOR2_X1 port map( A1 => n41, A2 => n40, ZN => Gout(23));
   U76 : INV_X1 port map( A => A(24), ZN => n43);
   U77 : INV_X1 port map( A => B(24), ZN => n42);
   U78 : NOR2_X1 port map( A1 => n43, A2 => n42, ZN => Gout(24));
   U79 : INV_X1 port map( A => A(25), ZN => n45);
   U80 : INV_X1 port map( A => B(25), ZN => n44);
   U81 : NOR2_X1 port map( A1 => n45, A2 => n44, ZN => Gout(25));
   U82 : INV_X1 port map( A => A(26), ZN => n47);
   U83 : INV_X1 port map( A => B(26), ZN => n46);
   U84 : NOR2_X1 port map( A1 => n47, A2 => n46, ZN => Gout(26));
   U85 : INV_X1 port map( A => A(27), ZN => n49);
   U86 : INV_X1 port map( A => B(27), ZN => n48);
   U87 : NOR2_X1 port map( A1 => n49, A2 => n48, ZN => Gout(27));
   U88 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U89 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U90 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U91 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U92 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U93 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U94 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U95 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U96 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U97 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U98 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U99 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U100 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U101 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U102 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U103 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U104 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U105 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U106 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U107 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U108 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U109 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U110 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U111 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U112 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U113 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_3;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => A(14), A2 => B(14), ZN => Gout(14));
   U2 : XNOR2_X1 port map( A => n34, B => A(19), ZN => Pout(19));
   U3 : XNOR2_X1 port map( A => A(9), B => n16, ZN => Pout(9));
   U4 : XNOR2_X1 port map( A => A(21), B => n38, ZN => Pout(21));
   U5 : XNOR2_X1 port map( A => n48, B => A(27), ZN => Pout(27));
   U6 : INV_X1 port map( A => B(23), ZN => n1);
   U7 : AND2_X1 port map( A1 => A(23), A2 => B(23), ZN => Gout(23));
   U8 : OR2_X1 port map( A1 => A(23), A2 => n1, ZN => n2);
   U9 : NAND2_X1 port map( A1 => A(23), A2 => n1, ZN => n3);
   U10 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Pout(23));
   U11 : AND2_X1 port map( A1 => A(5), A2 => B(5), ZN => Gout(5));
   U12 : AND2_X1 port map( A1 => A(4), A2 => B(4), ZN => Gout(4));
   U13 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => Gout(0));
   U14 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U15 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U16 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U17 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U18 : INV_X1 port map( A => A(1), ZN => n5);
   U19 : INV_X1 port map( A => B(1), ZN => n4);
   U20 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Gout(1));
   U21 : INV_X1 port map( A => A(2), ZN => n7);
   U22 : INV_X1 port map( A => B(2), ZN => n6);
   U23 : NOR2_X1 port map( A1 => n7, A2 => n6, ZN => Gout(2));
   U24 : INV_X1 port map( A => A(3), ZN => n9);
   U25 : INV_X1 port map( A => B(3), ZN => n8);
   U26 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => Gout(3));
   U27 : INV_X1 port map( A => A(6), ZN => n11);
   U28 : INV_X1 port map( A => B(6), ZN => n10);
   U29 : NOR2_X1 port map( A1 => n11, A2 => n10, ZN => Gout(6));
   U30 : INV_X1 port map( A => A(7), ZN => n13);
   U31 : INV_X1 port map( A => B(7), ZN => n12);
   U32 : NOR2_X1 port map( A1 => n13, A2 => n12, ZN => Gout(7));
   U33 : INV_X1 port map( A => A(8), ZN => n15);
   U34 : INV_X1 port map( A => B(8), ZN => n14);
   U35 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => Gout(8));
   U36 : INV_X1 port map( A => A(9), ZN => n17);
   U37 : INV_X1 port map( A => B(9), ZN => n16);
   U38 : NOR2_X1 port map( A1 => n17, A2 => n16, ZN => Gout(9));
   U39 : INV_X1 port map( A => A(10), ZN => n19);
   U42 : INV_X1 port map( A => B(10), ZN => n18);
   U45 : NOR2_X1 port map( A1 => n19, A2 => n18, ZN => Gout(10));
   U46 : INV_X1 port map( A => A(11), ZN => n21);
   U47 : INV_X1 port map( A => B(11), ZN => n20);
   U48 : NOR2_X1 port map( A1 => n21, A2 => n20, ZN => Gout(11));
   U49 : INV_X1 port map( A => A(12), ZN => n23);
   U50 : INV_X1 port map( A => B(12), ZN => n22);
   U51 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => Gout(12));
   U52 : INV_X1 port map( A => A(13), ZN => n25);
   U53 : INV_X1 port map( A => B(13), ZN => n24);
   U54 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => Gout(13));
   U55 : INV_X1 port map( A => A(15), ZN => n27);
   U56 : INV_X1 port map( A => B(15), ZN => n26);
   U57 : NOR2_X1 port map( A1 => n27, A2 => n26, ZN => Gout(15));
   U58 : INV_X1 port map( A => A(16), ZN => n29);
   U59 : INV_X1 port map( A => B(16), ZN => n28);
   U60 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => Gout(16));
   U61 : INV_X1 port map( A => A(17), ZN => n31);
   U62 : INV_X1 port map( A => B(17), ZN => n30);
   U63 : NOR2_X1 port map( A1 => n31, A2 => n30, ZN => Gout(17));
   U65 : INV_X1 port map( A => A(18), ZN => n33);
   U66 : INV_X1 port map( A => B(18), ZN => n32);
   U67 : NOR2_X1 port map( A1 => n33, A2 => n32, ZN => Gout(18));
   U68 : INV_X1 port map( A => A(19), ZN => n35);
   U69 : INV_X1 port map( A => B(19), ZN => n34);
   U70 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => Gout(19));
   U71 : INV_X1 port map( A => A(20), ZN => n37);
   U72 : INV_X1 port map( A => B(20), ZN => n36);
   U73 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => Gout(20));
   U74 : INV_X1 port map( A => A(21), ZN => n39);
   U75 : INV_X1 port map( A => B(21), ZN => n38);
   U76 : NOR2_X1 port map( A1 => n39, A2 => n38, ZN => Gout(21));
   U77 : INV_X1 port map( A => A(22), ZN => n41);
   U78 : INV_X1 port map( A => B(22), ZN => n40);
   U79 : NOR2_X1 port map( A1 => n41, A2 => n40, ZN => Gout(22));
   U80 : INV_X1 port map( A => A(24), ZN => n43);
   U81 : INV_X1 port map( A => B(24), ZN => n42);
   U82 : NOR2_X1 port map( A1 => n43, A2 => n42, ZN => Gout(24));
   U83 : INV_X1 port map( A => A(25), ZN => n45);
   U84 : INV_X1 port map( A => B(25), ZN => n44);
   U85 : NOR2_X1 port map( A1 => n45, A2 => n44, ZN => Gout(25));
   U86 : INV_X1 port map( A => A(26), ZN => n47);
   U87 : INV_X1 port map( A => B(26), ZN => n46);
   U88 : NOR2_X1 port map( A1 => n47, A2 => n46, ZN => Gout(26));
   U89 : INV_X1 port map( A => A(27), ZN => n49);
   U90 : INV_X1 port map( A => B(27), ZN => n48);
   U91 : NOR2_X1 port map( A1 => n49, A2 => n48, ZN => Gout(27));
   U92 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U93 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U94 : XOR2_X1 port map( A => A(3), B => B(3), Z => Pout(3));
   U95 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U96 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U97 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U98 : XOR2_X1 port map( A => A(7), B => B(7), Z => Pout(7));
   U99 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U100 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U101 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U102 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U103 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U104 : XOR2_X1 port map( A => A(14), B => B(14), Z => Pout(14));
   U105 : XOR2_X1 port map( A => A(15), B => B(15), Z => Pout(15));
   U106 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U107 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U108 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U109 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U110 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U111 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U112 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U113 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_2;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => A(4), A2 => B(4), ZN => Gout(4));
   U2 : AND2_X1 port map( A1 => A(5), A2 => B(5), ZN => Gout(5));
   U3 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U4 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U5 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U6 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U7 : INV_X1 port map( A => A(0), ZN => n2);
   U8 : INV_X1 port map( A => B(0), ZN => n1);
   U9 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Gout(0));
   U10 : INV_X1 port map( A => A(1), ZN => n4);
   U11 : INV_X1 port map( A => B(1), ZN => n3);
   U12 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Gout(1));
   U13 : INV_X1 port map( A => A(2), ZN => n6);
   U14 : INV_X1 port map( A => B(2), ZN => n5);
   U15 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Gout(2));
   U16 : INV_X1 port map( A => A(3), ZN => n8);
   U17 : INV_X1 port map( A => B(3), ZN => n7);
   U18 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => Gout(3));
   U19 : INV_X1 port map( A => A(6), ZN => n10);
   U20 : INV_X1 port map( A => B(6), ZN => n9);
   U21 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => Gout(6));
   U22 : INV_X1 port map( A => A(7), ZN => n12);
   U23 : INV_X1 port map( A => B(7), ZN => n11);
   U24 : NOR2_X1 port map( A1 => n12, A2 => n11, ZN => Gout(7));
   U25 : INV_X1 port map( A => A(8), ZN => n14);
   U26 : INV_X1 port map( A => B(8), ZN => n13);
   U27 : NOR2_X1 port map( A1 => n14, A2 => n13, ZN => Gout(8));
   U28 : INV_X1 port map( A => A(9), ZN => n16);
   U29 : INV_X1 port map( A => B(9), ZN => n15);
   U30 : NOR2_X1 port map( A1 => n16, A2 => n15, ZN => Gout(9));
   U31 : INV_X1 port map( A => A(10), ZN => n18);
   U32 : INV_X1 port map( A => B(10), ZN => n17);
   U33 : NOR2_X1 port map( A1 => n18, A2 => n17, ZN => Gout(10));
   U34 : INV_X1 port map( A => A(11), ZN => n20);
   U35 : INV_X1 port map( A => B(11), ZN => n19);
   U36 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => Gout(11));
   U37 : INV_X1 port map( A => A(12), ZN => n22);
   U38 : INV_X1 port map( A => B(12), ZN => n21);
   U39 : NOR2_X1 port map( A1 => n22, A2 => n21, ZN => Gout(12));
   U42 : INV_X1 port map( A => A(13), ZN => n24);
   U45 : INV_X1 port map( A => B(13), ZN => n23);
   U46 : NOR2_X1 port map( A1 => n24, A2 => n23, ZN => Gout(13));
   U47 : INV_X1 port map( A => A(14), ZN => n26);
   U48 : INV_X1 port map( A => B(14), ZN => n25);
   U49 : NOR2_X1 port map( A1 => n26, A2 => n25, ZN => Gout(14));
   U50 : INV_X1 port map( A => A(15), ZN => n28);
   U51 : INV_X1 port map( A => B(15), ZN => n27);
   U52 : NOR2_X1 port map( A1 => n28, A2 => n27, ZN => Gout(15));
   U53 : INV_X1 port map( A => A(16), ZN => n30);
   U54 : INV_X1 port map( A => B(16), ZN => n29);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n29, ZN => Gout(16));
   U56 : INV_X1 port map( A => A(17), ZN => n32);
   U57 : INV_X1 port map( A => B(17), ZN => n31);
   U58 : NOR2_X1 port map( A1 => n32, A2 => n31, ZN => Gout(17));
   U59 : INV_X1 port map( A => A(18), ZN => n34);
   U60 : INV_X1 port map( A => B(18), ZN => n33);
   U61 : NOR2_X1 port map( A1 => n34, A2 => n33, ZN => Gout(18));
   U62 : INV_X1 port map( A => A(19), ZN => n36);
   U63 : INV_X1 port map( A => B(19), ZN => n35);
   U65 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => Gout(19));
   U66 : INV_X1 port map( A => A(20), ZN => n38);
   U67 : INV_X1 port map( A => B(20), ZN => n37);
   U68 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => Gout(20));
   U69 : INV_X1 port map( A => A(21), ZN => n40);
   U70 : INV_X1 port map( A => B(21), ZN => n39);
   U71 : NOR2_X1 port map( A1 => n40, A2 => n39, ZN => Gout(21));
   U72 : INV_X1 port map( A => A(22), ZN => n42);
   U73 : INV_X1 port map( A => B(22), ZN => n41);
   U74 : NOR2_X1 port map( A1 => n42, A2 => n41, ZN => Gout(22));
   U75 : INV_X1 port map( A => A(23), ZN => n44);
   U76 : INV_X1 port map( A => B(23), ZN => n43);
   U77 : NOR2_X1 port map( A1 => n44, A2 => n43, ZN => Gout(23));
   U78 : INV_X1 port map( A => A(24), ZN => n46);
   U79 : INV_X1 port map( A => B(24), ZN => n45);
   U80 : NOR2_X1 port map( A1 => n46, A2 => n45, ZN => Gout(24));
   U81 : INV_X1 port map( A => A(25), ZN => n48);
   U82 : INV_X1 port map( A => B(25), ZN => n47);
   U83 : NOR2_X1 port map( A1 => n48, A2 => n47, ZN => Gout(25));
   U84 : INV_X1 port map( A => A(26), ZN => n50);
   U85 : INV_X1 port map( A => B(26), ZN => n49);
   U86 : NOR2_X1 port map( A1 => n50, A2 => n49, ZN => Gout(26));
   U87 : INV_X1 port map( A => A(27), ZN => n52);
   U88 : INV_X1 port map( A => B(27), ZN => n51);
   U89 : NOR2_X1 port map( A1 => n52, A2 => n51, ZN => Gout(27));
   U90 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U91 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U92 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U93 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U94 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U95 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U96 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U97 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U98 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U99 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U100 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U101 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U102 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U103 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U104 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U105 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U106 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U107 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U108 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U109 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U110 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U111 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U112 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U113 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U114 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U115 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U116 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_1;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50 : std_logic;

begin
   
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => A(4), A2 => B(4), ZN => Gout(4));
   U2 : AND2_X1 port map( A1 => A(5), A2 => B(5), ZN => Gout(5));
   U3 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => Gout(0));
   U4 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U5 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U6 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U7 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U8 : INV_X1 port map( A => A(1), ZN => n2);
   U9 : INV_X1 port map( A => B(1), ZN => n1);
   U10 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Gout(1));
   U11 : INV_X1 port map( A => A(2), ZN => n4);
   U12 : INV_X1 port map( A => B(2), ZN => n3);
   U13 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Gout(2));
   U14 : INV_X1 port map( A => A(3), ZN => n6);
   U15 : INV_X1 port map( A => B(3), ZN => n5);
   U16 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Gout(3));
   U17 : INV_X1 port map( A => A(6), ZN => n8);
   U18 : INV_X1 port map( A => B(6), ZN => n7);
   U19 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => Gout(6));
   U20 : INV_X1 port map( A => A(7), ZN => n10);
   U21 : INV_X1 port map( A => B(7), ZN => n9);
   U22 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => Gout(7));
   U23 : INV_X1 port map( A => A(8), ZN => n12);
   U24 : INV_X1 port map( A => B(8), ZN => n11);
   U25 : NOR2_X1 port map( A1 => n12, A2 => n11, ZN => Gout(8));
   U26 : INV_X1 port map( A => A(9), ZN => n14);
   U27 : INV_X1 port map( A => B(9), ZN => n13);
   U28 : NOR2_X1 port map( A1 => n14, A2 => n13, ZN => Gout(9));
   U29 : INV_X1 port map( A => A(10), ZN => n16);
   U30 : INV_X1 port map( A => B(10), ZN => n15);
   U31 : NOR2_X1 port map( A1 => n16, A2 => n15, ZN => Gout(10));
   U32 : INV_X1 port map( A => A(11), ZN => n18);
   U33 : INV_X1 port map( A => B(11), ZN => n17);
   U34 : NOR2_X1 port map( A1 => n18, A2 => n17, ZN => Gout(11));
   U35 : INV_X1 port map( A => A(12), ZN => n20);
   U36 : INV_X1 port map( A => B(12), ZN => n19);
   U37 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => Gout(12));
   U38 : INV_X1 port map( A => A(13), ZN => n22);
   U39 : INV_X1 port map( A => B(13), ZN => n21);
   U42 : NOR2_X1 port map( A1 => n22, A2 => n21, ZN => Gout(13));
   U45 : INV_X1 port map( A => A(14), ZN => n24);
   U46 : INV_X1 port map( A => B(14), ZN => n23);
   U47 : NOR2_X1 port map( A1 => n24, A2 => n23, ZN => Gout(14));
   U48 : INV_X1 port map( A => A(15), ZN => n26);
   U49 : INV_X1 port map( A => B(15), ZN => n25);
   U50 : NOR2_X1 port map( A1 => n26, A2 => n25, ZN => Gout(15));
   U51 : INV_X1 port map( A => A(16), ZN => n28);
   U52 : INV_X1 port map( A => B(16), ZN => n27);
   U53 : NOR2_X1 port map( A1 => n28, A2 => n27, ZN => Gout(16));
   U54 : INV_X1 port map( A => A(17), ZN => n30);
   U55 : INV_X1 port map( A => B(17), ZN => n29);
   U56 : NOR2_X1 port map( A1 => n30, A2 => n29, ZN => Gout(17));
   U57 : INV_X1 port map( A => A(18), ZN => n32);
   U58 : INV_X1 port map( A => B(18), ZN => n31);
   U59 : NOR2_X1 port map( A1 => n32, A2 => n31, ZN => Gout(18));
   U60 : INV_X1 port map( A => A(19), ZN => n34);
   U61 : INV_X1 port map( A => B(19), ZN => n33);
   U62 : NOR2_X1 port map( A1 => n34, A2 => n33, ZN => Gout(19));
   U63 : INV_X1 port map( A => A(20), ZN => n36);
   U65 : INV_X1 port map( A => B(20), ZN => n35);
   U66 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => Gout(20));
   U67 : INV_X1 port map( A => A(21), ZN => n38);
   U68 : INV_X1 port map( A => B(21), ZN => n37);
   U69 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => Gout(21));
   U70 : INV_X1 port map( A => A(22), ZN => n40);
   U71 : INV_X1 port map( A => B(22), ZN => n39);
   U72 : NOR2_X1 port map( A1 => n40, A2 => n39, ZN => Gout(22));
   U73 : INV_X1 port map( A => A(23), ZN => n42);
   U74 : INV_X1 port map( A => B(23), ZN => n41);
   U75 : NOR2_X1 port map( A1 => n42, A2 => n41, ZN => Gout(23));
   U76 : INV_X1 port map( A => A(24), ZN => n44);
   U77 : INV_X1 port map( A => B(24), ZN => n43);
   U78 : NOR2_X1 port map( A1 => n44, A2 => n43, ZN => Gout(24));
   U79 : INV_X1 port map( A => A(25), ZN => n46);
   U80 : INV_X1 port map( A => B(25), ZN => n45);
   U81 : NOR2_X1 port map( A1 => n46, A2 => n45, ZN => Gout(25));
   U82 : INV_X1 port map( A => A(26), ZN => n48);
   U83 : INV_X1 port map( A => B(26), ZN => n47);
   U84 : NOR2_X1 port map( A1 => n48, A2 => n47, ZN => Gout(26));
   U85 : INV_X1 port map( A => A(27), ZN => n50);
   U86 : INV_X1 port map( A => B(27), ZN => n49);
   U87 : NOR2_X1 port map( A1 => n50, A2 => n49, ZN => Gout(27));
   U88 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U89 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U90 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U91 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U92 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U93 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U94 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U95 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U96 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U97 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U98 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U99 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U100 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U101 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U102 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U103 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U104 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U105 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U106 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U107 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U108 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U109 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U110 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U111 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U112 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U113 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U114 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_7 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_7;

architecture SYN_BEHAVIORAL of ENCODER_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_6 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_6;

architecture SYN_BEHAVIORAL of ENCODER_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_5 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_5;

architecture SYN_BEHAVIORAL of ENCODER_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_4 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_4;

architecture SYN_BEHAVIORAL of ENCODER_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_3 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_3;

architecture SYN_BEHAVIORAL of ENCODER_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_2 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_2;

architecture SYN_BEHAVIORAL of ENCODER_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_1 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_1;

architecture SYN_BEHAVIORAL of ENCODER_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_31 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_31;

architecture SYN_ARCH1 of ND4_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_30 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_30;

architecture SYN_ARCH1 of ND4_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_29 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_29;

architecture SYN_ARCH1 of ND4_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_28 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_28;

architecture SYN_ARCH1 of ND4_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_27 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_27;

architecture SYN_ARCH1 of ND4_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_26 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_26;

architecture SYN_ARCH1 of ND4_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_25 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_25;

architecture SYN_ARCH1 of ND4_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_24 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_24;

architecture SYN_ARCH1 of ND4_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_23 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_23;

architecture SYN_ARCH1 of ND4_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_22 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_22;

architecture SYN_ARCH1 of ND4_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_21 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_21;

architecture SYN_ARCH1 of ND4_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_20 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_20;

architecture SYN_ARCH1 of ND4_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_19 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_19;

architecture SYN_ARCH1 of ND4_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_18 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_18;

architecture SYN_ARCH1 of ND4_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_17 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_17;

architecture SYN_ARCH1 of ND4_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_16 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_16;

architecture SYN_ARCH1 of ND4_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_15 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_15;

architecture SYN_ARCH1 of ND4_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_14 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_14;

architecture SYN_ARCH1 of ND4_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_13 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_13;

architecture SYN_ARCH1 of ND4_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_12 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_12;

architecture SYN_ARCH1 of ND4_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_11 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_11;

architecture SYN_ARCH1 of ND4_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_10 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_10;

architecture SYN_ARCH1 of ND4_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_9 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_9;

architecture SYN_ARCH1 of ND4_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_8 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_8;

architecture SYN_ARCH1 of ND4_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_7 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_7;

architecture SYN_ARCH1 of ND4_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_6 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_6;

architecture SYN_ARCH1 of ND4_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_5 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_5;

architecture SYN_ARCH1 of ND4_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_4 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_4;

architecture SYN_ARCH1 of ND4_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_3 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_3;

architecture SYN_ARCH1 of ND4_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_2 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_2;

architecture SYN_ARCH1 of ND4_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_1 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_1;

architecture SYN_ARCH1 of ND4_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_127 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_127;

architecture SYN_ARCH1 of ND3_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_126 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_126;

architecture SYN_ARCH1 of ND3_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_125 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_125;

architecture SYN_ARCH1 of ND3_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_124 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_124;

architecture SYN_ARCH1 of ND3_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_123 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_123;

architecture SYN_ARCH1 of ND3_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_122 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_122;

architecture SYN_ARCH1 of ND3_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_121 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_121;

architecture SYN_ARCH1 of ND3_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_120 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_120;

architecture SYN_ARCH1 of ND3_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_119 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_119;

architecture SYN_ARCH1 of ND3_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_118 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_118;

architecture SYN_ARCH1 of ND3_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_117 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_117;

architecture SYN_ARCH1 of ND3_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_116 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_116;

architecture SYN_ARCH1 of ND3_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_115 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_115;

architecture SYN_ARCH1 of ND3_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_114 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_114;

architecture SYN_ARCH1 of ND3_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_113 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_113;

architecture SYN_ARCH1 of ND3_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_112 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_112;

architecture SYN_ARCH1 of ND3_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_111 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_111;

architecture SYN_ARCH1 of ND3_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_110 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_110;

architecture SYN_ARCH1 of ND3_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_109 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_109;

architecture SYN_ARCH1 of ND3_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_108 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_108;

architecture SYN_ARCH1 of ND3_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_107 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_107;

architecture SYN_ARCH1 of ND3_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_106 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_106;

architecture SYN_ARCH1 of ND3_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_105 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_105;

architecture SYN_ARCH1 of ND3_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_104 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_104;

architecture SYN_ARCH1 of ND3_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_103 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_103;

architecture SYN_ARCH1 of ND3_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_102 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_102;

architecture SYN_ARCH1 of ND3_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_101 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_101;

architecture SYN_ARCH1 of ND3_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_100 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_100;

architecture SYN_ARCH1 of ND3_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_99 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_99;

architecture SYN_ARCH1 of ND3_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_98 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_98;

architecture SYN_ARCH1 of ND3_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_97 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_97;

architecture SYN_ARCH1 of ND3_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_96 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_96;

architecture SYN_ARCH1 of ND3_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_95 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_95;

architecture SYN_ARCH1 of ND3_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_94 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_94;

architecture SYN_ARCH1 of ND3_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_93 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_93;

architecture SYN_ARCH1 of ND3_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_92 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_92;

architecture SYN_ARCH1 of ND3_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_91 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_91;

architecture SYN_ARCH1 of ND3_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_90 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_90;

architecture SYN_ARCH1 of ND3_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_89 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_89;

architecture SYN_ARCH1 of ND3_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_88 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_88;

architecture SYN_ARCH1 of ND3_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_87 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_87;

architecture SYN_ARCH1 of ND3_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_86 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_86;

architecture SYN_ARCH1 of ND3_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_85 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_85;

architecture SYN_ARCH1 of ND3_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_84 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_84;

architecture SYN_ARCH1 of ND3_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_83 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_83;

architecture SYN_ARCH1 of ND3_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_82 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_82;

architecture SYN_ARCH1 of ND3_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_81 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_81;

architecture SYN_ARCH1 of ND3_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_80 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_80;

architecture SYN_ARCH1 of ND3_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_79 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_79;

architecture SYN_ARCH1 of ND3_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_78 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_78;

architecture SYN_ARCH1 of ND3_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_77 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_77;

architecture SYN_ARCH1 of ND3_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_76 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_76;

architecture SYN_ARCH1 of ND3_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_75 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_75;

architecture SYN_ARCH1 of ND3_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_74 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_74;

architecture SYN_ARCH1 of ND3_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_73 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_73;

architecture SYN_ARCH1 of ND3_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_72 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_72;

architecture SYN_ARCH1 of ND3_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_71 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_71;

architecture SYN_ARCH1 of ND3_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_70 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_70;

architecture SYN_ARCH1 of ND3_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_69 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_69;

architecture SYN_ARCH1 of ND3_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_68 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_68;

architecture SYN_ARCH1 of ND3_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_67 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_67;

architecture SYN_ARCH1 of ND3_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_66 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_66;

architecture SYN_ARCH1 of ND3_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_65 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_65;

architecture SYN_ARCH1 of ND3_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_64 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_64;

architecture SYN_ARCH1 of ND3_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_63 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_63;

architecture SYN_ARCH1 of ND3_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_62 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_62;

architecture SYN_ARCH1 of ND3_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_61 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_61;

architecture SYN_ARCH1 of ND3_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_60 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_60;

architecture SYN_ARCH1 of ND3_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_59 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_59;

architecture SYN_ARCH1 of ND3_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_58 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_58;

architecture SYN_ARCH1 of ND3_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_57 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_57;

architecture SYN_ARCH1 of ND3_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_56 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_56;

architecture SYN_ARCH1 of ND3_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_55 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_55;

architecture SYN_ARCH1 of ND3_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_54 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_54;

architecture SYN_ARCH1 of ND3_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_53 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_53;

architecture SYN_ARCH1 of ND3_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_52 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_52;

architecture SYN_ARCH1 of ND3_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_51 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_51;

architecture SYN_ARCH1 of ND3_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_50 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_50;

architecture SYN_ARCH1 of ND3_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_49 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_49;

architecture SYN_ARCH1 of ND3_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_48 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_48;

architecture SYN_ARCH1 of ND3_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_47 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_47;

architecture SYN_ARCH1 of ND3_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_46 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_46;

architecture SYN_ARCH1 of ND3_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_45 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_45;

architecture SYN_ARCH1 of ND3_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_44 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_44;

architecture SYN_ARCH1 of ND3_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_43 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_43;

architecture SYN_ARCH1 of ND3_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_42 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_42;

architecture SYN_ARCH1 of ND3_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_41 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_41;

architecture SYN_ARCH1 of ND3_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_40 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_40;

architecture SYN_ARCH1 of ND3_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_39 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_39;

architecture SYN_ARCH1 of ND3_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_38 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_38;

architecture SYN_ARCH1 of ND3_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_37 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_37;

architecture SYN_ARCH1 of ND3_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_36 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_36;

architecture SYN_ARCH1 of ND3_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_35 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_35;

architecture SYN_ARCH1 of ND3_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_34 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_34;

architecture SYN_ARCH1 of ND3_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_33 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_33;

architecture SYN_ARCH1 of ND3_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_32 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_32;

architecture SYN_ARCH1 of ND3_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_31 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_31;

architecture SYN_ARCH1 of ND3_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_30 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_30;

architecture SYN_ARCH1 of ND3_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_29 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_29;

architecture SYN_ARCH1 of ND3_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_28 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_28;

architecture SYN_ARCH1 of ND3_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_27 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_27;

architecture SYN_ARCH1 of ND3_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_26 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_26;

architecture SYN_ARCH1 of ND3_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_25 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_25;

architecture SYN_ARCH1 of ND3_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_24 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_24;

architecture SYN_ARCH1 of ND3_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_23 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_23;

architecture SYN_ARCH1 of ND3_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_22 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_22;

architecture SYN_ARCH1 of ND3_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_21 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_21;

architecture SYN_ARCH1 of ND3_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_20 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_20;

architecture SYN_ARCH1 of ND3_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_19 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_19;

architecture SYN_ARCH1 of ND3_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_18 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_18;

architecture SYN_ARCH1 of ND3_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_17 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_17;

architecture SYN_ARCH1 of ND3_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_16 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_16;

architecture SYN_ARCH1 of ND3_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_15 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_15;

architecture SYN_ARCH1 of ND3_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_14 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_14;

architecture SYN_ARCH1 of ND3_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_13 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_13;

architecture SYN_ARCH1 of ND3_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_12 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_12;

architecture SYN_ARCH1 of ND3_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_11 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_11;

architecture SYN_ARCH1 of ND3_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_10 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_10;

architecture SYN_ARCH1 of ND3_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_9 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_9;

architecture SYN_ARCH1 of ND3_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_8 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_8;

architecture SYN_ARCH1 of ND3_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_7 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_7;

architecture SYN_ARCH1 of ND3_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_6 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_6;

architecture SYN_ARCH1 of ND3_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_5 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_5;

architecture SYN_ARCH1 of ND3_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_4 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_4;

architecture SYN_ARCH1 of ND3_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_3 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_3;

architecture SYN_ARCH1 of ND3_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_2 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_2;

architecture SYN_ARCH1 of ND3_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_1 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_1;

architecture SYN_ARCH1 of ND3_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 is

   component CARRY_SEL_N_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_55 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_54 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_53 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_52 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_51 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_50 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_49 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 is

   component CARRY_SEL_N_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_47 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_46 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_45 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_44 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_43 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_42 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_41 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 is

   component CARRY_SEL_N_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_39 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_38 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_37 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_36 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_35 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_34 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_33 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 is

   component CARRY_SEL_N_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_31 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_30 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_29 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_28 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_27 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_26 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_25 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 is

   component CARRY_SEL_N_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_23 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_22 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_21 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_20 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_19 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_18 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_17 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 is

   component CARRY_SEL_N_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_15 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_14 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_13 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_12 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_11 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_10 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_9 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 is

   component CARRY_SEL_N_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_55
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_56
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_57
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_58
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_163
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_164
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_59
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_60
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_165
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_166
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_167
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_61
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_168
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_169
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_170
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_171
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_172
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_173
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_174
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_62
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_175
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_176
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_177
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_178
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_179
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_180
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_181
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_182
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_183
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_184
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_185
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_186
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_187
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_188
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_189
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_63
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n2, n3, n4, n5, n6, n_1154 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n6);
   pgnetwork_0 : PG_network_NBIT32_7 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1154, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_63 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_189 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_188 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_187 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_186 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_185 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_184 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_183 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_182 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_181 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_180 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_179 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_178 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_177 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_176 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_175 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_62 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_174 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_173 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_172 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_171 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_170 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_169 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_168 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_61 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_167 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_166 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_165 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_60 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_59 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_164 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_163 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_58 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_57 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_56 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_55 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Cin, A2 => n6, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => n4, A2 => n5, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_46
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_47
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_48
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_49
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_136
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_137
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_50
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_51
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_138
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_139
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_140
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_52
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_141
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_142
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_143
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_144
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_145
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_146
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_147
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_53
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_148
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_149
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_150
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_151
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_152
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_153
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_154
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_155
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_156
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_157
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_158
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_159
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_160
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_161
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_162
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_54
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, n11, Co_3_port, n12, n13,
      G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, G_16_9_port, 
      G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, G_12_12_port, 
      G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, G_10_9_port, 
      G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, G_6_6_port, 
      G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, G_2_2_port, 
      G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, G_32_25_port, 
      G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, G_29_29_port, 
      G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, G_27_27_port, 
      G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, G_24_23_port, 
      G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, G_22_21_port, 
      G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, G_19_19_port, 
      G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, P_32_32_port, P_32_31_port, P_32_29_port, 
      P_32_25_port, P_32_17_port, P_31_31_port, P_30_30_port, P_30_29_port, 
      P_29_29_port, P_28_28_port, P_28_27_port, P_28_25_port, P_28_17_port, 
      P_27_27_port, P_26_26_port, P_26_25_port, P_25_25_port, P_24_24_port, 
      P_24_23_port, P_24_21_port, P_24_17_port, P_23_23_port, P_22_22_port, 
      P_22_21_port, P_21_21_port, P_20_20_port, P_20_19_port, P_20_17_port, 
      P_19_19_port, P_18_18_port, P_18_17_port, P_17_17_port, n1, n2, Co_1_port
      , Co_4_port, Co_2_port, n6, n7, n8, n9, n10, n_1155 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_6 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => n2, Pout(31) => P_32_32_port, Pout(30)
                           => P_31_31_port, Pout(29) => P_30_30_port, Pout(28) 
                           => P_29_29_port, Pout(27) => P_28_28_port, Pout(26) 
                           => P_27_27_port, Pout(25) => P_26_26_port, Pout(24) 
                           => P_25_25_port, Pout(23) => P_24_24_port, Pout(22) 
                           => P_23_23_port, Pout(21) => P_22_22_port, Pout(20) 
                           => P_21_21_port, Pout(19) => P_20_20_port, Pout(18) 
                           => P_19_19_port, Pout(17) => P_18_18_port, Pout(16) 
                           => P_17_17_port, Pout(15) => P_16_16_port, Pout(14) 
                           => P_15_15_port, Pout(13) => P_14_14_port, Pout(12) 
                           => P_13_13_port, Pout(11) => P_12_12_port, Pout(10) 
                           => P_11_11_port, Pout(9) => P_10_10_port, Pout(8) =>
                           P_9_9_port, Pout(7) => P_8_8_port, Pout(6) => 
                           P_7_7_port, Pout(5) => P_6_6_port, Pout(4) => 
                           P_5_5_port, Pout(3) => P_4_4_port, Pout(2) => 
                           P_3_3_port, Pout(1) => P_2_2_port, Pout(0) => n_1155
                           , Gout(31) => G_32_32_port, Gout(30) => G_31_31_port
                           , Gout(29) => G_30_30_port, Gout(28) => G_29_29_port
                           , Gout(27) => G_28_28_port, Gout(26) => G_27_27_port
                           , Gout(25) => G_26_26_port, Gout(24) => G_25_25_port
                           , Gout(23) => G_24_24_port, Gout(22) => G_23_23_port
                           , Gout(21) => G_22_22_port, Gout(20) => G_21_21_port
                           , Gout(19) => G_20_20_port, Gout(18) => G_19_19_port
                           , Gout(17) => G_18_18_port, Gout(16) => G_17_17_port
                           , Gout(15) => G_16_16_port, Gout(14) => G_15_15_port
                           , Gout(13) => G_14_14_port, Gout(12) => G_13_13_port
                           , Gout(11) => G_12_12_port, Gout(10) => G_11_11_port
                           , Gout(9) => G_10_10_port, Gout(8) => G_9_9_port, 
                           Gout(7) => G_8_8_port, Gout(6) => G_7_7_port, 
                           Gout(5) => G_6_6_port, Gout(4) => G_5_5_port, 
                           Gout(3) => G_4_4_port, Gout(2) => G_3_3_port, 
                           Gout(1) => G_2_2_port, Gout(0) => n10);
   gblock1_1_1 : G_block_54 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_162 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_161 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_160 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_159 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_158 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_157 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_156 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_155 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_154 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_153 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_152 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_151 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_150 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_149 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_148 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_53 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => n13);
   pgblock1_2_2 : PG_block_147 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_146 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_145 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_144 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_143 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_142 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_141 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_52 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => n13, Gout => n12);
   pgblock1_3_2 : PG_block_140 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_139 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_138 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_51 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_50 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => n12, Gout => n11);
   pgblock2_4_28_2 : PG_block_137 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_136 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_49 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => n11, Gout => Co_5_port);
   gblock2_5_6 : G_block_48 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_47 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => n1, Gout => Co_7_port);
   gblock2_5_8 : G_block_46 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => n1, Gout => Co_8_port);
   U1 : CLKBUF_X3 port map( A => n11, Z => Co_4_port);
   U2 : BUF_X2 port map( A => n12, Z => Co_2_port);
   U3 : CLKBUF_X1 port map( A => B(0), Z => n2);
   U4 : CLKBUF_X1 port map( A => Co_4_port, Z => n1);
   U5 : CLKBUF_X1 port map( A => n13, Z => Co_1_port);
   U6 : INV_X1 port map( A => Cin, ZN => n8);
   U7 : INV_X1 port map( A => B(0), ZN => n7);
   U8 : INV_X1 port map( A => A(0), ZN => n6);
   U9 : OAI222_X1 port map( A1 => n8, A2 => n7, B1 => n6, B2 => n8, C1 => n7, 
                           C2 => n6, ZN => n9);
   U10 : AND2_X1 port map( A1 => n9, A2 => n10, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_37
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_38
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_39
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_40
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_109
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_110
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_41
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_42
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_111
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_112
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_113
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_43
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_114
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_115
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_116
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_117
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_118
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_119
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_120
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_44
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_121
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_122
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_123
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_124
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_125
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_126
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_127
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_128
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_129
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_130
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_131
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_132
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_133
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_134
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_135
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_45
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, n10, Co_3_port, Co_2_port
      , Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, 
      P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, 
      P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, 
      P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, 
      P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, 
      P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n1, Co_4_port, n3, n4, n5, n6, n7, n8, n9, n_1156 : 
      std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_5 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1156, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n9);
   gblock1_1_1 : G_block_45 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_135 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_134 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_133 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_132 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_131 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_130 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_129 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_128 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_127 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_126 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_125 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_124 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_123 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_122 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_121 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_44 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_120 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_119 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_118 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_117 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_116 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_115 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_114 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_43 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_113 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_112 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_111 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => n1, 
                           PGout(1) => P_32_25_port, PGout(0) => G_32_25_port);
   gblock2_4_3 : G_block_42 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_41 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => n10);
   pgblock2_4_28_2 : PG_block_110 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_109 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => n4, 
                           PGout(1) => P_32_17_port, PGout(0) => G_32_17_port);
   gblock2_5_5 : G_block_40 port map( A(1) => P_20_17_port, A(0) => n3, B => 
                           n10, Gout => Co_5_port);
   gblock2_5_6 : G_block_39 port map( A(1) => P_24_17_port, A(0) => n4, B => 
                           n10, Gout => Co_6_port);
   gblock2_5_7 : G_block_38 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => n10, Gout => Co_7_port);
   gblock2_5_8 : G_block_37 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : BUF_X1 port map( A => G_24_17_port, Z => n4);
   U2 : CLKBUF_X1 port map( A => n10, Z => Co_4_port);
   U3 : CLKBUF_X1 port map( A => G_28_25_port, Z => n1);
   U4 : CLKBUF_X1 port map( A => G_20_17_port, Z => n3);
   U5 : INV_X1 port map( A => B(0), ZN => n7);
   U6 : INV_X1 port map( A => Cin, ZN => n6);
   U7 : OAI21_X1 port map( B1 => Cin, B2 => B(0), A => A(0), ZN => n5);
   U8 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n5, ZN => n8);
   U9 : AND2_X1 port map( A1 => n9, A2 => n8, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_28
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_29
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_30
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_31
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_82
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_83
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_32
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_33
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_84
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_85
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_86
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_34
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_87
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_88
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_89
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_90
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_91
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_92
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_93
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_35
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_94
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_95
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_96
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_97
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_98
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_99
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_100
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_101
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_102
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_103
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_104
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_105
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_106
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_107
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_108
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_36
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, n12, Co_3_port, n13, n14,
      G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, G_16_9_port, 
      G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, G_12_12_port, 
      G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, G_10_9_port, 
      G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, G_6_6_port, 
      G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, G_2_2_port, 
      G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, G_32_25_port, 
      G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, G_29_29_port, 
      G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, G_27_27_port, 
      G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, G_24_23_port, 
      G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, G_22_21_port, 
      G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, G_19_19_port, 
      G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, P_32_32_port, P_32_31_port, P_32_29_port, 
      P_32_25_port, P_32_17_port, P_31_31_port, P_30_30_port, P_30_29_port, 
      P_29_29_port, P_28_28_port, P_28_27_port, P_28_25_port, P_28_17_port, 
      P_27_27_port, P_26_26_port, P_26_25_port, P_25_25_port, P_24_24_port, 
      P_24_23_port, P_24_21_port, P_24_17_port, P_23_23_port, P_22_22_port, 
      P_22_21_port, P_21_21_port, P_20_20_port, P_20_19_port, P_20_17_port, 
      P_19_19_port, P_18_18_port, P_18_17_port, P_17_17_port, n1, n2, n3, 
      Co_2_port, Co_4_port, n6, Co_1_port, n8, n9, n10, n11, n_1157 : std_logic
      ;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_4 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => n1, Pout(31) => P_32_32_port, Pout(30)
                           => P_31_31_port, Pout(29) => P_30_30_port, Pout(28) 
                           => P_29_29_port, Pout(27) => P_28_28_port, Pout(26) 
                           => P_27_27_port, Pout(25) => P_26_26_port, Pout(24) 
                           => P_25_25_port, Pout(23) => P_24_24_port, Pout(22) 
                           => P_23_23_port, Pout(21) => P_22_22_port, Pout(20) 
                           => P_21_21_port, Pout(19) => P_20_20_port, Pout(18) 
                           => P_19_19_port, Pout(17) => P_18_18_port, Pout(16) 
                           => P_17_17_port, Pout(15) => P_16_16_port, Pout(14) 
                           => P_15_15_port, Pout(13) => P_14_14_port, Pout(12) 
                           => P_13_13_port, Pout(11) => P_12_12_port, Pout(10) 
                           => P_11_11_port, Pout(9) => P_10_10_port, Pout(8) =>
                           P_9_9_port, Pout(7) => P_8_8_port, Pout(6) => 
                           P_7_7_port, Pout(5) => P_6_6_port, Pout(4) => 
                           P_5_5_port, Pout(3) => P_4_4_port, Pout(2) => 
                           P_3_3_port, Pout(1) => P_2_2_port, Pout(0) => n_1157
                           , Gout(31) => G_32_32_port, Gout(30) => G_31_31_port
                           , Gout(29) => G_30_30_port, Gout(28) => G_29_29_port
                           , Gout(27) => G_28_28_port, Gout(26) => G_27_27_port
                           , Gout(25) => G_26_26_port, Gout(24) => G_25_25_port
                           , Gout(23) => G_24_24_port, Gout(22) => G_23_23_port
                           , Gout(21) => G_22_22_port, Gout(20) => G_21_21_port
                           , Gout(19) => G_20_20_port, Gout(18) => G_19_19_port
                           , Gout(17) => G_18_18_port, Gout(16) => G_17_17_port
                           , Gout(15) => G_16_16_port, Gout(14) => G_15_15_port
                           , Gout(13) => G_14_14_port, Gout(12) => G_13_13_port
                           , Gout(11) => G_12_12_port, Gout(10) => G_11_11_port
                           , Gout(9) => G_10_10_port, Gout(8) => G_9_9_port, 
                           Gout(7) => G_8_8_port, Gout(6) => G_7_7_port, 
                           Gout(5) => G_6_6_port, Gout(4) => G_5_5_port, 
                           Gout(3) => G_4_4_port, Gout(2) => G_3_3_port, 
                           Gout(1) => G_2_2_port, Gout(0) => n11);
   gblock1_1_1 : G_block_36 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_108 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_107 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_106 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_105 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_104 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_103 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_102 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_101 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_100 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_99 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_98 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_97 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_96 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_95 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_94 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_35 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => n14);
   pgblock1_2_2 : PG_block_93 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_92 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_91 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_90 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_89 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_88 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_87 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_34 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => n14, Gout => n13);
   pgblock1_3_2 : PG_block_86 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_85 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_84 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_33 port map( A(1) => P_12_9_port, A(0) => n2, B => n13
                           , Gout => Co_3_port);
   gblock2_4_4 : G_block_32 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => n13, Gout => n12);
   pgblock2_4_28_2 : PG_block_83 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_82 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_31 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => n12, Gout => Co_5_port);
   gblock2_5_6 : G_block_30 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => n6, Gout => Co_6_port);
   gblock2_5_7 : G_block_29 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_28 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : BUF_X1 port map( A => n13, Z => Co_2_port);
   U2 : BUF_X2 port map( A => n12, Z => Co_4_port);
   U3 : CLKBUF_X1 port map( A => B(0), Z => n1);
   U4 : CLKBUF_X1 port map( A => G_12_9_port, Z => n2);
   U5 : INV_X1 port map( A => B(0), ZN => n3);
   U6 : CLKBUF_X1 port map( A => n12, Z => n6);
   U7 : CLKBUF_X1 port map( A => n14, Z => Co_1_port);
   U8 : INV_X1 port map( A => Cin, ZN => n9);
   U9 : INV_X1 port map( A => A(0), ZN => n8);
   U10 : OAI222_X1 port map( A1 => n9, A2 => n3, B1 => n8, B2 => n9, C1 => n3, 
                           C2 => n8, ZN => n10);
   U11 : AND2_X1 port map( A1 => n11, A2 => n10, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_19
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_20
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_21
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_22
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_55
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_56
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_23
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_24
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_57
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_58
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_59
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_25
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_60
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_61
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_62
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_63
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_64
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_65
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_66
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_26
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_67
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_68
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_69
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_70
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_71
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_72
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_73
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_74
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_75
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_76
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_77
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_78
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_79
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_80
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_81
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_27
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n1, n2, n3, n4, n5, n6, n7, n8, n_1158 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_3 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1158, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n8);
   gblock1_1_1 : G_block_27 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_81 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_80 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_79 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_78 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_77 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_76 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_75 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_74 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_73 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_72 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_71 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_70 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_69 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_68 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_67 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_26 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_66 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_65 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_64 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_63 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_62 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_61 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_60 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_25 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_59 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_58 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_57 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_24 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_23 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_56 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_55 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => n1, 
                           PGout(1) => P_32_17_port, PGout(0) => G_32_17_port);
   gblock2_5_5 : G_block_22 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_21 port map( A(1) => P_24_17_port, A(0) => n3, B => 
                           Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_20 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_19 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => n2, Gout => Co_8_port);
   U1 : CLKBUF_X1 port map( A => n3, Z => n1);
   U2 : CLKBUF_X1 port map( A => Co_4_port, Z => n2);
   U3 : BUF_X1 port map( A => G_24_17_port, Z => n3);
   U4 : INV_X1 port map( A => B(0), ZN => n6);
   U5 : INV_X1 port map( A => Cin, ZN => n5);
   U6 : OAI21_X1 port map( B1 => Cin, B2 => B(0), A => A(0), ZN => n4);
   U7 : OAI21_X1 port map( B1 => n6, B2 => n5, A => n4, ZN => n7);
   U8 : AND2_X1 port map( A1 => n8, A2 => n7, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_10
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_11
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_12
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_13
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_28
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_29
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_14
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_15
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_30
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_31
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_32
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_16
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_33
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_34
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_35
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_36
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_37
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_38
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_39
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_17
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_40
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_41
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_42
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_43
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_44
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_45
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_46
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_47
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_48
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_49
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_50
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_51
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_52
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_53
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_54
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_18
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n1, n2, n3, n4, n5, n_1159 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_2 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1159, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_18 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_54 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_53 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_52 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_51 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_50 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_49 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_48 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_47 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_46 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_45 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_44 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_43 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_42 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_41 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_40 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_17 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_39 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_38 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_37 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_36 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_35 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_34 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_33 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_16 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_32 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_31 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_30 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_15 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_14 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_29 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_28 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_13 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_12 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_11 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_10 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : INV_X1 port map( A => B(0), ZN => n3);
   U2 : INV_X1 port map( A => Cin, ZN => n2);
   U3 : INV_X1 port map( A => A(0), ZN => n1);
   U4 : OAI222_X1 port map( A1 => n3, A2 => n2, B1 => n1, B2 => n2, C1 => n3, 
                           C2 => n1, ZN => n4);
   U5 : AND2_X1 port map( A1 => n5, A2 => n4, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_1
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_2
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_3
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_4
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_1
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_2
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_5
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_6
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_3
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_4
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_5
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_7
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_6
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_7
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_8
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_9
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_10
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_11
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_12
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_8
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_13
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_14
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_15
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_16
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_17
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_18
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_19
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_20
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_21
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_22
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_23
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_24
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_25
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_26
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_27
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_9
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n1, n2, n3, n4, n5, n_1160 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_1 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1160, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_9 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B 
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_27 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_26 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_25 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_24 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_23 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_22 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_21 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_20 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_19 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_18 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_17 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_16 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_15 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_14 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_13 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_8 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B 
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_12 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_11 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_10 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_9 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_8 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_7 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_6 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_7 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B 
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_5 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_4 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_3 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_6 port map( A(1) => P_12_9_port, A(0) => G_12_9_port, 
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_5 port map( A(1) => P_16_9_port, A(0) => G_16_9_port, 
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_2 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_1 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_4 port map( A(1) => P_20_17_port, A(0) => G_20_17_port
                           , B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_3 port map( A(1) => P_24_17_port, A(0) => G_24_17_port
                           , B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_2 port map( A(1) => P_28_17_port, A(0) => G_28_17_port
                           , B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_1 port map( A(1) => P_32_17_port, A(0) => G_32_17_port
                           , B => Co_4_port, Gout => Co_8_port);
   U1 : INV_X1 port map( A => B(0), ZN => n3);
   U2 : INV_X1 port map( A => Cin, ZN => n2);
   U3 : OAI21_X1 port map( B1 => Cin, B2 => B(0), A => A(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => n4);
   U5 : AND2_X1 port map( A1 => n5, A2 => n4, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_7 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_7;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_6 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_6;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal C_internal, B_in_30_port, B_in_29_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46 : std_logic;

begin
   
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => n40, 
                           B(30) => B_in_30_port, B(29) => B_in_29_port, B(28) 
                           => n39, B(27) => n35, B(26) => n38, B(25) => n37, 
                           B(24) => n36, B(23) => n27, B(22) => n33, B(21) => 
                           n30, B(20) => n28, B(19) => n29, B(18) => n34, B(17)
                           => n32, B(16) => n31, B(15) => n17, B(14) => n23, 
                           B(13) => n21, B(12) => n26, B(11) => n20, B(10) => 
                           n25, B(9) => n22, B(8) => n24, B(7) => n15, B(6) => 
                           n19, B(5) => n16, B(4) => n18, B(3) => n12, B(2) => 
                           n13, B(1) => n14, B(0) => n11, Cin => C_internal, 
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => n1, B(31) => n40, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => n39, 
                           B(27) => n35, B(26) => n38, B(25) => n37, B(24) => 
                           n36, B(23) => n27, B(22) => n33, B(21) => n30, B(20)
                           => n28, B(19) => n29, B(18) => n34, B(17) => n32, 
                           B(16) => n31, B(15) => n9, B(14) => n23, B(13) => n6
                           , B(12) => n26, B(11) => n8, B(10) => n25, B(9) => 
                           n5, B(8) => n24, B(7) => n7, B(6) => n19, B(5) => n4
                           , B(4) => n18, B(3) => n2, B(2) => n13, B(1) => n14,
                           B(0) => n10, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : XNOR2_X2 port map( A => n41, B => B(1), ZN => n14);
   U5 : CLKBUF_X1 port map( A => n11, Z => n10);
   U6 : CLKBUF_X1 port map( A => A(0), Z => n1);
   U7 : CLKBUF_X1 port map( A => n12, Z => n2);
   U8 : XNOR2_X1 port map( A => n41, B => B(3), ZN => n12);
   U9 : INV_X1 port map( A => n16, ZN => n3);
   U10 : INV_X1 port map( A => n3, ZN => n4);
   U11 : XNOR2_X1 port map( A => n41, B => B(5), ZN => n16);
   U12 : BUF_X1 port map( A => n22, Z => n5);
   U13 : XNOR2_X1 port map( A => n41, B => B(9), ZN => n22);
   U14 : CLKBUF_X1 port map( A => n21, Z => n6);
   U15 : XNOR2_X1 port map( A => n42, B => B(13), ZN => n21);
   U16 : CLKBUF_X1 port map( A => n15, Z => n7);
   U17 : XNOR2_X1 port map( A => n41, B => B(7), ZN => n15);
   U18 : CLKBUF_X1 port map( A => n20, Z => n8);
   U19 : XNOR2_X1 port map( A => n41, B => B(11), ZN => n20);
   U20 : CLKBUF_X1 port map( A => n17, Z => n9);
   U21 : XNOR2_X1 port map( A => B(15), B => n42, ZN => n17);
   U22 : XNOR2_X2 port map( A => n42, B => B(20), ZN => n28);
   U23 : XNOR2_X1 port map( A => B(0), B => n41, ZN => n11);
   U24 : BUF_X1 port map( A => n46, Z => n41);
   U25 : BUF_X1 port map( A => n46, Z => n42);
   U26 : BUF_X1 port map( A => n46, Z => n43);
   U27 : XNOR2_X2 port map( A => n41, B => B(2), ZN => n13);
   U28 : XNOR2_X2 port map( A => n41, B => B(4), ZN => n18);
   U29 : XNOR2_X2 port map( A => n41, B => B(6), ZN => n19);
   U30 : XNOR2_X2 port map( A => n42, B => B(14), ZN => n23);
   U31 : XNOR2_X2 port map( A => n41, B => B(8), ZN => n24);
   U32 : XNOR2_X2 port map( A => n41, B => B(10), ZN => n25);
   U33 : XNOR2_X2 port map( A => n42, B => B(12), ZN => n26);
   U34 : XNOR2_X2 port map( A => n42, B => B(23), ZN => n27);
   U35 : XNOR2_X2 port map( A => n42, B => B(19), ZN => n29);
   U36 : XNOR2_X2 port map( A => n42, B => B(21), ZN => n30);
   U37 : XNOR2_X2 port map( A => n42, B => B(16), ZN => n31);
   U38 : XNOR2_X2 port map( A => n42, B => B(17), ZN => n32);
   U39 : XNOR2_X2 port map( A => n42, B => B(22), ZN => n33);
   U40 : XNOR2_X2 port map( A => n42, B => B(18), ZN => n34);
   U41 : XNOR2_X1 port map( A => n43, B => B(27), ZN => n35);
   U42 : XNOR2_X1 port map( A => n43, B => B(24), ZN => n36);
   U43 : XNOR2_X1 port map( A => n43, B => B(25), ZN => n37);
   U44 : XNOR2_X1 port map( A => n43, B => B(26), ZN => n38);
   U45 : XNOR2_X1 port map( A => n43, B => B(28), ZN => n39);
   U46 : XNOR2_X1 port map( A => n43, B => B(31), ZN => n40);
   U47 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U48 : INV_X1 port map( A => ADD_SUB, ZN => n46);
   U49 : XOR2_X1 port map( A => n43, B => B(29), Z => n44);
   U50 : INV_X1 port map( A => n44, ZN => B_in_29_port);
   U51 : XOR2_X1 port map( A => n43, B => B(30), Z => n45);
   U52 : INV_X1 port map( A => n45, ZN => B_in_30_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_5 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_5;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53 : std_logic;

begin
   
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => n4, A(27) 
                           => A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => n49, B(28) => n48, B(27) 
                           => n44, B(26) => n46, B(25) => n45, B(24) => n47, 
                           B(23) => n33, B(22) => n40, B(21) => n37, B(20) => 
                           n42, B(19) => n36, B(18) => n41, B(17) => n39, B(16)
                           => n43, B(15) => n26, B(14) => n32, B(13) => n30, 
                           B(12) => n38, B(11) => n29, B(10) => n35, B(9) => 
                           n31, B(8) => n34, B(7) => n23, B(6) => n28, B(5) => 
                           n24, B(4) => n27, B(3) => n21, B(2) => n25, B(1) => 
                           n22, B(0) => n20, Cin => C_internal, Co(8) => Cout, 
                           Co(7) => carry_7_port, Co(6) => carry_6_port, Co(5) 
                           => carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => n17,
                           A(26) => n9, A(25) => n18, A(24) => A(24), A(23) => 
                           n19, A(22) => n11, A(21) => n15, A(20) => A(20), 
                           A(19) => n13, A(18) => A(18), A(17) => n7, A(16) => 
                           A(16), A(15) => n14, A(14) => n3, A(13) => n5, A(12)
                           => A(12), A(11) => A(11), A(10) => A(10), A(9) => 
                           A(9), A(8) => A(8), A(7) => n2, A(6) => A(6), A(5) 
                           => A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), 
                           A(1) => A(1), A(0) => A(0), B(31) => B_in_31_port, 
                           B(30) => B_in_30_port, B(29) => n49, B(28) => n48, 
                           B(27) => n44, B(26) => n46, B(25) => n45, B(24) => 
                           n47, B(23) => n33, B(22) => n40, B(21) => n37, B(20)
                           => n42, B(19) => n36, B(18) => n41, B(17) => n39, 
                           B(16) => n43, B(15) => n26, B(14) => n32, B(13) => 
                           n30, B(12) => n38, B(11) => n29, B(10) => n35, B(9) 
                           => n31, B(8) => n34, B(7) => n23, B(6) => n28, B(5) 
                           => n24, B(4) => n27, B(3) => n21, B(2) => n25, B(1) 
                           => n22, B(0) => n20, Ci(7) => carry_7_port, Ci(6) =>
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : XNOR2_X2 port map( A => n51, B => B(15), ZN => n26);
   U5 : INV_X1 port map( A => A(7), ZN => n1);
   U6 : INV_X1 port map( A => n1, ZN => n2);
   U7 : BUF_X1 port map( A => A(14), Z => n3);
   U8 : INV_X1 port map( A => n6, ZN => n44);
   U9 : CLKBUF_X1 port map( A => A(15), Z => n14);
   U10 : CLKBUF_X1 port map( A => A(28), Z => n4);
   U11 : XNOR2_X2 port map( A => n51, B => B(19), ZN => n36);
   U14 : BUF_X2 port map( A => A(13), Z => n5);
   U15 : XNOR2_X1 port map( A => ADD_SUB, B => B(27), ZN => n6);
   U16 : XNOR2_X2 port map( A => n52, B => B(25), ZN => n45);
   U17 : XNOR2_X2 port map( A => n51, B => B(13), ZN => n30);
   U18 : CLKBUF_X1 port map( A => A(21), Z => n15);
   U19 : BUF_X2 port map( A => A(17), Z => n7);
   U20 : INV_X1 port map( A => A(26), ZN => n8);
   U21 : INV_X1 port map( A => n8, ZN => n9);
   U22 : INV_X1 port map( A => A(22), ZN => n10);
   U23 : INV_X1 port map( A => n10, ZN => n11);
   U24 : INV_X1 port map( A => A(19), ZN => n12);
   U25 : INV_X1 port map( A => n12, ZN => n13);
   U26 : CLKBUF_X1 port map( A => A(23), Z => n19);
   U27 : INV_X1 port map( A => A(27), ZN => n16);
   U28 : INV_X1 port map( A => n16, ZN => n17);
   U29 : BUF_X2 port map( A => A(25), Z => n18);
   U30 : XNOR2_X2 port map( A => n51, B => B(21), ZN => n37);
   U31 : BUF_X1 port map( A => n53, Z => n50);
   U32 : BUF_X1 port map( A => n53, Z => n51);
   U33 : BUF_X1 port map( A => n53, Z => n52);
   U34 : XNOR2_X1 port map( A => n50, B => B(0), ZN => n20);
   U35 : XNOR2_X1 port map( A => n50, B => B(3), ZN => n21);
   U36 : XNOR2_X1 port map( A => n50, B => B(1), ZN => n22);
   U37 : XNOR2_X1 port map( A => n50, B => B(7), ZN => n23);
   U38 : XNOR2_X1 port map( A => n50, B => B(5), ZN => n24);
   U39 : XNOR2_X1 port map( A => n50, B => B(2), ZN => n25);
   U40 : XNOR2_X1 port map( A => n50, B => B(4), ZN => n27);
   U41 : XNOR2_X1 port map( A => n50, B => B(6), ZN => n28);
   U42 : XNOR2_X1 port map( A => n50, B => B(11), ZN => n29);
   U43 : XNOR2_X1 port map( A => n50, B => B(9), ZN => n31);
   U44 : XNOR2_X1 port map( A => n51, B => B(14), ZN => n32);
   U45 : XNOR2_X2 port map( A => n51, B => B(23), ZN => n33);
   U46 : XNOR2_X1 port map( A => n50, B => B(8), ZN => n34);
   U47 : XNOR2_X1 port map( A => n50, B => B(10), ZN => n35);
   U48 : XNOR2_X1 port map( A => n51, B => B(12), ZN => n38);
   U49 : XNOR2_X1 port map( A => n51, B => B(17), ZN => n39);
   U50 : XNOR2_X1 port map( A => n51, B => B(22), ZN => n40);
   U51 : XNOR2_X1 port map( A => n51, B => B(18), ZN => n41);
   U52 : XNOR2_X1 port map( A => n51, B => B(20), ZN => n42);
   U53 : XNOR2_X1 port map( A => n51, B => B(16), ZN => n43);
   U54 : XNOR2_X1 port map( A => n52, B => B(26), ZN => n46);
   U55 : XNOR2_X1 port map( A => n52, B => B(24), ZN => n47);
   U56 : XNOR2_X1 port map( A => n52, B => B(28), ZN => n48);
   U57 : XNOR2_X1 port map( A => n52, B => B(29), ZN => n49);
   U58 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U59 : INV_X1 port map( A => ADD_SUB, ZN => n53);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_4 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_4;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal C_internal, B_in_30_port, B_in_29_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49 : std_logic;

begin
   
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => n43, 
                           B(30) => B_in_30_port, B(29) => B_in_29_port, B(28) 
                           => n42, B(27) => n38, B(26) => n41, B(25) => n40, 
                           B(24) => n39, B(23) => n30, B(22) => n36, B(21) => 
                           n33, B(20) => n31, B(19) => n32, B(18) => n37, B(17)
                           => n35, B(16) => n34, B(15) => n20, B(14) => n26, 
                           B(13) => n24, B(12) => n29, B(11) => n23, B(10) => 
                           n28, B(9) => n25, B(8) => n27, B(7) => n18, B(6) => 
                           n22, B(5) => n19, B(4) => n21, B(3) => n15, B(2) => 
                           n16, B(1) => n17, B(0) => n14, Cin => C_internal, 
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => n6, B(31) => n43, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => n42, 
                           B(27) => n38, B(26) => n41, B(25) => n40, B(24) => 
                           n39, B(23) => n30, B(22) => n36, B(21) => n33, B(20)
                           => n31, B(19) => n32, B(18) => n37, B(17) => n35, 
                           B(16) => n34, B(15) => n11, B(14) => n26, B(13) => 
                           n9, B(12) => n29, B(11) => n10, B(10) => n28, B(9) 
                           => n5, B(8) => n27, B(7) => n12, B(6) => n4, B(5) =>
                           n8, B(4) => n21, B(3) => n2, B(2) => n16, B(1) => n1
                           , B(0) => n13, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : XNOR2_X1 port map( A => n44, B => B(1), ZN => n1);
   U5 : XNOR2_X1 port map( A => n44, B => B(1), ZN => n17);
   U6 : XNOR2_X1 port map( A => n44, B => B(3), ZN => n2);
   U7 : XNOR2_X1 port map( A => n44, B => B(3), ZN => n15);
   U8 : CLKBUF_X1 port map( A => B(7), Z => n3);
   U9 : XNOR2_X1 port map( A => n44, B => B(6), ZN => n4);
   U10 : XNOR2_X1 port map( A => n44, B => B(6), ZN => n22);
   U11 : BUF_X1 port map( A => n25, Z => n5);
   U12 : XNOR2_X1 port map( A => n44, B => B(9), ZN => n25);
   U13 : BUF_X1 port map( A => A(0), Z => n6);
   U14 : INV_X1 port map( A => n19, ZN => n7);
   U15 : INV_X1 port map( A => n7, ZN => n8);
   U16 : XNOR2_X1 port map( A => n44, B => B(5), ZN => n19);
   U17 : CLKBUF_X1 port map( A => n24, Z => n9);
   U18 : XNOR2_X1 port map( A => n45, B => B(13), ZN => n24);
   U19 : XNOR2_X1 port map( A => B(11), B => n44, ZN => n10);
   U20 : XNOR2_X1 port map( A => B(11), B => n44, ZN => n23);
   U21 : XNOR2_X1 port map( A => B(15), B => n45, ZN => n11);
   U22 : XNOR2_X1 port map( A => B(15), B => n45, ZN => n20);
   U23 : XNOR2_X1 port map( A => n3, B => n44, ZN => n12);
   U24 : XNOR2_X1 port map( A => B(7), B => n44, ZN => n18);
   U25 : XNOR2_X2 port map( A => n45, B => B(20), ZN => n31);
   U26 : CLKBUF_X1 port map( A => n14, Z => n13);
   U27 : XNOR2_X1 port map( A => B(0), B => n44, ZN => n14);
   U28 : BUF_X1 port map( A => n49, Z => n44);
   U29 : BUF_X1 port map( A => n49, Z => n45);
   U30 : BUF_X1 port map( A => n49, Z => n46);
   U31 : XNOR2_X2 port map( A => n44, B => B(2), ZN => n16);
   U32 : XNOR2_X2 port map( A => n44, B => B(4), ZN => n21);
   U33 : XNOR2_X2 port map( A => n45, B => B(14), ZN => n26);
   U34 : XNOR2_X2 port map( A => n44, B => B(8), ZN => n27);
   U35 : XNOR2_X2 port map( A => n44, B => B(10), ZN => n28);
   U36 : XNOR2_X2 port map( A => n45, B => B(12), ZN => n29);
   U37 : XNOR2_X2 port map( A => n45, B => B(23), ZN => n30);
   U38 : XNOR2_X2 port map( A => n45, B => B(19), ZN => n32);
   U39 : XNOR2_X2 port map( A => n45, B => B(21), ZN => n33);
   U40 : XNOR2_X2 port map( A => n45, B => B(16), ZN => n34);
   U41 : XNOR2_X2 port map( A => n45, B => B(17), ZN => n35);
   U42 : XNOR2_X2 port map( A => n45, B => B(22), ZN => n36);
   U43 : XNOR2_X2 port map( A => n45, B => B(18), ZN => n37);
   U44 : XNOR2_X1 port map( A => n46, B => B(27), ZN => n38);
   U45 : XNOR2_X1 port map( A => n46, B => B(24), ZN => n39);
   U46 : XNOR2_X1 port map( A => n46, B => B(25), ZN => n40);
   U47 : XNOR2_X1 port map( A => n46, B => B(26), ZN => n41);
   U48 : XNOR2_X1 port map( A => n46, B => B(28), ZN => n42);
   U49 : XNOR2_X1 port map( A => n46, B => B(31), ZN => n43);
   U50 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U51 : INV_X1 port map( A => ADD_SUB, ZN => n49);
   U52 : XOR2_X1 port map( A => n46, B => B(29), Z => n47);
   U53 : INV_X1 port map( A => n47, ZN => B_in_29_port);
   U54 : XOR2_X1 port map( A => n46, B => B(30), Z => n48);
   U55 : INV_X1 port map( A => n48, ZN => B_in_30_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54 : std_logic;

begin
   
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => n50, 
                           B(28) => n49, B(27) => n45, B(26) => n47, B(25) => 
                           n46, B(24) => n48, B(23) => n34, B(22) => n41, B(21)
                           => n38, B(20) => n43, B(19) => n37, B(18) => n42, 
                           B(17) => n40, B(16) => n44, B(15) => n27, B(14) => 
                           n33, B(13) => n31, B(12) => n39, B(11) => n30, B(10)
                           => n36, B(9) => n32, B(8) => n35, B(7) => n24, B(6) 
                           => n29, B(5) => n25, B(4) => n28, B(3) => n22, B(2) 
                           => n26, B(1) => n23, B(0) => n21, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => n19,
                           A(26) => n2, A(25) => n13, A(24) => A(24), A(23) => 
                           n20, A(22) => n11, A(21) => n16, A(20) => n3, A(19) 
                           => n18, A(18) => A(18), A(17) => n7, A(16) => A(16),
                           A(15) => n14, A(14) => A(14), A(13) => n9, A(12) => 
                           A(12), A(11) => n5, A(10) => A(10), A(9) => A(9), 
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => n50, B(28) => n49, B(27) 
                           => n45, B(26) => n47, B(25) => n46, B(24) => n48, 
                           B(23) => n34, B(22) => n41, B(21) => n38, B(20) => 
                           n43, B(19) => n37, B(18) => n42, B(17) => n40, B(16)
                           => n44, B(15) => n27, B(14) => n33, B(13) => n31, 
                           B(12) => n39, B(11) => n30, B(10) => n36, B(9) => 
                           n32, B(8) => n35, B(7) => n24, B(6) => n29, B(5) => 
                           n25, B(4) => n28, B(3) => n22, B(2) => n26, B(1) => 
                           n23, B(0) => n21, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : BUF_X1 port map( A => A(15), Z => n14);
   U5 : XNOR2_X2 port map( A => n52, B => B(19), ZN => n37);
   U6 : CLKBUF_X1 port map( A => A(23), Z => n20);
   U7 : XNOR2_X2 port map( A => n51, B => B(9), ZN => n32);
   U8 : INV_X1 port map( A => A(26), ZN => n1);
   U9 : INV_X1 port map( A => n1, ZN => n2);
   U10 : XNOR2_X2 port map( A => n52, B => B(21), ZN => n38);
   U11 : XNOR2_X2 port map( A => n53, B => B(27), ZN => n45);
   U14 : BUF_X2 port map( A => A(20), Z => n3);
   U15 : INV_X1 port map( A => A(11), ZN => n4);
   U16 : INV_X1 port map( A => n4, ZN => n5);
   U17 : INV_X1 port map( A => A(17), ZN => n6);
   U18 : INV_X1 port map( A => n6, ZN => n7);
   U19 : INV_X1 port map( A => A(13), ZN => n8);
   U20 : INV_X1 port map( A => n8, ZN => n9);
   U21 : INV_X1 port map( A => A(22), ZN => n10);
   U22 : INV_X1 port map( A => n10, ZN => n11);
   U23 : INV_X1 port map( A => A(25), ZN => n12);
   U24 : INV_X1 port map( A => n12, ZN => n13);
   U25 : INV_X1 port map( A => A(21), ZN => n15);
   U26 : INV_X1 port map( A => n15, ZN => n16);
   U27 : INV_X1 port map( A => A(19), ZN => n17);
   U28 : INV_X1 port map( A => n17, ZN => n18);
   U29 : BUF_X2 port map( A => A(27), Z => n19);
   U30 : BUF_X1 port map( A => n54, Z => n51);
   U31 : BUF_X1 port map( A => n54, Z => n52);
   U32 : BUF_X1 port map( A => n54, Z => n53);
   U33 : XNOR2_X1 port map( A => n51, B => B(0), ZN => n21);
   U34 : XNOR2_X1 port map( A => n51, B => B(3), ZN => n22);
   U35 : XNOR2_X1 port map( A => n51, B => B(1), ZN => n23);
   U36 : XNOR2_X1 port map( A => n51, B => B(7), ZN => n24);
   U37 : XNOR2_X1 port map( A => n51, B => B(5), ZN => n25);
   U38 : XNOR2_X1 port map( A => n51, B => B(2), ZN => n26);
   U39 : XNOR2_X1 port map( A => n52, B => B(15), ZN => n27);
   U40 : XNOR2_X1 port map( A => n51, B => B(4), ZN => n28);
   U41 : XNOR2_X1 port map( A => n51, B => B(6), ZN => n29);
   U42 : XNOR2_X1 port map( A => n51, B => B(11), ZN => n30);
   U43 : XNOR2_X1 port map( A => n52, B => B(13), ZN => n31);
   U44 : XNOR2_X1 port map( A => n52, B => B(14), ZN => n33);
   U45 : XNOR2_X2 port map( A => n52, B => B(23), ZN => n34);
   U46 : XNOR2_X1 port map( A => n51, B => B(8), ZN => n35);
   U47 : XNOR2_X1 port map( A => n51, B => B(10), ZN => n36);
   U48 : XNOR2_X1 port map( A => n52, B => B(12), ZN => n39);
   U49 : XNOR2_X1 port map( A => n52, B => B(17), ZN => n40);
   U50 : XNOR2_X1 port map( A => n52, B => B(22), ZN => n41);
   U51 : XNOR2_X1 port map( A => n52, B => B(18), ZN => n42);
   U52 : XNOR2_X1 port map( A => n52, B => B(20), ZN => n43);
   U53 : XNOR2_X1 port map( A => n52, B => B(16), ZN => n44);
   U54 : XNOR2_X1 port map( A => n53, B => B(25), ZN => n46);
   U55 : XNOR2_X1 port map( A => n53, B => B(26), ZN => n47);
   U56 : XNOR2_X1 port map( A => n53, B => B(24), ZN => n48);
   U57 : XNOR2_X1 port map( A => n53, B => B(28), ZN => n49);
   U58 : XNOR2_X1 port map( A => n53, B => B(29), ZN => n50);
   U59 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U60 : INV_X1 port map( A => ADD_SUB, ZN => n54);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal C_internal, B_in_5_port, B_in_3_port, B_in_0_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, carry_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36 : std_logic;

begin
   
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => n29, 
                           B(30) => n2, B(29) => n1, B(28) => n28, B(27) => n24
                           , B(26) => n27, B(25) => n26, B(24) => n25, B(23) =>
                           n17, B(22) => n22, B(21) => n20, B(20) => n16, B(19)
                           => n19, B(18) => n23, B(17) => n21, B(16) => n18, 
                           B(15) => n8, B(14) => n12, B(13) => n10, B(12) => 
                           n15, B(11) => n9, B(10) => n14, B(9) => n11, B(8) =>
                           n13, B(7) => n4, B(6) => n7, B(5) => B_in_5_port, 
                           B(4) => n6, B(3) => B_in_3_port, B(2) => n3, B(1) =>
                           n5, B(0) => B_in_0_port, Cin => C_internal, Co(8) =>
                           Cout, Co(7) => carry_7_port, Co(6) => carry_6_port, 
                           Co(5) => carry_5_port, Co(4) => carry_4_port, Co(3) 
                           => carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => n29, B(30) => n2, 
                           B(29) => n1, B(28) => n28, B(27) => n24, B(26) => 
                           n27, B(25) => n26, B(24) => n25, B(23) => n17, B(22)
                           => n22, B(21) => n20, B(20) => n16, B(19) => n19, 
                           B(18) => n23, B(17) => n21, B(16) => n18, B(15) => 
                           n8, B(14) => n12, B(13) => n10, B(12) => n15, B(11) 
                           => n9, B(10) => n14, B(9) => n11, B(8) => n13, B(7) 
                           => n4, B(6) => n7, B(5) => n34, B(4) => n6, B(3) => 
                           n35, B(2) => n3, B(1) => n5, B(0) => n36, Ci(7) => 
                           carry_7_port, Ci(6) => carry_6_port, Ci(5) => 
                           carry_5_port, Ci(4) => carry_4_port, Ci(3) => 
                           carry_3_port, Ci(2) => carry_2_port, Ci(1) => 
                           carry_1_port, Ci(0) => carry_0_port, S(31) => S(31),
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U4 : XNOR2_X1 port map( A => n32, B => B(29), ZN => n1);
   U5 : XNOR2_X1 port map( A => n32, B => B(30), ZN => n2);
   U6 : BUF_X1 port map( A => n33, Z => n30);
   U7 : BUF_X1 port map( A => n33, Z => n31);
   U8 : BUF_X1 port map( A => n33, Z => n32);
   U9 : XNOR2_X1 port map( A => n30, B => B(2), ZN => n3);
   U10 : XNOR2_X1 port map( A => n30, B => B(7), ZN => n4);
   U11 : XNOR2_X1 port map( A => n30, B => B(1), ZN => n5);
   U12 : XNOR2_X1 port map( A => n30, B => B(4), ZN => n6);
   U13 : XNOR2_X1 port map( A => n30, B => B(6), ZN => n7);
   U14 : XNOR2_X1 port map( A => n31, B => B(15), ZN => n8);
   U15 : XNOR2_X1 port map( A => n30, B => B(11), ZN => n9);
   U16 : XNOR2_X1 port map( A => n30, B => B(13), ZN => n10);
   U17 : XNOR2_X1 port map( A => n30, B => B(9), ZN => n11);
   U18 : XNOR2_X1 port map( A => n30, B => B(14), ZN => n12);
   U19 : XNOR2_X1 port map( A => n30, B => B(8), ZN => n13);
   U20 : XNOR2_X1 port map( A => n30, B => B(10), ZN => n14);
   U21 : XNOR2_X1 port map( A => n30, B => B(12), ZN => n15);
   U22 : XNOR2_X1 port map( A => n31, B => B(20), ZN => n16);
   U23 : XNOR2_X1 port map( A => n31, B => B(23), ZN => n17);
   U24 : XNOR2_X1 port map( A => n31, B => B(16), ZN => n18);
   U25 : XNOR2_X1 port map( A => n31, B => B(19), ZN => n19);
   U26 : XNOR2_X1 port map( A => n31, B => B(21), ZN => n20);
   U27 : XNOR2_X1 port map( A => n31, B => B(17), ZN => n21);
   U28 : XNOR2_X1 port map( A => n31, B => B(22), ZN => n22);
   U29 : XNOR2_X1 port map( A => n31, B => B(18), ZN => n23);
   U30 : XNOR2_X1 port map( A => n32, B => B(27), ZN => n24);
   U31 : XNOR2_X1 port map( A => n31, B => B(24), ZN => n25);
   U32 : XNOR2_X1 port map( A => n31, B => B(25), ZN => n26);
   U33 : XNOR2_X1 port map( A => n31, B => B(26), ZN => n27);
   U34 : XNOR2_X1 port map( A => n32, B => B(28), ZN => n28);
   U35 : XNOR2_X1 port map( A => n32, B => B(31), ZN => n29);
   U36 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U37 : XOR2_X1 port map( A => ADD_SUB, B => B(0), Z => B_in_0_port);
   U38 : INV_X1 port map( A => ADD_SUB, ZN => n33);
   U39 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U40 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U41 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => n34);
   U42 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => n35);
   U43 : XOR2_X1 port map( A => ADD_SUB, B => B(0), Z => n36);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, carry_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35 : std_logic;

begin
   
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => n31, B(29) => n30, B(28) => 
                           n29, B(27) => n26, B(26) => n1, B(25) => n27, B(24) 
                           => n28, B(23) => n19, B(22) => n2, B(21) => n21, 
                           B(20) => n24, B(19) => n20, B(18) => n23, B(17) => 
                           n22, B(16) => n25, B(15) => n11, B(14) => n18, B(13)
                           => n14, B(12) => n17, B(11) => n13, B(10) => n16, 
                           B(9) => n12, B(8) => n15, B(7) => n7, B(6) => n10, 
                           B(5) => n6, B(4) => n9, B(3) => n4, B(2) => n8, B(1)
                           => n5, B(0) => n3, Cin => C_internal, Co(8) => Cout,
                           Co(7) => carry_7_port, Co(6) => carry_6_port, Co(5) 
                           => carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => n31, B(29) => n30, B(28) => n29, B(27) => n26, 
                           B(26) => n1, B(25) => n27, B(24) => n28, B(23) => 
                           n19, B(22) => n2, B(21) => n21, B(20) => n24, B(19) 
                           => n20, B(18) => n23, B(17) => n22, B(16) => n25, 
                           B(15) => n11, B(14) => n18, B(13) => n14, B(12) => 
                           n17, B(11) => n13, B(10) => n16, B(9) => n12, B(8) 
                           => n15, B(7) => n7, B(6) => n10, B(5) => n6, B(4) =>
                           n9, B(3) => n4, B(2) => n8, B(1) => n5, B(0) => n3, 
                           Ci(7) => carry_7_port, Ci(6) => carry_6_port, Ci(5) 
                           => carry_5_port, Ci(4) => carry_4_port, Ci(3) => 
                           carry_3_port, Ci(2) => carry_2_port, Ci(1) => 
                           carry_1_port, Ci(0) => carry_0_port, S(31) => S(31),
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U4 : XNOR2_X1 port map( A => n34, B => B(26), ZN => n1);
   U5 : XNOR2_X1 port map( A => n33, B => B(22), ZN => n2);
   U6 : BUF_X1 port map( A => n35, Z => n32);
   U7 : BUF_X1 port map( A => n35, Z => n33);
   U8 : BUF_X1 port map( A => n35, Z => n34);
   U9 : XNOR2_X1 port map( A => n32, B => B(0), ZN => n3);
   U10 : XNOR2_X1 port map( A => n32, B => B(3), ZN => n4);
   U11 : XNOR2_X1 port map( A => n32, B => B(1), ZN => n5);
   U13 : XNOR2_X1 port map( A => n32, B => B(5), ZN => n6);
   U14 : XNOR2_X1 port map( A => n32, B => B(7), ZN => n7);
   U15 : XNOR2_X1 port map( A => n32, B => B(2), ZN => n8);
   U16 : XNOR2_X1 port map( A => n32, B => B(4), ZN => n9);
   U17 : XNOR2_X1 port map( A => n32, B => B(6), ZN => n10);
   U18 : XNOR2_X1 port map( A => n33, B => B(15), ZN => n11);
   U19 : XNOR2_X1 port map( A => n32, B => B(9), ZN => n12);
   U20 : XNOR2_X1 port map( A => n32, B => B(11), ZN => n13);
   U21 : XNOR2_X1 port map( A => n33, B => B(13), ZN => n14);
   U22 : XNOR2_X1 port map( A => n32, B => B(8), ZN => n15);
   U23 : XNOR2_X1 port map( A => n32, B => B(10), ZN => n16);
   U24 : XNOR2_X1 port map( A => n33, B => B(12), ZN => n17);
   U25 : XNOR2_X1 port map( A => n33, B => B(14), ZN => n18);
   U26 : XNOR2_X1 port map( A => n33, B => B(23), ZN => n19);
   U27 : XNOR2_X1 port map( A => n33, B => B(19), ZN => n20);
   U28 : XNOR2_X1 port map( A => n33, B => B(21), ZN => n21);
   U29 : XNOR2_X1 port map( A => n33, B => B(17), ZN => n22);
   U30 : XNOR2_X1 port map( A => n33, B => B(18), ZN => n23);
   U31 : XNOR2_X1 port map( A => n33, B => B(20), ZN => n24);
   U32 : XNOR2_X1 port map( A => n33, B => B(16), ZN => n25);
   U33 : XNOR2_X1 port map( A => n34, B => B(27), ZN => n26);
   U34 : XNOR2_X1 port map( A => n34, B => B(25), ZN => n27);
   U35 : XNOR2_X1 port map( A => n34, B => B(24), ZN => n28);
   U36 : XNOR2_X1 port map( A => n34, B => B(28), ZN => n29);
   U37 : XNOR2_X1 port map( A => n34, B => B(29), ZN => n30);
   U38 : XNOR2_X1 port map( A => n34, B => B(30), ZN => n31);
   U39 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U40 : INV_X1 port map( A => ADD_SUB, ZN => n35);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_228;

architecture SYN_Behavioral of AND2_228 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_227;

architecture SYN_Behavioral of AND2_227 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_226;

architecture SYN_Behavioral of AND2_226 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_225;

architecture SYN_Behavioral of AND2_225 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_224;

architecture SYN_Behavioral of AND2_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_223;

architecture SYN_Behavioral of AND2_223 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_222;

architecture SYN_Behavioral of AND2_222 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_221;

architecture SYN_Behavioral of AND2_221 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_220;

architecture SYN_Behavioral of AND2_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_219;

architecture SYN_Behavioral of AND2_219 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_218;

architecture SYN_Behavioral of AND2_218 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_217;

architecture SYN_Behavioral of AND2_217 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_216;

architecture SYN_Behavioral of AND2_216 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_215;

architecture SYN_Behavioral of AND2_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_214;

architecture SYN_Behavioral of AND2_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_213;

architecture SYN_Behavioral of AND2_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_212;

architecture SYN_Behavioral of AND2_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_211;

architecture SYN_Behavioral of AND2_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_210;

architecture SYN_Behavioral of AND2_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_209;

architecture SYN_Behavioral of AND2_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_208;

architecture SYN_Behavioral of AND2_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_207;

architecture SYN_Behavioral of AND2_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_206;

architecture SYN_Behavioral of AND2_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_205;

architecture SYN_Behavioral of AND2_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_204;

architecture SYN_Behavioral of AND2_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_203;

architecture SYN_Behavioral of AND2_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_202;

architecture SYN_Behavioral of AND2_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_201;

architecture SYN_Behavioral of AND2_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_200;

architecture SYN_Behavioral of AND2_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_199;

architecture SYN_Behavioral of AND2_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_198;

architecture SYN_Behavioral of AND2_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_197;

architecture SYN_Behavioral of AND2_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_196;

architecture SYN_Behavioral of AND2_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_195;

architecture SYN_Behavioral of AND2_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_194;

architecture SYN_Behavioral of AND2_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_193;

architecture SYN_Behavioral of AND2_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_192;

architecture SYN_Behavioral of AND2_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_191;

architecture SYN_Behavioral of AND2_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_190;

architecture SYN_Behavioral of AND2_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_189;

architecture SYN_Behavioral of AND2_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_188;

architecture SYN_Behavioral of AND2_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_187;

architecture SYN_Behavioral of AND2_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_186;

architecture SYN_Behavioral of AND2_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_185;

architecture SYN_Behavioral of AND2_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_184;

architecture SYN_Behavioral of AND2_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_183;

architecture SYN_Behavioral of AND2_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_182;

architecture SYN_Behavioral of AND2_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_181;

architecture SYN_Behavioral of AND2_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_180;

architecture SYN_Behavioral of AND2_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_179;

architecture SYN_Behavioral of AND2_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_178;

architecture SYN_Behavioral of AND2_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_177;

architecture SYN_Behavioral of AND2_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_176;

architecture SYN_Behavioral of AND2_176 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_175;

architecture SYN_Behavioral of AND2_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_174;

architecture SYN_Behavioral of AND2_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_173;

architecture SYN_Behavioral of AND2_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_172;

architecture SYN_Behavioral of AND2_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_171;

architecture SYN_Behavioral of AND2_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_170;

architecture SYN_Behavioral of AND2_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_169;

architecture SYN_Behavioral of AND2_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_168;

architecture SYN_Behavioral of AND2_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_167;

architecture SYN_Behavioral of AND2_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_166;

architecture SYN_Behavioral of AND2_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_165;

architecture SYN_Behavioral of AND2_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_164;

architecture SYN_Behavioral of AND2_164 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_163;

architecture SYN_Behavioral of AND2_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_162;

architecture SYN_Behavioral of AND2_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_161;

architecture SYN_Behavioral of AND2_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_160;

architecture SYN_Behavioral of AND2_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_159;

architecture SYN_Behavioral of AND2_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_158;

architecture SYN_Behavioral of AND2_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_157;

architecture SYN_Behavioral of AND2_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_156;

architecture SYN_Behavioral of AND2_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_155;

architecture SYN_Behavioral of AND2_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_154;

architecture SYN_Behavioral of AND2_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_153;

architecture SYN_Behavioral of AND2_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_152;

architecture SYN_Behavioral of AND2_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_151;

architecture SYN_Behavioral of AND2_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_150;

architecture SYN_Behavioral of AND2_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_149;

architecture SYN_Behavioral of AND2_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_148;

architecture SYN_Behavioral of AND2_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_147;

architecture SYN_Behavioral of AND2_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_146;

architecture SYN_Behavioral of AND2_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_145;

architecture SYN_Behavioral of AND2_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_144;

architecture SYN_Behavioral of AND2_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_143;

architecture SYN_Behavioral of AND2_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_142;

architecture SYN_Behavioral of AND2_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_141;

architecture SYN_Behavioral of AND2_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_140;

architecture SYN_Behavioral of AND2_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_139;

architecture SYN_Behavioral of AND2_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_138;

architecture SYN_Behavioral of AND2_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_137;

architecture SYN_Behavioral of AND2_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_136;

architecture SYN_Behavioral of AND2_136 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_135;

architecture SYN_Behavioral of AND2_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_134;

architecture SYN_Behavioral of AND2_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_133;

architecture SYN_Behavioral of AND2_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_132;

architecture SYN_Behavioral of AND2_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_131;

architecture SYN_Behavioral of AND2_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_130;

architecture SYN_Behavioral of AND2_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_129;

architecture SYN_Behavioral of AND2_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_128;

architecture SYN_Behavioral of AND2_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_127;

architecture SYN_Behavioral of AND2_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_126;

architecture SYN_Behavioral of AND2_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_125;

architecture SYN_Behavioral of AND2_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_124;

architecture SYN_Behavioral of AND2_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_123;

architecture SYN_Behavioral of AND2_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_122;

architecture SYN_Behavioral of AND2_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_121;

architecture SYN_Behavioral of AND2_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_120;

architecture SYN_Behavioral of AND2_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_119;

architecture SYN_Behavioral of AND2_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_118;

architecture SYN_Behavioral of AND2_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_117;

architecture SYN_Behavioral of AND2_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_116;

architecture SYN_Behavioral of AND2_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_115;

architecture SYN_Behavioral of AND2_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_114;

architecture SYN_Behavioral of AND2_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_113;

architecture SYN_Behavioral of AND2_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_112;

architecture SYN_Behavioral of AND2_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_111;

architecture SYN_Behavioral of AND2_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_110;

architecture SYN_Behavioral of AND2_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_109;

architecture SYN_Behavioral of AND2_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_108;

architecture SYN_Behavioral of AND2_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_107;

architecture SYN_Behavioral of AND2_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_106;

architecture SYN_Behavioral of AND2_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_105;

architecture SYN_Behavioral of AND2_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_104;

architecture SYN_Behavioral of AND2_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_103;

architecture SYN_Behavioral of AND2_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_102;

architecture SYN_Behavioral of AND2_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_101;

architecture SYN_Behavioral of AND2_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_100;

architecture SYN_Behavioral of AND2_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_99;

architecture SYN_Behavioral of AND2_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_98;

architecture SYN_Behavioral of AND2_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_97;

architecture SYN_Behavioral of AND2_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_96;

architecture SYN_Behavioral of AND2_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_95;

architecture SYN_Behavioral of AND2_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_94;

architecture SYN_Behavioral of AND2_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_93;

architecture SYN_Behavioral of AND2_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_92;

architecture SYN_Behavioral of AND2_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_91;

architecture SYN_Behavioral of AND2_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_90;

architecture SYN_Behavioral of AND2_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_89;

architecture SYN_Behavioral of AND2_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_88;

architecture SYN_Behavioral of AND2_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_87;

architecture SYN_Behavioral of AND2_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_86;

architecture SYN_Behavioral of AND2_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_85;

architecture SYN_Behavioral of AND2_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_84;

architecture SYN_Behavioral of AND2_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_83;

architecture SYN_Behavioral of AND2_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_82;

architecture SYN_Behavioral of AND2_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_81;

architecture SYN_Behavioral of AND2_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_80;

architecture SYN_Behavioral of AND2_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_79;

architecture SYN_Behavioral of AND2_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_78;

architecture SYN_Behavioral of AND2_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_77;

architecture SYN_Behavioral of AND2_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_76;

architecture SYN_Behavioral of AND2_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_75;

architecture SYN_Behavioral of AND2_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_74;

architecture SYN_Behavioral of AND2_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_73;

architecture SYN_Behavioral of AND2_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_72;

architecture SYN_Behavioral of AND2_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_71;

architecture SYN_Behavioral of AND2_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_70;

architecture SYN_Behavioral of AND2_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_69;

architecture SYN_Behavioral of AND2_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_68;

architecture SYN_Behavioral of AND2_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_67;

architecture SYN_Behavioral of AND2_67 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_66;

architecture SYN_Behavioral of AND2_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_65;

architecture SYN_Behavioral of AND2_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_64;

architecture SYN_Behavioral of AND2_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_63;

architecture SYN_Behavioral of AND2_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_62;

architecture SYN_Behavioral of AND2_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_61;

architecture SYN_Behavioral of AND2_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_60;

architecture SYN_Behavioral of AND2_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_59;

architecture SYN_Behavioral of AND2_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_58;

architecture SYN_Behavioral of AND2_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_57;

architecture SYN_Behavioral of AND2_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_56;

architecture SYN_Behavioral of AND2_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_55;

architecture SYN_Behavioral of AND2_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_54;

architecture SYN_Behavioral of AND2_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_53;

architecture SYN_Behavioral of AND2_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_52;

architecture SYN_Behavioral of AND2_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_51;

architecture SYN_Behavioral of AND2_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_50;

architecture SYN_Behavioral of AND2_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_49;

architecture SYN_Behavioral of AND2_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_48;

architecture SYN_Behavioral of AND2_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_47;

architecture SYN_Behavioral of AND2_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_46;

architecture SYN_Behavioral of AND2_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_45;

architecture SYN_Behavioral of AND2_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_44;

architecture SYN_Behavioral of AND2_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_43;

architecture SYN_Behavioral of AND2_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_42;

architecture SYN_Behavioral of AND2_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_41;

architecture SYN_Behavioral of AND2_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_40;

architecture SYN_Behavioral of AND2_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_39;

architecture SYN_Behavioral of AND2_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_38;

architecture SYN_Behavioral of AND2_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_37;

architecture SYN_Behavioral of AND2_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_36;

architecture SYN_Behavioral of AND2_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_35;

architecture SYN_Behavioral of AND2_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_34;

architecture SYN_Behavioral of AND2_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_33;

architecture SYN_Behavioral of AND2_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_32;

architecture SYN_Behavioral of AND2_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_31;

architecture SYN_Behavioral of AND2_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_30;

architecture SYN_Behavioral of AND2_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_29;

architecture SYN_Behavioral of AND2_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_28;

architecture SYN_Behavioral of AND2_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_27;

architecture SYN_Behavioral of AND2_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_26;

architecture SYN_Behavioral of AND2_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_25;

architecture SYN_Behavioral of AND2_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_24;

architecture SYN_Behavioral of AND2_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_23;

architecture SYN_Behavioral of AND2_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_22;

architecture SYN_Behavioral of AND2_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_21;

architecture SYN_Behavioral of AND2_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_20;

architecture SYN_Behavioral of AND2_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_19;

architecture SYN_Behavioral of AND2_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_18;

architecture SYN_Behavioral of AND2_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_17;

architecture SYN_Behavioral of AND2_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_16;

architecture SYN_Behavioral of AND2_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_15;

architecture SYN_Behavioral of AND2_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_14;

architecture SYN_Behavioral of AND2_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_13;

architecture SYN_Behavioral of AND2_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_12;

architecture SYN_Behavioral of AND2_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_11;

architecture SYN_Behavioral of AND2_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_10;

architecture SYN_Behavioral of AND2_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_9;

architecture SYN_Behavioral of AND2_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_8;

architecture SYN_Behavioral of AND2_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_7;

architecture SYN_Behavioral of AND2_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_6;

architecture SYN_Behavioral of AND2_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_5;

architecture SYN_Behavioral of AND2_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_4;

architecture SYN_Behavioral of AND2_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_3;

architecture SYN_Behavioral of AND2_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_2;

architecture SYN_Behavioral of AND2_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_1;

architecture SYN_Behavioral of AND2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX4to1_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX4to1_NBIT32_1;

architecture SYN_Behavioral of MUX4to1_NBIT32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n3, Z => n11);
   U2 : BUF_X1 port map( A => n4, Z => n15);
   U3 : AND2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n1);
   U4 : AND2_X1 port map( A1 => SEL(0), A2 => n20, ZN => n2);
   U5 : BUF_X1 port map( A => n11, Z => n10);
   U6 : BUF_X1 port map( A => n15, Z => n14);
   U7 : BUF_X1 port map( A => n15, Z => n13);
   U8 : BUF_X1 port map( A => n11, Z => n8);
   U9 : CLKBUF_X1 port map( A => n11, Z => n9);
   U10 : CLKBUF_X1 port map( A => n15, Z => n12);
   U11 : BUF_X1 port map( A => n2, Z => n18);
   U12 : BUF_X1 port map( A => n2, Z => n16);
   U13 : BUF_X1 port map( A => n2, Z => n17);
   U14 : BUF_X1 port map( A => n1, Z => n5);
   U15 : AND2_X1 port map( A1 => n19, A2 => n20, ZN => n3);
   U16 : AND2_X1 port map( A1 => SEL(1), A2 => n19, ZN => n4);
   U17 : BUF_X1 port map( A => n1, Z => n6);
   U18 : BUF_X1 port map( A => n1, Z => n7);
   U19 : INV_X1 port map( A => SEL(0), ZN => n19);
   U20 : AOI22_X1 port map( A1 => C(0), A2 => n12, B1 => D(0), B2 => n6, ZN => 
                           n22);
   U21 : INV_X1 port map( A => SEL(1), ZN => n20);
   U22 : AOI22_X1 port map( A1 => A(0), A2 => n8, B1 => B(0), B2 => n16, ZN => 
                           n21);
   U23 : NAND2_X1 port map( A1 => n22, A2 => n21, ZN => Y(0));
   U24 : AOI22_X1 port map( A1 => C(1), A2 => n13, B1 => D(1), B2 => n6, ZN => 
                           n24);
   U25 : AOI22_X1 port map( A1 => A(1), A2 => n10, B1 => B(1), B2 => n18, ZN =>
                           n23);
   U26 : NAND2_X1 port map( A1 => n24, A2 => n23, ZN => Y(1));
   U27 : AOI22_X1 port map( A1 => C(2), A2 => n13, B1 => D(2), B2 => n7, ZN => 
                           n26);
   U28 : AOI22_X1 port map( A1 => A(2), A2 => n10, B1 => B(2), B2 => n18, ZN =>
                           n25);
   U29 : NAND2_X1 port map( A1 => n26, A2 => n25, ZN => Y(2));
   U30 : AOI22_X1 port map( A1 => C(3), A2 => n13, B1 => D(3), B2 => n7, ZN => 
                           n28);
   U31 : AOI22_X1 port map( A1 => A(3), A2 => n10, B1 => B(3), B2 => n18, ZN =>
                           n27);
   U32 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => Y(3));
   U33 : AOI22_X1 port map( A1 => C(4), A2 => n13, B1 => D(4), B2 => n7, ZN => 
                           n30);
   U34 : AOI22_X1 port map( A1 => A(4), A2 => n10, B1 => B(4), B2 => n17, ZN =>
                           n29);
   U35 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => Y(4));
   U36 : AOI22_X1 port map( A1 => C(5), A2 => n13, B1 => D(5), B2 => n7, ZN => 
                           n32);
   U37 : AOI22_X1 port map( A1 => A(5), A2 => n9, B1 => B(5), B2 => n18, ZN => 
                           n31);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => Y(5));
   U39 : AOI22_X1 port map( A1 => C(6), A2 => n13, B1 => D(6), B2 => n7, ZN => 
                           n34);
   U40 : AOI22_X1 port map( A1 => A(6), A2 => n9, B1 => B(6), B2 => n18, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y(6));
   U42 : AOI22_X1 port map( A1 => C(7), A2 => n13, B1 => D(7), B2 => n7, ZN => 
                           n36);
   U43 : AOI22_X1 port map( A1 => A(7), A2 => n9, B1 => B(7), B2 => n17, ZN => 
                           n35);
   U44 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => Y(7));
   U45 : AOI22_X1 port map( A1 => C(8), A2 => n13, B1 => D(8), B2 => n7, ZN => 
                           n38);
   U46 : AOI22_X1 port map( A1 => A(8), A2 => n9, B1 => B(8), B2 => n17, ZN => 
                           n37);
   U47 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => Y(8));
   U48 : AOI22_X1 port map( A1 => C(9), A2 => n12, B1 => D(9), B2 => n7, ZN => 
                           n40);
   U49 : AOI22_X1 port map( A1 => A(9), A2 => n9, B1 => B(9), B2 => n17, ZN => 
                           n39);
   U50 : NAND2_X1 port map( A1 => n40, A2 => n39, ZN => Y(9));
   U51 : AOI22_X1 port map( A1 => C(10), A2 => n12, B1 => D(10), B2 => n6, ZN 
                           => n42);
   U52 : AOI22_X1 port map( A1 => A(10), A2 => n9, B1 => B(10), B2 => n17, ZN 
                           => n41);
   U53 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => Y(10));
   U54 : AOI22_X1 port map( A1 => C(11), A2 => n12, B1 => D(11), B2 => n6, ZN 
                           => n44);
   U55 : AOI22_X1 port map( A1 => A(11), A2 => n9, B1 => B(11), B2 => n17, ZN 
                           => n43);
   U56 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => Y(11));
   U57 : AOI22_X1 port map( A1 => C(12), A2 => n12, B1 => D(12), B2 => n6, ZN 
                           => n46);
   U58 : AOI22_X1 port map( A1 => A(12), A2 => n9, B1 => B(12), B2 => n17, ZN 
                           => n45);
   U59 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => Y(12));
   U60 : AOI22_X1 port map( A1 => C(13), A2 => n12, B1 => D(13), B2 => n6, ZN 
                           => n48);
   U61 : AOI22_X1 port map( A1 => A(13), A2 => n9, B1 => B(13), B2 => n17, ZN 
                           => n47);
   U62 : NAND2_X1 port map( A1 => n48, A2 => n47, ZN => Y(13));
   U63 : AOI22_X1 port map( A1 => C(14), A2 => n12, B1 => D(14), B2 => n6, ZN 
                           => n50);
   U64 : AOI22_X1 port map( A1 => A(14), A2 => n9, B1 => B(14), B2 => n17, ZN 
                           => n49);
   U65 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => Y(14));
   U66 : AOI22_X1 port map( A1 => C(15), A2 => n12, B1 => D(15), B2 => n6, ZN 
                           => n52);
   U67 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => B(15), B2 => n17, ZN 
                           => n51);
   U68 : NAND2_X1 port map( A1 => n52, A2 => n51, ZN => Y(15));
   U69 : AOI22_X1 port map( A1 => C(16), A2 => n12, B1 => D(16), B2 => n6, ZN 
                           => n54);
   U70 : AOI22_X1 port map( A1 => A(16), A2 => n8, B1 => B(16), B2 => n17, ZN 
                           => n53);
   U71 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => Y(16));
   U72 : AOI22_X1 port map( A1 => C(17), A2 => n12, B1 => D(17), B2 => n6, ZN 
                           => n56);
   U73 : AOI22_X1 port map( A1 => A(17), A2 => n8, B1 => B(17), B2 => n16, ZN 
                           => n55);
   U74 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => Y(17));
   U75 : AOI22_X1 port map( A1 => C(18), A2 => n12, B1 => D(18), B2 => n6, ZN 
                           => n58);
   U76 : AOI22_X1 port map( A1 => A(18), A2 => n8, B1 => B(18), B2 => n16, ZN 
                           => n57);
   U77 : NAND2_X1 port map( A1 => n58, A2 => n57, ZN => Y(18));
   U78 : AOI22_X1 port map( A1 => C(19), A2 => n12, B1 => D(19), B2 => n6, ZN 
                           => n60);
   U79 : AOI22_X1 port map( A1 => A(19), A2 => n8, B1 => B(19), B2 => n16, ZN 
                           => n59);
   U80 : NAND2_X1 port map( A1 => n60, A2 => n59, ZN => Y(19));
   U81 : AOI222_X1 port map( A1 => A(20), A2 => n8, B1 => B(20), B2 => n18, C1 
                           => C(20), C2 => n14, ZN => n62);
   U82 : NAND2_X1 port map( A1 => D(20), A2 => n5, ZN => n61);
   U83 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => Y(20));
   U84 : AOI222_X1 port map( A1 => A(21), A2 => n8, B1 => B(21), B2 => n18, C1 
                           => C(21), C2 => n14, ZN => n64);
   U85 : NAND2_X1 port map( A1 => D(21), A2 => n5, ZN => n63);
   U86 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => Y(21));
   U87 : AOI222_X1 port map( A1 => A(22), A2 => n8, B1 => B(22), B2 => n18, C1 
                           => C(22), C2 => n14, ZN => n66);
   U88 : NAND2_X1 port map( A1 => D(22), A2 => n5, ZN => n65);
   U89 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => Y(22));
   U90 : AOI22_X1 port map( A1 => D(23), A2 => n5, B1 => C(23), B2 => n13, ZN 
                           => n68);
   U91 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => B(23), B2 => n17, ZN 
                           => n67);
   U92 : NAND2_X1 port map( A1 => n68, A2 => n67, ZN => Y(23));
   U93 : AOI22_X1 port map( A1 => D(24), A2 => n5, B1 => C(24), B2 => n13, ZN 
                           => n70);
   U94 : AOI22_X1 port map( A1 => A(24), A2 => n8, B1 => B(24), B2 => n16, ZN 
                           => n69);
   U95 : NAND2_X1 port map( A1 => n70, A2 => n69, ZN => Y(24));
   U96 : AOI22_X1 port map( A1 => D(25), A2 => n5, B1 => C(25), B2 => n13, ZN 
                           => n72);
   U97 : AOI22_X1 port map( A1 => A(25), A2 => n8, B1 => B(25), B2 => n16, ZN 
                           => n71);
   U98 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => Y(25));
   U99 : AOI22_X1 port map( A1 => D(26), A2 => n5, B1 => C(26), B2 => n13, ZN 
                           => n74);
   U100 : AOI22_X1 port map( A1 => A(26), A2 => n8, B1 => B(26), B2 => n16, ZN 
                           => n73);
   U101 : NAND2_X1 port map( A1 => n74, A2 => n73, ZN => Y(26));
   U102 : AOI22_X1 port map( A1 => D(27), A2 => n5, B1 => C(27), B2 => n14, ZN 
                           => n76);
   U103 : AOI22_X1 port map( A1 => A(27), A2 => n8, B1 => B(27), B2 => n16, ZN 
                           => n75);
   U104 : NAND2_X1 port map( A1 => n76, A2 => n75, ZN => Y(27));
   U105 : NAND2_X1 port map( A1 => D(28), A2 => n5, ZN => n78);
   U106 : AOI222_X1 port map( A1 => B(28), A2 => n16, B1 => C(28), B2 => n14, 
                           C1 => A(28), C2 => n10, ZN => n77);
   U107 : NAND2_X1 port map( A1 => n78, A2 => n77, ZN => Y(28));
   U108 : NAND2_X1 port map( A1 => D(29), A2 => n5, ZN => n80);
   U109 : AOI222_X1 port map( A1 => B(29), A2 => n16, B1 => C(29), B2 => n14, 
                           C1 => A(29), C2 => n10, ZN => n79);
   U110 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => Y(29));
   U111 : NAND2_X1 port map( A1 => D(30), A2 => n5, ZN => n82);
   U112 : AOI222_X1 port map( A1 => B(30), A2 => n16, B1 => C(30), B2 => n14, 
                           C1 => A(30), C2 => n10, ZN => n81);
   U113 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => Y(30));
   U114 : NAND2_X1 port map( A1 => D(31), A2 => n5, ZN => n84);
   U115 : AOI222_X1 port map( A1 => B(31), A2 => n16, B1 => C(31), B2 => n14, 
                           C1 => A(31), C2 => n10, ZN => n83);
   U116 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => Y(31));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_8 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_8;

architecture SYN_Behavioral of MUX5to1_NBIT32_8 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n164, Z => n90);
   U6 : BUF_X1 port map( A => n161, Z => n78);
   U7 : BUF_X1 port map( A => n160, Z => n74);
   U8 : BUF_X1 port map( A => n163, Z => n83);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : INV_X1 port map( A => SEL(1), ZN => n95);
   U15 : INV_X1 port map( A => SEL(0), ZN => n96);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n74, Z => n2);
   U19 : BUF_X1 port map( A => n74, Z => n1);
   U20 : BUF_X1 port map( A => n83, Z => n85);
   U21 : BUF_X1 port map( A => n83, Z => n84);
   U22 : BUF_X1 port map( A => n82, Z => n80);
   U23 : BUF_X1 port map( A => n82, Z => n79);
   U24 : BUF_X1 port map( A => n90, Z => n88);
   U25 : BUF_X1 port map( A => n90, Z => n87);
   U26 : BUF_X1 port map( A => n78, Z => n77);
   U27 : BUF_X1 port map( A => n74, Z => n73);
   U28 : BUF_X1 port map( A => n83, Z => n86);
   U29 : BUF_X1 port map( A => n82, Z => n81);
   U30 : BUF_X1 port map( A => n90, Z => n89);
   U31 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U32 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U34 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U35 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U36 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U37 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN =>
                           n101);
   U38 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U39 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U40 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN =>
                           n103);
   U41 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U42 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U43 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN =>
                           n105);
   U44 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U45 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U46 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN =>
                           n107);
   U47 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U48 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U49 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n109);
   U50 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U51 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U52 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n111);
   U53 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U54 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U55 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n113);
   U56 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U57 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U58 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n115);
   U59 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U60 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U61 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n117);
   U62 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U63 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U64 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U65 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n80, ZN => n118);
   U66 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U67 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U68 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n120);
   U69 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U70 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U71 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U72 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U73 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U74 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U75 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U76 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U77 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U78 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U79 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U80 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U81 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U82 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U83 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U84 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U85 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U86 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U87 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U88 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U89 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U90 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U91 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U92 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U93 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U94 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U95 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U96 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U97 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U98 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U99 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U100 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U101 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, 
                           C1 => D(22), C2 => n79, ZN => n142);
   U102 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U103 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U104 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, 
                           C1 => D(23), C2 => n79, ZN => n144);
   U105 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U106 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U107 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, 
                           C1 => D(24), C2 => n79, ZN => n146);
   U108 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U109 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U110 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n79, ZN => n148);
   U111 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U112 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U113 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n79, ZN => n150);
   U114 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U115 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U116 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n79, ZN => n152);
   U117 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U118 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U119 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n79, ZN => n154);
   U120 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U121 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U122 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n79, ZN => n156);
   U123 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U124 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U125 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n79, ZN => n158);
   U126 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U127 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U128 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n79, ZN => n165);
   U129 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U130 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n99);
   U131 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_7 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_7;

architecture SYN_Behavioral of MUX5to1_NBIT32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U37 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN =>
                           n105);
   U38 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U39 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U40 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN =>
                           n107);
   U41 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U42 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U43 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n109);
   U44 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U45 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U46 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n111);
   U47 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U48 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U49 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n113);
   U50 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U51 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U52 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n115);
   U53 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U54 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U55 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n117);
   U56 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U57 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U58 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U59 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n80, ZN => n118);
   U60 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U61 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U62 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n120);
   U63 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U64 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U65 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U66 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U67 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U68 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U69 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U70 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U71 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U72 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U73 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U74 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U75 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U76 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U77 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U78 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U79 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U80 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U81 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U82 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U83 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U84 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U85 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U86 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U87 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U88 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U89 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U90 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U91 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U92 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U93 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U94 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U95 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U96 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U97 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U98 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U99 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U100 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U101 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, 
                           C1 => D(24), C2 => n79, ZN => n146);
   U102 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U103 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U104 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n79, ZN => n148);
   U105 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U106 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U107 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n79, ZN => n150);
   U108 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U109 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U110 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n79, ZN => n152);
   U111 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U112 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U113 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n79, ZN => n154);
   U114 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U115 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U116 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n79, ZN => n156);
   U117 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U118 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U119 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n79, ZN => n158);
   U120 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U121 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U122 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n79, ZN => n165);
   U123 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U124 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n103);
   U125 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U126 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U127 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n99);
   U128 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U129 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U130 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n101);
   U131 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_6 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_6;

architecture SYN_Behavioral of MUX5to1_NBIT32_6 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U37 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n109);
   U38 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U39 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U40 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n111);
   U41 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U42 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U43 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n113);
   U44 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U45 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U46 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n115);
   U47 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U48 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U49 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n117);
   U50 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U51 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U52 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U53 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n80, ZN => n118);
   U54 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U55 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U56 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n120);
   U57 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U58 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U59 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U60 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U61 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U62 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U63 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U64 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U65 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U66 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U67 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U68 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U69 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U70 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U71 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U72 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U73 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U74 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U75 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U76 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U77 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U78 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U79 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U80 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U81 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U82 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U83 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U84 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U85 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U86 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U87 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U88 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U89 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U90 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U91 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U92 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U93 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U94 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U95 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n79, ZN => n146);
   U96 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U97 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U98 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n79, ZN => n148);
   U99 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U100 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U101 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n79, ZN => n150);
   U102 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U103 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U104 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n79, ZN => n152);
   U105 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U106 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U107 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n79, ZN => n154);
   U108 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U109 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U110 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n79, ZN => n156);
   U111 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U112 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U113 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n79, ZN => n158);
   U114 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U115 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U116 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n79, ZN => n165);
   U117 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U118 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n107);
   U119 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U120 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U121 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n99);
   U122 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U123 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U124 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n101);
   U125 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U126 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U127 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n103);
   U128 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U129 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U130 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n105);
   U131 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_5 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_5;

architecture SYN_Behavioral of MUX5to1_NBIT32_5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U37 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n113);
   U38 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U39 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U40 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n115);
   U41 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U42 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U43 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n117);
   U44 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U45 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U46 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U47 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n80, ZN => n118);
   U48 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U49 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U50 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n120);
   U51 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U52 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U53 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U54 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U55 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U56 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U57 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U58 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U59 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U60 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U61 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U62 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U63 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U64 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U65 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U66 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U67 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U68 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U69 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U70 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U71 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U72 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U73 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U74 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U75 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U76 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U77 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U78 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U79 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U80 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U81 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U82 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U83 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U84 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U85 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U86 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U87 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U88 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U89 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n79, ZN => n146);
   U90 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U91 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U92 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n79, ZN => n148);
   U93 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U94 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U95 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n79, ZN => n150);
   U96 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U97 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U98 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n79, ZN => n152);
   U99 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U100 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U101 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n79, ZN => n154);
   U102 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U103 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U104 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n79, ZN => n156);
   U105 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U106 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U107 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n79, ZN => n158);
   U108 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U109 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U110 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n79, ZN => n165);
   U111 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U112 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n111);
   U113 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U114 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U115 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n99);
   U116 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U117 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U118 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n101);
   U119 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U120 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U121 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n103);
   U122 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U123 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U124 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n105);
   U125 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U126 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U127 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n107);
   U128 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U129 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U130 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n109);
   U131 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_4 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_4;

architecture SYN_Behavioral of MUX5to1_NBIT32_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U37 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n117);
   U38 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U39 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U40 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U41 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n80, ZN => n118);
   U42 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U43 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U44 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n120);
   U45 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U46 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U47 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U48 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U49 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U50 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U51 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U52 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U53 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U54 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U55 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U56 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U57 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U58 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U59 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U60 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U61 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U62 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U63 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U64 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U65 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U66 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U67 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U68 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U69 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U70 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U71 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U72 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U73 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U74 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U75 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U76 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U77 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U78 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U79 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U80 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U81 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U82 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U83 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n79, ZN => n146);
   U84 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U85 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U86 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n79, ZN => n148);
   U87 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U88 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U89 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n79, ZN => n150);
   U90 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U91 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U92 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n79, ZN => n152);
   U93 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U94 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U95 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n79, ZN => n154);
   U96 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U97 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U98 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n79, ZN => n156);
   U99 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U100 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U101 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n79, ZN => n158);
   U102 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U103 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U104 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n79, ZN => n165);
   U105 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U106 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n115);
   U107 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U108 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U109 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n99);
   U110 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U111 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U112 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n101);
   U113 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U114 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U115 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n103);
   U116 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U117 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U118 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n105);
   U119 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U120 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U121 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n107);
   U122 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U123 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U124 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n109);
   U125 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U126 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U127 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n111);
   U128 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U129 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U130 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n113);
   U131 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_3 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_3;

architecture SYN_Behavioral of MUX5to1_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U37 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U38 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n120);
   U39 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U40 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U41 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U42 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U43 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U44 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U45 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U46 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U47 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U48 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U49 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U50 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U51 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U52 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U53 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U54 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U55 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U56 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U57 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U58 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U59 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U60 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U61 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U62 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U63 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U64 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U65 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U66 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U67 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U68 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U69 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U70 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U71 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U72 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U73 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U74 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U75 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U76 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U77 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n79, ZN => n146);
   U78 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U79 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U80 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n79, ZN => n148);
   U81 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U82 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U83 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n79, ZN => n150);
   U84 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U85 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U86 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n79, ZN => n152);
   U87 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U88 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U89 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n79, ZN => n154);
   U90 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U91 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U92 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n79, ZN => n156);
   U93 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U94 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U95 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, C1
                           => D(30), C2 => n79, ZN => n158);
   U96 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U97 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U98 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, C1
                           => D(31), C2 => n79, ZN => n165);
   U99 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U100 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U101 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, 
                           C1 => D(10), C2 => n80, ZN => n118);
   U102 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U103 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n99);
   U104 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U105 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U106 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n101);
   U107 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U108 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U109 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n103);
   U110 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U111 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U112 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n105);
   U113 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U114 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U115 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n107);
   U116 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U117 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U118 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n109);
   U119 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U120 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U121 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n111);
   U122 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U123 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U124 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n113);
   U125 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U126 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U127 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n115);
   U128 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U129 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U130 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN =>
                           n117);
   U131 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_2 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_2;

architecture SYN_Behavioral of MUX5to1_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U37 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U38 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n124);
   U39 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U40 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U41 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U42 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U43 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U44 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U45 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U46 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U47 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U48 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U49 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U50 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U51 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U52 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U53 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U54 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U55 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U56 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U57 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U58 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U59 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U60 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U61 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U62 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U63 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U64 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U65 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U66 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U67 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U68 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U69 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U70 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U71 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n79, ZN => n146);
   U72 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U73 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U74 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n79, ZN => n148);
   U75 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U76 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U77 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n79, ZN => n150);
   U78 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U79 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U80 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n79, ZN => n152);
   U81 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U82 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U83 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n79, ZN => n154);
   U84 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U85 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U86 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n79, ZN => n156);
   U87 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U88 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U89 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, C1
                           => D(30), C2 => n79, ZN => n158);
   U90 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U91 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U92 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, C1
                           => D(31), C2 => n79, ZN => n165);
   U93 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U94 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U95 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n122);
   U96 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U97 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN =>
                           n99);
   U98 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U99 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U100 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n101);
   U101 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U102 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U103 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n103);
   U104 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U105 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U106 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n105);
   U107 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U108 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U109 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n107);
   U110 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U111 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U112 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n109);
   U113 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U114 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U115 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n111);
   U116 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U117 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U118 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n113);
   U119 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U120 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U121 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n115);
   U122 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U123 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U124 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN =>
                           n117);
   U125 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U126 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U127 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U128 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, 
                           C1 => D(10), C2 => n80, ZN => n118);
   U129 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U130 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U131 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, 
                           C1 => D(11), C2 => n80, ZN => n120);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_1 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_1;

architecture SYN_Behavioral of MUX5to1_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n162, Z => n82);
   U5 : BUF_X1 port map( A => n161, Z => n78);
   U6 : BUF_X1 port map( A => n163, Z => n83);
   U7 : BUF_X1 port map( A => n164, Z => n90);
   U8 : BUF_X1 port map( A => n160, Z => n74);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n97, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n97);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n83, Z => n85);
   U17 : BUF_X1 port map( A => n83, Z => n84);
   U18 : BUF_X1 port map( A => n82, Z => n80);
   U19 : BUF_X1 port map( A => n82, Z => n79);
   U20 : BUF_X1 port map( A => n78, Z => n77);
   U21 : BUF_X1 port map( A => n83, Z => n86);
   U22 : BUF_X1 port map( A => n82, Z => n81);
   U23 : INV_X1 port map( A => SEL(1), ZN => n95);
   U24 : NOR3_X1 port map( A1 => n96, A2 => SEL(2), A3 => n95, ZN => n162);
   U25 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n96, ZN => n161);
   U26 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => SEL(2), ZN => n163);
   U27 : BUF_X1 port map( A => n74, Z => n2);
   U28 : BUF_X1 port map( A => n74, Z => n1);
   U29 : BUF_X1 port map( A => n90, Z => n88);
   U30 : BUF_X1 port map( A => n90, Z => n87);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : INV_X1 port map( A => SEL(0), ZN => n96);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n95, ZN => n164);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n160
                           );
   U36 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N41);
   U37 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n129);
   U38 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n128);
   U39 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N42);
   U40 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n131);
   U41 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n130);
   U42 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N43);
   U43 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n133);
   U44 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n132);
   U45 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N44);
   U46 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n135);
   U47 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n134);
   U48 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N45);
   U49 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n137);
   U50 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n136);
   U51 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N46);
   U52 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n139);
   U53 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n138);
   U54 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N47);
   U55 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n141);
   U56 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n79, ZN => n140);
   U57 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N48);
   U58 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n143);
   U59 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n79, ZN => n142);
   U60 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N49);
   U61 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n145);
   U62 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n79, ZN => n144);
   U63 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N50);
   U64 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n147);
   U65 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n79, ZN => n146);
   U66 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N51);
   U67 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n149);
   U68 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n79, ZN => n148);
   U69 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N52);
   U70 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n151);
   U71 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n79, ZN => n150);
   U72 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N53);
   U73 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n153);
   U74 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n79, ZN => n152);
   U75 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N54);
   U76 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n155);
   U77 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n79, ZN => n154);
   U78 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N55);
   U79 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n157);
   U80 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n79, ZN => n156);
   U81 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N56);
   U82 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n159);
   U83 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, C1
                           => D(30), C2 => n79, ZN => n158);
   U84 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => N57);
   U85 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n166);
   U86 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, C1
                           => D(31), C2 => n79, ZN => n165);
   U87 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N40);
   U88 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n127);
   U89 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n126);
   U90 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => N26);
   U91 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN =>
                           n99);
   U92 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n98);
   U93 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N27);
   U94 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN =>
                           n101);
   U95 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n100);
   U96 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N28);
   U97 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN =>
                           n103);
   U98 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n102);
   U99 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N29);
   U100 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n105);
   U101 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n104);
   U102 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N30);
   U103 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n107);
   U104 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n106);
   U105 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N31);
   U106 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n109);
   U107 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n108);
   U108 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N32);
   U109 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n111);
   U110 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n110);
   U111 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N33);
   U112 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n113);
   U113 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n112);
   U114 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N34);
   U115 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n115);
   U116 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n114);
   U117 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N35);
   U118 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN =>
                           n117);
   U119 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n116);
   U120 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N36);
   U121 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n119);
   U122 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, 
                           C1 => D(10), C2 => n80, ZN => n118);
   U123 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N37);
   U124 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n121);
   U125 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, 
                           C1 => D(11), C2 => n80, ZN => n120);
   U126 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N38);
   U127 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n123);
   U128 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, 
                           C1 => D(12), C2 => n80, ZN => n122);
   U129 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N39);
   U130 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n125);
   U131 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, 
                           C1 => D(13), C2 => n80, ZN => n124);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_8 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_8;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n80, ZN => Y(1));
   U2 : BUF_X1 port map( A => n68, Z => n1);
   U3 : BUF_X1 port map( A => n68, Z => n2);
   U4 : BUF_X1 port map( A => n68, Z => n3);
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => SEL, ZN => 
                           n80);
   U6 : INV_X1 port map( A => n91, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => SEL, ZN => 
                           n91);
   U8 : INV_X1 port map( A => n94, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => SEL, ZN => 
                           n94);
   U10 : INV_X1 port map( A => n95, ZN => Y(4));
   U11 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => SEL, ZN => 
                           n95);
   U12 : INV_X1 port map( A => n96, ZN => Y(5));
   U13 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => SEL, ZN => 
                           n96);
   U14 : INV_X1 port map( A => n97, ZN => Y(6));
   U15 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => SEL, ZN => 
                           n97);
   U16 : INV_X1 port map( A => n98, ZN => Y(7));
   U17 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => SEL, ZN => 
                           n98);
   U18 : INV_X1 port map( A => n99, ZN => Y(8));
   U19 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => SEL, ZN => 
                           n99);
   U20 : INV_X1 port map( A => n100, ZN => Y(9));
   U21 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => SEL, B2 => B(9), ZN => 
                           n100);
   U22 : INV_X1 port map( A => n70, ZN => Y(10));
   U23 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => SEL, ZN 
                           => n70);
   U24 : INV_X1 port map( A => n71, ZN => Y(11));
   U25 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => SEL, ZN 
                           => n71);
   U26 : INV_X1 port map( A => n72, ZN => Y(12));
   U27 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => SEL, ZN 
                           => n72);
   U28 : INV_X1 port map( A => n73, ZN => Y(13));
   U29 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => SEL, ZN 
                           => n73);
   U30 : INV_X1 port map( A => n74, ZN => Y(14));
   U31 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => SEL, ZN 
                           => n74);
   U32 : INV_X1 port map( A => n75, ZN => Y(15));
   U33 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => SEL, ZN 
                           => n75);
   U34 : INV_X1 port map( A => n76, ZN => Y(16));
   U35 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => SEL, ZN 
                           => n76);
   U36 : INV_X1 port map( A => n77, ZN => Y(17));
   U37 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => SEL, ZN 
                           => n77);
   U38 : INV_X1 port map( A => n78, ZN => Y(18));
   U39 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => SEL, ZN 
                           => n78);
   U40 : INV_X1 port map( A => n79, ZN => Y(19));
   U41 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => SEL, ZN 
                           => n79);
   U42 : INV_X1 port map( A => n81, ZN => Y(20));
   U43 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => SEL, ZN 
                           => n81);
   U44 : INV_X1 port map( A => n82, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => SEL, ZN 
                           => n82);
   U46 : INV_X1 port map( A => n83, ZN => Y(22));
   U47 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => SEL, ZN 
                           => n83);
   U48 : INV_X1 port map( A => n84, ZN => Y(23));
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => SEL, ZN 
                           => n84);
   U50 : INV_X1 port map( A => n85, ZN => Y(24));
   U51 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => SEL, ZN 
                           => n85);
   U52 : INV_X1 port map( A => n86, ZN => Y(25));
   U53 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => SEL, ZN 
                           => n86);
   U54 : INV_X1 port map( A => n87, ZN => Y(26));
   U55 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => SEL, ZN 
                           => n87);
   U56 : INV_X1 port map( A => n88, ZN => Y(27));
   U57 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => SEL, ZN 
                           => n88);
   U58 : INV_X1 port map( A => n89, ZN => Y(28));
   U59 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => SEL, ZN 
                           => n89);
   U60 : INV_X1 port map( A => n90, ZN => Y(29));
   U61 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => SEL, ZN 
                           => n90);
   U62 : INV_X1 port map( A => n92, ZN => Y(30));
   U63 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => SEL, ZN 
                           => n92);
   U64 : INV_X1 port map( A => n69, ZN => Y(0));
   U65 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => SEL, ZN => 
                           n69);
   U66 : INV_X1 port map( A => SEL, ZN => n68);
   U67 : INV_X1 port map( A => n93, ZN => Y(31));
   U68 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => SEL, ZN 
                           => n93);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_7;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n1);
   U2 : CLKBUF_X1 port map( A => n4, Z => n2);
   U3 : CLKBUF_X1 port map( A => n4, Z => n3);
   U4 : BUF_X1 port map( A => SEL, Z => n4);
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U6 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U7 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U8 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U9 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U10 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U11 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U12 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U13 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U14 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U15 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U16 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U17 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U18 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U19 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U20 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U21 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U22 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U23 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U24 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U25 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U26 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U27 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U28 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U29 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U30 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U31 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U32 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U33 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U34 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U35 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U36 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_6;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n1);
   U2 : BUF_X1 port map( A => n4, Z => n2);
   U3 : BUF_X1 port map( A => n4, Z => n3);
   U4 : BUF_X1 port map( A => SEL, Z => n4);
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U6 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U7 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U8 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U9 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U10 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U11 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U12 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U13 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U14 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U15 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U16 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U17 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U18 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U19 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U20 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U21 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U22 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U23 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U24 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U25 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U26 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U27 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U28 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U29 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U30 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U31 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U32 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U33 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U34 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U35 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U36 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_5;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U4 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U5 : MUX2_X1 port map( A => A(2), B => B(2), S => n2, Z => Y(2));
   U6 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U7 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U8 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U9 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U10 : MUX2_X1 port map( A => A(7), B => B(7), S => n2, Z => Y(7));
   U11 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U12 : MUX2_X1 port map( A => A(9), B => B(9), S => n2, Z => Y(9));
   U13 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U14 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U15 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U16 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U17 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U18 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U19 : MUX2_X1 port map( A => A(16), B => B(16), S => n1, Z => Y(16));
   U20 : MUX2_X1 port map( A => A(17), B => B(17), S => n1, Z => Y(17));
   U21 : MUX2_X1 port map( A => A(18), B => B(18), S => n1, Z => Y(18));
   U22 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U23 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U24 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U25 : MUX2_X1 port map( A => A(22), B => B(22), S => n1, Z => Y(22));
   U26 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U27 : MUX2_X1 port map( A => A(24), B => B(24), S => n1, Z => Y(24));
   U28 : MUX2_X1 port map( A => A(25), B => B(25), S => n2, Z => Y(25));
   U29 : MUX2_X1 port map( A => A(26), B => B(26), S => n1, Z => Y(26));
   U30 : MUX2_X1 port map( A => A(27), B => B(27), S => n2, Z => Y(27));
   U31 : MUX2_X1 port map( A => A(28), B => B(28), S => n2, Z => Y(28));
   U32 : MUX2_X1 port map( A => A(29), B => B(29), S => n2, Z => Y(29));
   U33 : MUX2_X1 port map( A => A(30), B => B(30), S => n1, Z => Y(30));
   U34 : MUX2_X1 port map( A => A(31), B => B(31), S => n1, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_4;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n7);
   U2 : BUF_X1 port map( A => n4, Z => n8);
   U3 : BUF_X1 port map( A => n8, Z => n1);
   U4 : BUF_X1 port map( A => n8, Z => n2);
   U5 : INV_X1 port map( A => n7, ZN => n5);
   U6 : INV_X1 port map( A => n7, ZN => n6);
   U7 : BUF_X1 port map( A => n8, Z => n3);
   U8 : BUF_X1 port map( A => SEL, Z => n4);
   U9 : INV_X1 port map( A => n73, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n73);
   U11 : INV_X1 port map( A => n84, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U13 : INV_X1 port map( A => n95, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U15 : INV_X1 port map( A => n98, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U17 : INV_X1 port map( A => n99, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U19 : INV_X1 port map( A => n100, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U21 : INV_X1 port map( A => n101, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U23 : INV_X1 port map( A => n102, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U25 : INV_X1 port map( A => n103, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U27 : INV_X1 port map( A => n104, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U29 : INV_X1 port map( A => n74, ZN => Y(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U31 : INV_X1 port map( A => n75, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U33 : INV_X1 port map( A => n76, ZN => Y(12));
   U34 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U35 : INV_X1 port map( A => n77, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U37 : INV_X1 port map( A => n78, ZN => Y(14));
   U38 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U39 : INV_X1 port map( A => n79, ZN => Y(15));
   U40 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U41 : INV_X1 port map( A => n80, ZN => Y(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U43 : INV_X1 port map( A => n81, ZN => Y(17));
   U44 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U45 : INV_X1 port map( A => n82, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U47 : INV_X1 port map( A => n83, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U49 : INV_X1 port map( A => n85, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U51 : INV_X1 port map( A => n86, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U53 : INV_X1 port map( A => n87, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U55 : INV_X1 port map( A => n88, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U57 : INV_X1 port map( A => n89, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U59 : INV_X1 port map( A => n90, ZN => Y(25));
   U60 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U61 : INV_X1 port map( A => n91, ZN => Y(26));
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U63 : INV_X1 port map( A => n92, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U65 : INV_X1 port map( A => n93, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U67 : INV_X1 port map( A => n94, ZN => Y(29));
   U68 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U69 : INV_X1 port map( A => n96, ZN => Y(30));
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U71 : INV_X1 port map( A => n97, ZN => Y(31));
   U72 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n3, ZN =>
                           n97);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_3;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n9);
   U2 : BUF_X1 port map( A => n4, Z => n8);
   U3 : BUF_X1 port map( A => SEL, Z => n4);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : BUF_X1 port map( A => n9, Z => n1);
   U8 : BUF_X1 port map( A => n9, Z => n3);
   U9 : BUF_X1 port map( A => n9, Z => n2);
   U10 : INV_X1 port map( A => n103, ZN => Y(7));
   U11 : AOI22_X1 port map( A1 => A(7), A2 => n7, B1 => B(7), B2 => n3, ZN => 
                           n103);
   U12 : INV_X1 port map( A => n75, ZN => Y(10));
   U13 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n75);
   U14 : INV_X1 port map( A => n76, ZN => Y(11));
   U15 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n76);
   U16 : INV_X1 port map( A => n77, ZN => Y(12));
   U17 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n77);
   U18 : INV_X1 port map( A => n78, ZN => Y(13));
   U19 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n78);
   U20 : INV_X1 port map( A => n79, ZN => Y(14));
   U21 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n79);
   U22 : INV_X1 port map( A => n80, ZN => Y(15));
   U23 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n80);
   U24 : INV_X1 port map( A => n81, ZN => Y(16));
   U25 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n81);
   U26 : INV_X1 port map( A => n82, ZN => Y(17));
   U27 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n82);
   U28 : INV_X1 port map( A => n83, ZN => Y(18));
   U29 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n83);
   U30 : INV_X1 port map( A => n84, ZN => Y(19));
   U31 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n84);
   U32 : INV_X1 port map( A => n86, ZN => Y(20));
   U33 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n86);
   U34 : INV_X1 port map( A => n87, ZN => Y(21));
   U35 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n87);
   U36 : INV_X1 port map( A => n88, ZN => Y(22));
   U37 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n88);
   U38 : INV_X1 port map( A => n89, ZN => Y(23));
   U39 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n89);
   U40 : INV_X1 port map( A => n90, ZN => Y(24));
   U41 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n90);
   U42 : INV_X1 port map( A => n91, ZN => Y(25));
   U43 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n91);
   U44 : INV_X1 port map( A => n92, ZN => Y(26));
   U45 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n92);
   U46 : INV_X1 port map( A => n93, ZN => Y(27));
   U47 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n93);
   U48 : INV_X1 port map( A => n94, ZN => Y(28));
   U49 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n94);
   U50 : INV_X1 port map( A => n95, ZN => Y(29));
   U51 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n95);
   U52 : INV_X1 port map( A => n97, ZN => Y(30));
   U53 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n97);
   U54 : INV_X1 port map( A => n98, ZN => Y(31));
   U55 : AOI22_X1 port map( A1 => A(31), A2 => n7, B1 => B(31), B2 => n3, ZN =>
                           n98);
   U56 : INV_X1 port map( A => n105, ZN => Y(9));
   U57 : AOI22_X1 port map( A1 => A(9), A2 => n7, B1 => n3, B2 => B(9), ZN => 
                           n105);
   U58 : INV_X1 port map( A => n85, ZN => Y(1));
   U59 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n85);
   U60 : INV_X1 port map( A => n96, ZN => Y(2));
   U61 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n96);
   U62 : INV_X1 port map( A => n99, ZN => Y(3));
   U63 : AOI22_X1 port map( A1 => A(3), A2 => n7, B1 => B(3), B2 => n3, ZN => 
                           n99);
   U64 : INV_X1 port map( A => n100, ZN => Y(4));
   U65 : AOI22_X1 port map( A1 => A(4), A2 => n7, B1 => B(4), B2 => n3, ZN => 
                           n100);
   U66 : INV_X1 port map( A => n101, ZN => Y(5));
   U67 : AOI22_X1 port map( A1 => A(5), A2 => n7, B1 => B(5), B2 => n3, ZN => 
                           n101);
   U68 : INV_X1 port map( A => n102, ZN => Y(6));
   U69 : AOI22_X1 port map( A1 => A(6), A2 => n7, B1 => B(6), B2 => n3, ZN => 
                           n102);
   U70 : INV_X1 port map( A => n104, ZN => Y(8));
   U71 : AOI22_X1 port map( A1 => A(8), A2 => n7, B1 => B(8), B2 => n3, ZN => 
                           n104);
   U72 : INV_X1 port map( A => n74, ZN => Y(0));
   U73 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n74);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_2;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n7);
   U2 : BUF_X1 port map( A => n4, Z => n8);
   U3 : BUF_X1 port map( A => n8, Z => n1);
   U4 : BUF_X1 port map( A => n8, Z => n2);
   U5 : INV_X1 port map( A => n7, ZN => n5);
   U6 : INV_X1 port map( A => n7, ZN => n6);
   U7 : BUF_X1 port map( A => n8, Z => n3);
   U8 : BUF_X1 port map( A => SEL, Z => n4);
   U9 : INV_X1 port map( A => n73, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n73);
   U11 : INV_X1 port map( A => n84, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U13 : INV_X1 port map( A => n95, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U15 : INV_X1 port map( A => n98, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U17 : INV_X1 port map( A => n99, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U19 : INV_X1 port map( A => n100, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U21 : INV_X1 port map( A => n101, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U23 : INV_X1 port map( A => n102, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U25 : INV_X1 port map( A => n103, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U27 : INV_X1 port map( A => n104, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U29 : INV_X1 port map( A => n74, ZN => Y(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U31 : INV_X1 port map( A => n75, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U33 : INV_X1 port map( A => n76, ZN => Y(12));
   U34 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U35 : INV_X1 port map( A => n77, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U37 : INV_X1 port map( A => n78, ZN => Y(14));
   U38 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U39 : INV_X1 port map( A => n79, ZN => Y(15));
   U40 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U41 : INV_X1 port map( A => n80, ZN => Y(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U43 : INV_X1 port map( A => n81, ZN => Y(17));
   U44 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U45 : INV_X1 port map( A => n82, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U47 : INV_X1 port map( A => n83, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U49 : INV_X1 port map( A => n85, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U51 : INV_X1 port map( A => n86, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U53 : INV_X1 port map( A => n87, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U55 : INV_X1 port map( A => n88, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U57 : INV_X1 port map( A => n89, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U59 : INV_X1 port map( A => n90, ZN => Y(25));
   U60 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U61 : INV_X1 port map( A => n91, ZN => Y(26));
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U63 : INV_X1 port map( A => n92, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U65 : INV_X1 port map( A => n93, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U67 : INV_X1 port map( A => n94, ZN => Y(29));
   U68 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U69 : INV_X1 port map( A => n96, ZN => Y(30));
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U71 : INV_X1 port map( A => n97, ZN => Y(31));
   U72 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n3, ZN =>
                           n97);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_1;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => SEL, Z => n4);
   U2 : BUF_X2 port map( A => n4, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n9);
   U4 : INV_X1 port map( A => n8, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : BUF_X1 port map( A => n9, Z => n3);
   U8 : BUF_X1 port map( A => n9, Z => n1);
   U9 : BUF_X1 port map( A => n9, Z => n2);
   U10 : INV_X1 port map( A => n105, ZN => Y(9));
   U11 : AOI22_X1 port map( A1 => A(9), A2 => n7, B1 => n3, B2 => B(9), ZN => 
                           n105);
   U12 : INV_X1 port map( A => n99, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n7, B1 => B(3), B2 => n3, ZN => 
                           n99);
   U14 : INV_X1 port map( A => n100, ZN => Y(4));
   U15 : AOI22_X1 port map( A1 => A(4), A2 => n7, B1 => B(4), B2 => n3, ZN => 
                           n100);
   U16 : INV_X1 port map( A => n101, ZN => Y(5));
   U17 : AOI22_X1 port map( A1 => A(5), A2 => n7, B1 => B(5), B2 => n3, ZN => 
                           n101);
   U18 : INV_X1 port map( A => n102, ZN => Y(6));
   U19 : AOI22_X1 port map( A1 => A(6), A2 => n7, B1 => B(6), B2 => n3, ZN => 
                           n102);
   U20 : INV_X1 port map( A => n103, ZN => Y(7));
   U21 : AOI22_X1 port map( A1 => A(7), A2 => n7, B1 => B(7), B2 => n3, ZN => 
                           n103);
   U22 : INV_X1 port map( A => n104, ZN => Y(8));
   U23 : AOI22_X1 port map( A1 => A(8), A2 => n7, B1 => B(8), B2 => n3, ZN => 
                           n104);
   U24 : INV_X1 port map( A => n98, ZN => Y(31));
   U25 : AOI22_X1 port map( A1 => A(31), A2 => n7, B1 => B(31), B2 => n3, ZN =>
                           n98);
   U26 : INV_X1 port map( A => n74, ZN => Y(0));
   U27 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n74);
   U28 : INV_X1 port map( A => n85, ZN => Y(1));
   U29 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n85);
   U30 : INV_X1 port map( A => n96, ZN => Y(2));
   U31 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n96);
   U32 : INV_X1 port map( A => n75, ZN => Y(10));
   U33 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n75);
   U34 : INV_X1 port map( A => n76, ZN => Y(11));
   U35 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n76);
   U36 : INV_X1 port map( A => n77, ZN => Y(12));
   U37 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n77);
   U38 : INV_X1 port map( A => n78, ZN => Y(13));
   U39 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n78);
   U40 : INV_X1 port map( A => n79, ZN => Y(14));
   U41 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n79);
   U42 : INV_X1 port map( A => n80, ZN => Y(15));
   U43 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n80);
   U44 : INV_X1 port map( A => n81, ZN => Y(16));
   U45 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n81);
   U46 : INV_X1 port map( A => n82, ZN => Y(17));
   U47 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n82);
   U48 : INV_X1 port map( A => n83, ZN => Y(18));
   U49 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n83);
   U50 : INV_X1 port map( A => n84, ZN => Y(19));
   U51 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n84);
   U52 : INV_X1 port map( A => n86, ZN => Y(20));
   U53 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n86);
   U54 : INV_X1 port map( A => n87, ZN => Y(21));
   U55 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n87);
   U56 : INV_X1 port map( A => n88, ZN => Y(22));
   U57 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n88);
   U58 : INV_X1 port map( A => n89, ZN => Y(23));
   U59 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n89);
   U60 : INV_X1 port map( A => n90, ZN => Y(24));
   U61 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n90);
   U62 : INV_X1 port map( A => n91, ZN => Y(25));
   U63 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n91);
   U64 : INV_X1 port map( A => n92, ZN => Y(26));
   U65 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n92);
   U66 : INV_X1 port map( A => n93, ZN => Y(27));
   U67 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n93);
   U68 : INV_X1 port map( A => n94, ZN => Y(28));
   U69 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n94);
   U70 : INV_X1 port map( A => n95, ZN => Y(29));
   U71 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n95);
   U72 : INV_X1 port map( A => n97, ZN => Y(30));
   U73 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n97);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_3 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_3;

architecture SYN_Behavioral of MUX3to1_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12_port, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n16, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n17, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n18, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n27, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n28, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n73, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U4 : BUF_X1 port map( A => n117, Z => n12_port);
   U5 : BUF_X1 port map( A => n116, Z => n8);
   U6 : BUF_X1 port map( A => n115, Z => n1);
   U7 : BUF_X1 port map( A => N12, Z => n14);
   U8 : BUF_X1 port map( A => N12, Z => n13);
   U9 : BUF_X1 port map( A => N12, Z => n15);
   U10 : BUF_X1 port map( A => n8, Z => n6);
   U11 : BUF_X1 port map( A => n8, Z => n5);
   U12 : BUF_X1 port map( A => n1, Z => n2);
   U13 : BUF_X1 port map( A => n1, Z => n3);
   U14 : BUF_X1 port map( A => n12_port, Z => n9);
   U15 : BUF_X1 port map( A => n12_port, Z => n10);
   U16 : BUF_X1 port map( A => n8, Z => n7);
   U17 : BUF_X1 port map( A => n1, Z => n4);
   U18 : BUF_X1 port map( A => n12_port, Z => n11);
   U19 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n117);
   U20 : NOR2_X1 port map( A1 => n83, A2 => SEL(0), ZN => n116);
   U21 : AND2_X1 port map( A1 => SEL(0), A2 => n83, ZN => n115);
   U22 : INV_X1 port map( A => SEL(1), ZN => n83);
   U23 : INV_X1 port map( A => n84, ZN => n82);
   U24 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n84);
   U25 : INV_X1 port map( A => n85, ZN => n81);
   U26 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n85);
   U27 : INV_X1 port map( A => n86, ZN => n80);
   U28 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n86);
   U29 : INV_X1 port map( A => n87, ZN => n79);
   U30 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n87);
   U31 : INV_X1 port map( A => n88, ZN => n78);
   U32 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n88);
   U33 : INV_X1 port map( A => n89, ZN => n77);
   U34 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n89);
   U35 : INV_X1 port map( A => n90, ZN => n76);
   U36 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n90);
   U37 : INV_X1 port map( A => n91, ZN => n75);
   U38 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n91);
   U39 : INV_X1 port map( A => n92, ZN => n74);
   U40 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n92);
   U41 : INV_X1 port map( A => n93, ZN => n73);
   U42 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n93);
   U43 : INV_X1 port map( A => n94, ZN => n72);
   U44 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n94);
   U45 : INV_X1 port map( A => n95, ZN => n71);
   U46 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n95);
   U47 : INV_X1 port map( A => n96, ZN => n70);
   U48 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n96);
   U49 : INV_X1 port map( A => n97, ZN => n69);
   U50 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n97);
   U51 : INV_X1 port map( A => n98, ZN => n33);
   U52 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n98);
   U53 : INV_X1 port map( A => n99, ZN => n32);
   U54 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n99);
   U55 : INV_X1 port map( A => n100, ZN => n31);
   U56 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n100);
   U57 : INV_X1 port map( A => n101, ZN => n30);
   U58 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n101);
   U59 : INV_X1 port map( A => n102, ZN => n29);
   U60 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n102);
   U61 : INV_X1 port map( A => n103, ZN => n28);
   U62 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n103);
   U63 : INV_X1 port map( A => n104, ZN => n27);
   U64 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n104);
   U65 : INV_X1 port map( A => n105, ZN => n26);
   U66 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n105);
   U67 : INV_X1 port map( A => n106, ZN => n25);
   U68 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n106);
   U69 : INV_X1 port map( A => n107, ZN => n24);
   U70 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n107);
   U71 : INV_X1 port map( A => n108, ZN => n23);
   U72 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n108);
   U73 : INV_X1 port map( A => n109, ZN => n22);
   U74 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n109);
   U75 : INV_X1 port map( A => n110, ZN => n21);
   U76 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n110);
   U77 : INV_X1 port map( A => n111, ZN => n20);
   U78 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n111);
   U79 : INV_X1 port map( A => n112, ZN => n19);
   U80 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n112);
   U81 : INV_X1 port map( A => n113, ZN => n18);
   U82 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n113);
   U83 : INV_X1 port map( A => n114, ZN => n17);
   U84 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n114);
   U85 : INV_X1 port map( A => n118, ZN => n16);
   U86 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n118);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_2 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_2;

architecture SYN_Behavioral of MUX3to1_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12_port, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n16, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n17, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n18, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n27, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n28, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n73, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U4 : BUF_X1 port map( A => n117, Z => n12_port);
   U5 : BUF_X1 port map( A => n116, Z => n8);
   U6 : BUF_X1 port map( A => n115, Z => n1);
   U7 : BUF_X1 port map( A => N12, Z => n14);
   U8 : BUF_X1 port map( A => N12, Z => n13);
   U9 : BUF_X1 port map( A => N12, Z => n15);
   U10 : BUF_X1 port map( A => n8, Z => n6);
   U11 : BUF_X1 port map( A => n8, Z => n5);
   U12 : BUF_X1 port map( A => n1, Z => n2);
   U13 : BUF_X1 port map( A => n1, Z => n3);
   U14 : BUF_X1 port map( A => n12_port, Z => n9);
   U15 : BUF_X1 port map( A => n12_port, Z => n10);
   U16 : BUF_X1 port map( A => n8, Z => n7);
   U17 : BUF_X1 port map( A => n1, Z => n4);
   U18 : BUF_X1 port map( A => n12_port, Z => n11);
   U19 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n117);
   U20 : NOR2_X1 port map( A1 => n83, A2 => SEL(0), ZN => n116);
   U21 : AND2_X1 port map( A1 => SEL(0), A2 => n83, ZN => n115);
   U22 : INV_X1 port map( A => SEL(1), ZN => n83);
   U23 : INV_X1 port map( A => n84, ZN => n82);
   U24 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n84);
   U25 : INV_X1 port map( A => n85, ZN => n81);
   U26 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n85);
   U27 : INV_X1 port map( A => n86, ZN => n80);
   U28 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n86);
   U29 : INV_X1 port map( A => n87, ZN => n79);
   U30 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n87);
   U31 : INV_X1 port map( A => n88, ZN => n78);
   U32 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n88);
   U33 : INV_X1 port map( A => n89, ZN => n77);
   U34 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n89);
   U35 : INV_X1 port map( A => n90, ZN => n76);
   U36 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n90);
   U37 : INV_X1 port map( A => n91, ZN => n75);
   U38 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n91);
   U39 : INV_X1 port map( A => n92, ZN => n74);
   U40 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n92);
   U41 : INV_X1 port map( A => n93, ZN => n73);
   U42 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n93);
   U43 : INV_X1 port map( A => n94, ZN => n72);
   U44 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n94);
   U45 : INV_X1 port map( A => n95, ZN => n71);
   U46 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n95);
   U47 : INV_X1 port map( A => n96, ZN => n70);
   U48 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n96);
   U49 : INV_X1 port map( A => n97, ZN => n69);
   U50 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n97);
   U51 : INV_X1 port map( A => n98, ZN => n33);
   U52 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n98);
   U53 : INV_X1 port map( A => n99, ZN => n32);
   U54 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n99);
   U55 : INV_X1 port map( A => n100, ZN => n31);
   U56 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n100);
   U57 : INV_X1 port map( A => n101, ZN => n30);
   U58 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n101);
   U59 : INV_X1 port map( A => n102, ZN => n29);
   U60 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n102);
   U61 : INV_X1 port map( A => n103, ZN => n28);
   U62 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n103);
   U63 : INV_X1 port map( A => n104, ZN => n27);
   U64 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n104);
   U65 : INV_X1 port map( A => n105, ZN => n26);
   U66 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n105);
   U67 : INV_X1 port map( A => n106, ZN => n25);
   U68 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n106);
   U69 : INV_X1 port map( A => n107, ZN => n24);
   U70 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n107);
   U71 : INV_X1 port map( A => n108, ZN => n23);
   U72 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n108);
   U73 : INV_X1 port map( A => n109, ZN => n22);
   U74 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n109);
   U75 : INV_X1 port map( A => n110, ZN => n21);
   U76 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n110);
   U77 : INV_X1 port map( A => n111, ZN => n20);
   U78 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n111);
   U79 : INV_X1 port map( A => n112, ZN => n19);
   U80 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n112);
   U81 : INV_X1 port map( A => n113, ZN => n18);
   U82 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n113);
   U83 : INV_X1 port map( A => n114, ZN => n17);
   U84 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n114);
   U85 : INV_X1 port map( A => n118, ZN => n16);
   U86 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n118);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_1 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_1;

architecture SYN_Behavioral of MUX3to1_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12_port, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n16, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n17, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n18, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n27, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n28, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n73, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U4 : BUF_X1 port map( A => n117, Z => n12_port);
   U5 : BUF_X1 port map( A => n116, Z => n8);
   U6 : BUF_X1 port map( A => n115, Z => n1);
   U7 : BUF_X1 port map( A => N12, Z => n14);
   U8 : BUF_X1 port map( A => N12, Z => n13);
   U9 : BUF_X1 port map( A => N12, Z => n15);
   U10 : BUF_X1 port map( A => n8, Z => n6);
   U11 : BUF_X1 port map( A => n8, Z => n5);
   U12 : BUF_X1 port map( A => n1, Z => n2);
   U13 : BUF_X1 port map( A => n1, Z => n3);
   U14 : BUF_X1 port map( A => n12_port, Z => n9);
   U15 : BUF_X1 port map( A => n12_port, Z => n10);
   U16 : BUF_X1 port map( A => n8, Z => n7);
   U17 : BUF_X1 port map( A => n1, Z => n4);
   U18 : BUF_X1 port map( A => n12_port, Z => n11);
   U19 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n117);
   U20 : NOR2_X1 port map( A1 => n83, A2 => SEL(0), ZN => n116);
   U21 : INV_X1 port map( A => SEL(1), ZN => n83);
   U22 : AND2_X1 port map( A1 => SEL(0), A2 => n83, ZN => n115);
   U23 : INV_X1 port map( A => n84, ZN => n82);
   U24 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n84);
   U25 : INV_X1 port map( A => n85, ZN => n81);
   U26 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n85);
   U27 : INV_X1 port map( A => n86, ZN => n80);
   U28 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n86);
   U29 : INV_X1 port map( A => n87, ZN => n79);
   U30 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n87);
   U31 : INV_X1 port map( A => n88, ZN => n78);
   U32 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n88);
   U33 : INV_X1 port map( A => n89, ZN => n77);
   U34 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n89);
   U35 : INV_X1 port map( A => n90, ZN => n76);
   U36 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n90);
   U37 : INV_X1 port map( A => n91, ZN => n75);
   U38 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n91);
   U39 : INV_X1 port map( A => n92, ZN => n74);
   U40 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n92);
   U41 : INV_X1 port map( A => n93, ZN => n73);
   U42 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n93);
   U43 : INV_X1 port map( A => n94, ZN => n72);
   U44 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n94);
   U45 : INV_X1 port map( A => n95, ZN => n71);
   U46 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n95);
   U47 : INV_X1 port map( A => n96, ZN => n70);
   U48 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n96);
   U49 : INV_X1 port map( A => n97, ZN => n69);
   U50 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n97);
   U51 : INV_X1 port map( A => n98, ZN => n33);
   U52 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n98);
   U53 : INV_X1 port map( A => n99, ZN => n32);
   U54 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n99);
   U55 : INV_X1 port map( A => n100, ZN => n31);
   U56 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n100);
   U57 : INV_X1 port map( A => n101, ZN => n30);
   U58 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n101);
   U59 : INV_X1 port map( A => n102, ZN => n29);
   U60 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n102);
   U61 : INV_X1 port map( A => n103, ZN => n28);
   U62 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n103);
   U63 : INV_X1 port map( A => n104, ZN => n27);
   U64 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n104);
   U65 : INV_X1 port map( A => n105, ZN => n26);
   U66 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n105);
   U67 : INV_X1 port map( A => n106, ZN => n25);
   U68 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n106);
   U69 : INV_X1 port map( A => n107, ZN => n24);
   U70 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n107);
   U71 : INV_X1 port map( A => n108, ZN => n23);
   U72 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n108);
   U73 : INV_X1 port map( A => n109, ZN => n22);
   U74 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n109);
   U75 : INV_X1 port map( A => n110, ZN => n21);
   U76 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n110);
   U77 : INV_X1 port map( A => n111, ZN => n20);
   U78 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n111);
   U79 : INV_X1 port map( A => n112, ZN => n19);
   U80 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n112);
   U81 : INV_X1 port map( A => n113, ZN => n18);
   U82 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n113);
   U83 : INV_X1 port map( A => n114, ZN => n17);
   U84 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n114);
   U85 : INV_X1 port map( A => n118, ZN => n16);
   U86 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n118);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Sum : out std_logic_vector 
         (31 downto 0));

end PC_adder_1;

architecture SYN_Behavioral of PC_adder_1 is

   component PC_adder_1_DW01_add_0_DW01_add_128
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1161 : std_logic;

begin
   
   n2 <= '0';
   add_16 : PC_adder_1_DW01_add_0_DW01_add_128 port map( A(31) => A(31), A(30) 
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => n2, SUM(31) => Sum(31),
                           SUM(30) => Sum(30), SUM(29) => Sum(29), SUM(28) => 
                           Sum(28), SUM(27) => Sum(27), SUM(26) => Sum(26), 
                           SUM(25) => Sum(25), SUM(24) => Sum(24), SUM(23) => 
                           Sum(23), SUM(22) => Sum(22), SUM(21) => Sum(21), 
                           SUM(20) => Sum(20), SUM(19) => Sum(19), SUM(18) => 
                           Sum(18), SUM(17) => Sum(17), SUM(16) => Sum(16), 
                           SUM(15) => Sum(15), SUM(14) => Sum(14), SUM(13) => 
                           Sum(13), SUM(12) => Sum(12), SUM(11) => Sum(11), 
                           SUM(10) => Sum(10), SUM(9) => Sum(9), SUM(8) => 
                           Sum(8), SUM(7) => Sum(7), SUM(6) => Sum(6), SUM(5) 
                           => Sum(5), SUM(4) => Sum(4), SUM(3) => Sum(3), 
                           SUM(2) => Sum(2), SUM(1) => Sum(1), SUM(0) => Sum(0)
                           , CO => n_1161);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FFD_1;

architecture SYN_BEHAVIORAL of FFD_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n3, n_1162 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFRS_X1 port map( D => n3, CK => CK, RN => n2, SN => n1, Q => 
                           Q_port, QN => n_1162);
   n1 <= '1';
   U3 : INV_X1 port map( A => RESET, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_17 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_17;

architecture SYN_Behavioral of REG_NBIT32_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_28_port, 
      data_out_27_port, data_out_26_port, data_out_25_port, data_out_24_port, 
      data_out_23_port, data_out_22_port, data_out_21_port, data_out_20_port, 
      data_out_19_port, data_out_18_port, data_out_17_port, data_out_16_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, data_out_0_port, data_out_1_port, 
      data_out_2_port, data_out_3_port, data_out_4_port, data_out_5_port, 
      data_out_6_port, data_out_7_port, data_out_8_port, data_out_9_port, 
      data_out_10_port, data_out_11_port, data_out_12_port, data_out_13_port, 
      data_out_14_port, data_out_15_port, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, data_out_29_port, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n55, n56, n57, n61, n62, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183 : 
      std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_31_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n5, Q => 
                           data_out_31_port, QN => n95);
   reg_reg_30_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n5, Q => 
                           data_out_30_port, QN => n96);
   reg_reg_29_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n5, Q => 
                           data_out_29_port, QN => n_1163);
   reg_reg_28_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n5, Q => 
                           data_out_28_port, QN => n_1164);
   reg_reg_27_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n5, Q => 
                           data_out_27_port, QN => n97);
   reg_reg_26_inst : DFFR_X1 port map( D => n42, CK => clk, RN => n5, Q => 
                           data_out_26_port, QN => n98);
   reg_reg_25_inst : DFFR_X1 port map( D => n43, CK => clk, RN => n5, Q => 
                           data_out_25_port, QN => n99);
   reg_reg_24_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n5, Q => 
                           data_out_24_port, QN => n_1165);
   reg_reg_23_inst : DFFR_X1 port map( D => n45, CK => clk, RN => n5, Q => 
                           data_out_23_port, QN => n_1166);
   reg_reg_22_inst : DFFR_X1 port map( D => n46, CK => clk, RN => n5, Q => 
                           data_out_22_port, QN => n_1167);
   reg_reg_21_inst : DFFR_X1 port map( D => n47, CK => clk, RN => n5, Q => 
                           data_out_21_port, QN => n100);
   reg_reg_20_inst : DFFR_X1 port map( D => n48, CK => clk, RN => n5, Q => 
                           data_out_20_port, QN => n101);
   reg_reg_19_inst : DFFR_X1 port map( D => n55, CK => clk, RN => n6, Q => 
                           data_out_19_port, QN => n102);
   reg_reg_18_inst : DFFR_X1 port map( D => n56, CK => clk, RN => n6, Q => 
                           data_out_18_port, QN => n103);
   reg_reg_17_inst : DFFR_X1 port map( D => n57, CK => clk, RN => n6, Q => 
                           data_out_17_port, QN => n104);
   reg_reg_16_inst : DFFR_X1 port map( D => n61, CK => clk, RN => n6, Q => 
                           data_out_16_port, QN => n105);
   reg_reg_15_inst : DFFR_X1 port map( D => n62, CK => clk, RN => n8, Q => 
                           data_out_15_port, QN => n_1168);
   reg_reg_14_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n8, Q => 
                           data_out_14_port, QN => n_1169);
   reg_reg_13_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n8, Q => 
                           data_out_13_port, QN => n_1170);
   reg_reg_12_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n8, Q => 
                           data_out_12_port, QN => n_1171);
   reg_reg_11_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n8, Q => 
                           data_out_11_port, QN => n_1172);
   reg_reg_10_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n8, Q => 
                           data_out_10_port, QN => n_1173);
   reg_reg_9_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n8, Q => 
                           data_out_9_port, QN => n_1174);
   reg_reg_8_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n8, Q => 
                           data_out_8_port, QN => n_1175);
   reg_reg_7_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n8, Q => 
                           data_out_7_port, QN => n_1176);
   reg_reg_6_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n8, Q => 
                           data_out_6_port, QN => n_1177);
   reg_reg_5_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n8, Q => 
                           data_out_5_port, QN => n_1178);
   reg_reg_4_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n8, Q => 
                           data_out_4_port, QN => n_1179);
   reg_reg_3_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n8, Q => 
                           data_out_3_port, QN => n_1180);
   reg_reg_2_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n8, Q => 
                           data_out_2_port, QN => n_1181);
   reg_reg_1_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n8, Q => 
                           data_out_1_port, QN => n_1182);
   reg_reg_0_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n8, Q => 
                           data_out_0_port, QN => n_1183);
   U2 : BUF_X1 port map( A => enable, Z => n4);
   U3 : BUF_X1 port map( A => n8, Z => n7);
   U4 : BUF_X1 port map( A => n4, Z => n3);
   U5 : BUF_X1 port map( A => n4, Z => n1);
   U6 : BUF_X1 port map( A => n4, Z => n2);
   U7 : BUF_X1 port map( A => n7, Z => n6);
   U8 : BUF_X1 port map( A => n7, Z => n5);
   U9 : INV_X1 port map( A => reset, ZN => n8);
   U10 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => n1, Z =>
                           n94);
   U11 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n1, Z =>
                           n93);
   U12 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => n1, Z =>
                           n92);
   U13 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => n1, Z =>
                           n91);
   U14 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => n1, Z =>
                           n90);
   U15 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n1, Z =>
                           n89);
   U16 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n1, Z =>
                           n88);
   U17 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => n1, Z =>
                           n87);
   U18 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => n1, Z =>
                           n86);
   U19 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n1, Z =>
                           n85);
   U20 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => n1, Z 
                           => n84);
   U21 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => n1, Z 
                           => n83);
   U22 : MUX2_X1 port map( A => data_out_12_port, B => data_in(12), S => n2, Z 
                           => n82);
   U23 : MUX2_X1 port map( A => data_out_13_port, B => data_in(13), S => n2, Z 
                           => n81);
   U24 : MUX2_X1 port map( A => data_out_14_port, B => data_in(14), S => n2, Z 
                           => n80);
   U25 : MUX2_X1 port map( A => data_out_15_port, B => data_in(15), S => n2, Z 
                           => n62);
   U26 : INV_X1 port map( A => n105, ZN => n25);
   U27 : MUX2_X1 port map( A => n25, B => data_in(16), S => n2, Z => n61);
   U28 : INV_X1 port map( A => n104, ZN => n26);
   U29 : MUX2_X1 port map( A => n26, B => data_in(17), S => n2, Z => n57);
   U30 : INV_X1 port map( A => n103, ZN => n27);
   U31 : MUX2_X1 port map( A => n27, B => data_in(18), S => n2, Z => n56);
   U32 : INV_X1 port map( A => n102, ZN => n28);
   U33 : MUX2_X1 port map( A => n28, B => data_in(19), S => n2, Z => n55);
   U34 : INV_X1 port map( A => n101, ZN => n29);
   U35 : MUX2_X1 port map( A => n29, B => data_in(20), S => n2, Z => n48);
   U36 : INV_X1 port map( A => n100, ZN => n30);
   U37 : MUX2_X1 port map( A => n30, B => data_in(21), S => n2, Z => n47);
   U38 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => n2, Z 
                           => n46);
   U39 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => n2, Z 
                           => n45);
   U40 : MUX2_X1 port map( A => data_out_24_port, B => data_in(24), S => n3, Z 
                           => n44);
   U41 : INV_X1 port map( A => n99, ZN => n31);
   U42 : MUX2_X1 port map( A => n31, B => data_in(25), S => n3, Z => n43);
   U43 : INV_X1 port map( A => n98, ZN => n32);
   U44 : MUX2_X1 port map( A => n32, B => data_in(26), S => n3, Z => n42);
   U45 : INV_X1 port map( A => n97, ZN => n33);
   U46 : MUX2_X1 port map( A => n33, B => data_in(27), S => n3, Z => n41);
   U47 : MUX2_X1 port map( A => data_out_28_port, B => data_in(28), S => n3, Z 
                           => n40);
   U48 : MUX2_X1 port map( A => data_out_29_port, B => data_in(29), S => n3, Z 
                           => n39);
   U49 : INV_X1 port map( A => n96, ZN => n35);
   U50 : MUX2_X1 port map( A => n35, B => data_in(30), S => n3, Z => n38);
   U51 : INV_X1 port map( A => n95, ZN => n36);
   U52 : MUX2_X1 port map( A => n36, B => data_in(31), S => n3, Z => n37);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_16 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_16;

architecture SYN_Behavioral of REG_NBIT32_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, data_out_0_port, data_out_1_port, data_out_2_port
      , data_out_3_port, data_out_4_port, data_out_5_port, data_out_6_port, 
      data_out_7_port, data_out_8_port, data_out_9_port, data_out_10_port, 
      data_out_11_port, data_out_12_port, data_out_13_port, data_out_14_port, 
      data_out_15_port, data_out_16_port, data_out_17_port, data_out_18_port, 
      data_out_19_port, data_out_20_port, data_out_21_port, data_out_22_port, 
      data_out_23_port, data_out_24_port, data_out_25_port, data_out_26_port, 
      data_out_27_port, data_out_28_port, data_out_29_port, data_out_30_port, 
      data_out_31_port, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n70, n71, n72, n73, n74, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215 : 
      std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_0_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n5, Q => 
                           data_out_0_port, QN => n_1184);
   reg_reg_1_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n5, Q => 
                           data_out_1_port, QN => n_1185);
   reg_reg_2_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n5, Q => 
                           data_out_2_port, QN => n_1186);
   reg_reg_3_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n5, Q => 
                           data_out_3_port, QN => n_1187);
   reg_reg_4_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n5, Q => 
                           data_out_4_port, QN => n_1188);
   reg_reg_5_inst : DFFR_X1 port map( D => n64, CK => clk, RN => n5, Q => 
                           data_out_5_port, QN => n_1189);
   reg_reg_8_inst : DFFR_X1 port map( D => n61, CK => clk, RN => n5, Q => 
                           data_out_8_port, QN => n_1190);
   reg_reg_9_inst : DFFR_X1 port map( D => n60, CK => clk, RN => n5, Q => 
                           data_out_9_port, QN => n_1191);
   reg_reg_12_inst : DFFR_X1 port map( D => n57, CK => clk, RN => n5, Q => 
                           data_out_12_port, QN => n_1192);
   reg_reg_6_inst : DFFR_X1 port map( D => n63, CK => clk, RN => n5, Q => 
                           data_out_6_port, QN => n_1193);
   reg_reg_13_inst : DFFR_X1 port map( D => n56, CK => clk, RN => n5, Q => 
                           data_out_13_port, QN => n_1194);
   reg_reg_16_inst : DFFR_X1 port map( D => n53, CK => clk, RN => n5, Q => 
                           data_out_16_port, QN => n_1195);
   reg_reg_10_inst : DFFR_X1 port map( D => n59, CK => clk, RN => n5, Q => 
                           data_out_10_port, QN => n_1196);
   reg_reg_11_inst : DFFR_X1 port map( D => n58, CK => clk, RN => n5, Q => 
                           data_out_11_port, QN => n_1197);
   reg_reg_7_inst : DFFR_X1 port map( D => n62, CK => clk, RN => n5, Q => 
                           data_out_7_port, QN => n_1198);
   reg_reg_14_inst : DFFR_X1 port map( D => n55, CK => clk, RN => n5, Q => 
                           data_out_14_port, QN => n_1199);
   reg_reg_15_inst : DFFR_X1 port map( D => n54, CK => clk, RN => n5, Q => 
                           data_out_15_port, QN => n_1200);
   reg_reg_21_inst : DFFR_X1 port map( D => n48, CK => clk, RN => n5, Q => 
                           data_out_21_port, QN => n_1201);
   reg_reg_24_inst : DFFR_X1 port map( D => n45, CK => clk, RN => n5, Q => 
                           data_out_24_port, QN => n_1202);
   reg_reg_28_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n5, Q => 
                           data_out_28_port, QN => n_1203);
   reg_reg_17_inst : DFFR_X1 port map( D => n52, CK => clk, RN => n5, Q => 
                           data_out_17_port, QN => n_1204);
   reg_reg_20_inst : DFFR_X1 port map( D => n49, CK => clk, RN => n5, Q => 
                           data_out_20_port, QN => n_1205);
   reg_reg_18_inst : DFFR_X1 port map( D => n51, CK => clk, RN => n5, Q => 
                           data_out_18_port, QN => n_1206);
   reg_reg_25_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n5, Q => 
                           data_out_25_port, QN => n_1207);
   reg_reg_26_inst : DFFR_X1 port map( D => n43, CK => clk, RN => n5, Q => 
                           data_out_26_port, QN => n_1208);
   reg_reg_29_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n5, Q => 
                           data_out_29_port, QN => n_1209);
   reg_reg_23_inst : DFFR_X1 port map( D => n46, CK => clk, RN => n5, Q => 
                           data_out_23_port, QN => n_1210);
   reg_reg_27_inst : DFFR_X1 port map( D => n42, CK => clk, RN => n5, Q => 
                           data_out_27_port, QN => n_1211);
   reg_reg_31_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n5, Q => 
                           data_out_31_port, QN => n_1212);
   reg_reg_22_inst : DFFR_X1 port map( D => n47, CK => clk, RN => n5, Q => 
                           data_out_22_port, QN => n_1213);
   reg_reg_19_inst : DFFR_X1 port map( D => n50, CK => clk, RN => n5, Q => 
                           data_out_19_port, QN => n_1214);
   reg_reg_30_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n5, Q => 
                           data_out_30_port, QN => n_1215);
   U2 : INV_X2 port map( A => reset, ZN => n5);
   U3 : BUF_X1 port map( A => enable, Z => n4);
   U4 : BUF_X1 port map( A => n4, Z => n3);
   U5 : BUF_X1 port map( A => n4, Z => n1);
   U6 : BUF_X1 port map( A => n4, Z => n2);
   U7 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => n1, Z => 
                           n74);
   U8 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n1, Z => 
                           n73);
   U9 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => n1, Z => 
                           n72);
   U10 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => n1, Z =>
                           n71);
   U11 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => n1, Z =>
                           n70);
   U12 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n1, Z =>
                           n64);
   U13 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n1, Z =>
                           n63);
   U14 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => n1, Z =>
                           n62);
   U15 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => n1, Z =>
                           n61);
   U16 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n1, Z =>
                           n60);
   U17 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => n1, Z 
                           => n59);
   U18 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => n1, Z 
                           => n58);
   U19 : MUX2_X1 port map( A => data_out_12_port, B => data_in(12), S => n2, Z 
                           => n57);
   U20 : MUX2_X1 port map( A => data_out_13_port, B => data_in(13), S => n2, Z 
                           => n56);
   U21 : MUX2_X1 port map( A => data_out_14_port, B => data_in(14), S => n2, Z 
                           => n55);
   U22 : MUX2_X1 port map( A => data_out_15_port, B => data_in(15), S => n2, Z 
                           => n54);
   U23 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => n2, Z 
                           => n53);
   U24 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => n2, Z 
                           => n52);
   U25 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => n2, Z 
                           => n51);
   U26 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => n2, Z 
                           => n50);
   U27 : MUX2_X1 port map( A => data_out_20_port, B => data_in(20), S => n2, Z 
                           => n49);
   U28 : MUX2_X1 port map( A => data_out_21_port, B => data_in(21), S => n2, Z 
                           => n48);
   U29 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => n2, Z 
                           => n47);
   U30 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => n2, Z 
                           => n46);
   U31 : MUX2_X1 port map( A => data_out_24_port, B => data_in(24), S => n3, Z 
                           => n45);
   U32 : MUX2_X1 port map( A => data_out_25_port, B => data_in(25), S => n3, Z 
                           => n44);
   U33 : MUX2_X1 port map( A => data_out_26_port, B => data_in(26), S => n3, Z 
                           => n43);
   U34 : MUX2_X1 port map( A => data_out_27_port, B => data_in(27), S => n3, Z 
                           => n42);
   U35 : MUX2_X1 port map( A => data_out_28_port, B => data_in(28), S => n3, Z 
                           => n41);
   U36 : MUX2_X1 port map( A => data_out_29_port, B => data_in(29), S => n3, Z 
                           => n40);
   U37 : MUX2_X1 port map( A => data_out_30_port, B => data_in(30), S => n3, Z 
                           => n39);
   U38 : MUX2_X1 port map( A => data_out_31_port, B => data_in(31), S => n3, Z 
                           => n38);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_15 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_15;

architecture SYN_Behavioral of REG_NBIT32_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202 : 
      std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n102, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n102, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n102, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n102, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n102, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n102, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n102, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n102, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n102, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n102, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n102, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n102, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n103, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n103, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n103, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n103, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n103, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n103, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n103, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n103, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n103, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n103, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n103, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n103, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n104, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n104, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n104, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n104, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n104, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n104, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n104, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n104, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n1, Z => n100);
   U3 : BUF_X1 port map( A => n106, Z => n105);
   U4 : BUF_X1 port map( A => n101, Z => n3);
   U5 : BUF_X1 port map( A => n101, Z => n2);
   U6 : BUF_X1 port map( A => n100, Z => n96);
   U7 : BUF_X1 port map( A => n100, Z => n98);
   U8 : BUF_X1 port map( A => n100, Z => n99);
   U9 : BUF_X1 port map( A => n105, Z => n103);
   U10 : BUF_X1 port map( A => n105, Z => n102);
   U11 : BUF_X1 port map( A => n105, Z => n104);
   U12 : INV_X1 port map( A => reset, ZN => n106);
   U13 : BUF_X1 port map( A => n1, Z => n101);
   U14 : BUF_X1 port map( A => enable, Z => n1);
   U15 : OAI21_X1 port map( B1 => n170, B2 => n99, A => n202, ZN => n138);
   U16 : NAND2_X1 port map( A1 => data_in(3), A2 => n2, ZN => n202);
   U17 : OAI21_X1 port map( B1 => n169, B2 => n99, A => n201, ZN => n137);
   U18 : NAND2_X1 port map( A1 => data_in(4), A2 => n2, ZN => n201);
   U19 : OAI21_X1 port map( B1 => n168, B2 => n98, A => n200, ZN => n136);
   U20 : NAND2_X1 port map( A1 => data_in(5), A2 => n2, ZN => n200);
   U21 : OAI21_X1 port map( B1 => n167, B2 => n99, A => n199, ZN => n135);
   U22 : NAND2_X1 port map( A1 => data_in(6), A2 => n2, ZN => n199);
   U23 : OAI21_X1 port map( B1 => n166, B2 => n99, A => n198, ZN => n134);
   U24 : NAND2_X1 port map( A1 => data_in(7), A2 => n2, ZN => n198);
   U25 : OAI21_X1 port map( B1 => n165, B2 => n99, A => n197, ZN => n133);
   U26 : NAND2_X1 port map( A1 => data_in(8), A2 => n2, ZN => n197);
   U27 : OAI21_X1 port map( B1 => n164, B2 => n99, A => n196, ZN => n132);
   U28 : NAND2_X1 port map( A1 => data_in(9), A2 => n3, ZN => n196);
   U29 : OAI21_X1 port map( B1 => n163, B2 => n99, A => n195, ZN => n131);
   U30 : NAND2_X1 port map( A1 => data_in(10), A2 => n3, ZN => n195);
   U31 : OAI21_X1 port map( B1 => n162, B2 => n99, A => n194, ZN => n130);
   U32 : NAND2_X1 port map( A1 => data_in(11), A2 => n2, ZN => n194);
   U33 : OAI21_X1 port map( B1 => n161, B2 => n99, A => n193, ZN => n129);
   U34 : NAND2_X1 port map( A1 => data_in(12), A2 => n3, ZN => n193);
   U35 : OAI21_X1 port map( B1 => n160, B2 => n99, A => n192, ZN => n128);
   U36 : NAND2_X1 port map( A1 => data_in(13), A2 => n3, ZN => n192);
   U37 : OAI21_X1 port map( B1 => n159, B2 => n98, A => n191, ZN => n127);
   U38 : NAND2_X1 port map( A1 => data_in(14), A2 => n3, ZN => n191);
   U39 : OAI21_X1 port map( B1 => n158, B2 => n98, A => n190, ZN => n126);
   U40 : NAND2_X1 port map( A1 => data_in(15), A2 => n3, ZN => n190);
   U41 : OAI21_X1 port map( B1 => n157, B2 => n98, A => n189, ZN => n125);
   U42 : NAND2_X1 port map( A1 => data_in(16), A2 => n3, ZN => n189);
   U43 : OAI21_X1 port map( B1 => n156, B2 => n98, A => n188, ZN => n124);
   U44 : NAND2_X1 port map( A1 => data_in(17), A2 => n3, ZN => n188);
   U45 : OAI21_X1 port map( B1 => n155, B2 => n98, A => n187, ZN => n123);
   U46 : NAND2_X1 port map( A1 => data_in(18), A2 => n96, ZN => n187);
   U47 : OAI21_X1 port map( B1 => n154, B2 => n98, A => n186, ZN => n122);
   U48 : NAND2_X1 port map( A1 => data_in(19), A2 => n96, ZN => n186);
   U49 : OAI21_X1 port map( B1 => n153, B2 => n98, A => n185, ZN => n121);
   U50 : NAND2_X1 port map( A1 => data_in(20), A2 => n96, ZN => n185);
   U51 : OAI21_X1 port map( B1 => n152, B2 => n98, A => n184, ZN => n120);
   U52 : NAND2_X1 port map( A1 => data_in(21), A2 => n96, ZN => n184);
   U53 : OAI21_X1 port map( B1 => n151, B2 => n98, A => n183, ZN => n119);
   U54 : NAND2_X1 port map( A1 => data_in(22), A2 => n96, ZN => n183);
   U55 : OAI21_X1 port map( B1 => n150, B2 => n98, A => n182, ZN => n118);
   U56 : NAND2_X1 port map( A1 => data_in(23), A2 => n3, ZN => n182);
   U57 : OAI21_X1 port map( B1 => n149, B2 => n96, A => n181, ZN => n117);
   U58 : NAND2_X1 port map( A1 => data_in(24), A2 => n3, ZN => n181);
   U59 : OAI21_X1 port map( B1 => n148, B2 => n98, A => n180, ZN => n116);
   U60 : NAND2_X1 port map( A1 => data_in(25), A2 => n3, ZN => n180);
   U61 : OAI21_X1 port map( B1 => n147, B2 => n96, A => n179, ZN => n115);
   U62 : NAND2_X1 port map( A1 => data_in(26), A2 => n2, ZN => n179);
   U63 : OAI21_X1 port map( B1 => n146, B2 => n96, A => n178, ZN => n114);
   U64 : NAND2_X1 port map( A1 => data_in(27), A2 => n3, ZN => n178);
   U65 : OAI21_X1 port map( B1 => n145, B2 => n96, A => n177, ZN => n113);
   U66 : NAND2_X1 port map( A1 => data_in(28), A2 => n2, ZN => n177);
   U67 : OAI21_X1 port map( B1 => n144, B2 => n96, A => n176, ZN => n112);
   U68 : NAND2_X1 port map( A1 => data_in(29), A2 => n2, ZN => n176);
   U69 : OAI21_X1 port map( B1 => n143, B2 => n96, A => n175, ZN => n111);
   U70 : NAND2_X1 port map( A1 => data_in(30), A2 => n2, ZN => n175);
   U71 : OAI21_X1 port map( B1 => n142, B2 => n96, A => n174, ZN => n110);
   U72 : NAND2_X1 port map( A1 => data_in(31), A2 => n2, ZN => n174);
   U73 : INV_X1 port map( A => n173, ZN => n107);
   U74 : MUX2_X1 port map( A => n107, B => data_in(0), S => n99, Z => n141);
   U75 : INV_X1 port map( A => n172, ZN => n108);
   U76 : MUX2_X1 port map( A => n108, B => data_in(1), S => n99, Z => n140);
   U77 : INV_X1 port map( A => n171, ZN => n109);
   U78 : MUX2_X1 port map( A => n109, B => data_in(2), S => n99, Z => n139);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_14 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_14;

architecture SYN_Behavioral of REG_NBIT32_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n_1216
      , n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225,
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_31_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n5, Q => 
                           data_out_31_port, QN => n_1216);
   reg_reg_30_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n5, Q => 
                           data_out_30_port, QN => n_1217);
   reg_reg_29_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n5, Q => 
                           data_out_29_port, QN => n_1218);
   reg_reg_28_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n5, Q => 
                           data_out_28_port, QN => n_1219);
   reg_reg_27_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n5, Q => 
                           data_out_27_port, QN => n_1220);
   reg_reg_26_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n5, Q => 
                           data_out_26_port, QN => n_1221);
   reg_reg_25_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n5, Q => 
                           data_out_25_port, QN => n_1222);
   reg_reg_24_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n5, Q => 
                           data_out_24_port, QN => n_1223);
   reg_reg_23_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n5, Q => 
                           data_out_23_port, QN => n_1224);
   reg_reg_22_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n5, Q => 
                           data_out_22_port, QN => n_1225);
   reg_reg_21_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n5, Q => 
                           data_out_21_port, QN => n_1226);
   reg_reg_20_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n5, Q => 
                           data_out_20_port, QN => n_1227);
   reg_reg_19_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n6, Q => 
                           data_out_19_port, QN => n_1228);
   reg_reg_18_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n6, Q => 
                           data_out_18_port, QN => n_1229);
   reg_reg_17_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n6, Q => 
                           data_out_17_port, QN => n_1230);
   reg_reg_16_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n6, Q => 
                           data_out_16_port, QN => n_1231);
   reg_reg_15_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n6, Q => 
                           data_out_15_port, QN => n_1232);
   reg_reg_14_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n6, Q => 
                           data_out_14_port, QN => n_1233);
   reg_reg_13_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n6, Q => 
                           data_out_13_port, QN => n_1234);
   reg_reg_12_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n6, Q => 
                           data_out_12_port, QN => n_1235);
   reg_reg_11_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n6, Q => 
                           data_out_11_port, QN => n_1236);
   reg_reg_10_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n6, Q => 
                           data_out_10_port, QN => n_1237);
   reg_reg_9_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n6, Q => 
                           data_out_9_port, QN => n_1238);
   reg_reg_8_inst : DFFR_X1 port map( D => n33, CK => clk, RN => n6, Q => 
                           data_out_8_port, QN => n_1239);
   reg_reg_7_inst : DFFR_X1 port map( D => n34, CK => clk, RN => n7, Q => 
                           data_out_7_port, QN => n_1240);
   reg_reg_6_inst : DFFR_X1 port map( D => n35, CK => clk, RN => n7, Q => 
                           data_out_6_port, QN => n_1241);
   reg_reg_5_inst : DFFR_X1 port map( D => n36, CK => clk, RN => n7, Q => 
                           data_out_5_port, QN => n_1242);
   reg_reg_4_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n7, Q => 
                           data_out_4_port, QN => n_1243);
   reg_reg_3_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n7, Q => 
                           data_out_3_port, QN => n_1244);
   reg_reg_2_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n7, Q => 
                           data_out_2_port, QN => n_1245);
   reg_reg_1_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n7, Q => 
                           data_out_1_port, QN => n_1246);
   reg_reg_0_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n7, Q => 
                           data_out_0_port, QN => n_1247);
   U2 : BUF_X1 port map( A => n9, Z => n8);
   U3 : BUF_X1 port map( A => enable, Z => n4);
   U4 : BUF_X1 port map( A => n8, Z => n6);
   U5 : BUF_X1 port map( A => n8, Z => n5);
   U6 : BUF_X1 port map( A => n8, Z => n7);
   U7 : INV_X1 port map( A => reset, ZN => n9);
   U8 : BUF_X1 port map( A => n4, Z => n1);
   U9 : BUF_X1 port map( A => n4, Z => n2);
   U10 : BUF_X1 port map( A => n4, Z => n3);
   U11 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => n1, Z =>
                           n41);
   U12 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n1, Z =>
                           n40);
   U13 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => n1, Z =>
                           n39);
   U14 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => n1, Z =>
                           n38);
   U15 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => n1, Z =>
                           n37);
   U16 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n1, Z =>
                           n36);
   U17 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n1, Z =>
                           n35);
   U18 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => n1, Z =>
                           n34);
   U19 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => n1, Z =>
                           n33);
   U20 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n1, Z =>
                           n32);
   U21 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => n1, Z 
                           => n31);
   U22 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => n1, Z 
                           => n30);
   U23 : MUX2_X1 port map( A => data_out_12_port, B => data_in(12), S => n2, Z 
                           => n29);
   U24 : MUX2_X1 port map( A => data_out_13_port, B => data_in(13), S => n2, Z 
                           => n28);
   U25 : MUX2_X1 port map( A => data_out_14_port, B => data_in(14), S => n2, Z 
                           => n27);
   U26 : MUX2_X1 port map( A => data_out_15_port, B => data_in(15), S => n2, Z 
                           => n26);
   U27 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => n2, Z 
                           => n25);
   U28 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => n2, Z 
                           => n24);
   U29 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => n2, Z 
                           => n23);
   U30 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => n2, Z 
                           => n22);
   U31 : MUX2_X1 port map( A => data_out_20_port, B => data_in(20), S => n2, Z 
                           => n21);
   U32 : MUX2_X1 port map( A => data_out_21_port, B => data_in(21), S => n2, Z 
                           => n20);
   U33 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => n2, Z 
                           => n19);
   U34 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => n2, Z 
                           => n18);
   U35 : MUX2_X1 port map( A => data_out_24_port, B => data_in(24), S => n3, Z 
                           => n17);
   U36 : MUX2_X1 port map( A => data_out_25_port, B => data_in(25), S => n3, Z 
                           => n16);
   U37 : MUX2_X1 port map( A => data_out_26_port, B => data_in(26), S => n3, Z 
                           => n15);
   U38 : MUX2_X1 port map( A => data_out_27_port, B => data_in(27), S => n3, Z 
                           => n14);
   U39 : MUX2_X1 port map( A => data_out_28_port, B => data_in(28), S => n3, Z 
                           => n13);
   U40 : MUX2_X1 port map( A => data_out_29_port, B => data_in(29), S => n3, Z 
                           => n12);
   U41 : MUX2_X1 port map( A => data_out_30_port, B => data_in(30), S => n3, Z 
                           => n11);
   U42 : MUX2_X1 port map( A => data_out_31_port, B => data_in(31), S => n3, Z 
                           => n10);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_13 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_13;

architecture SYN_Behavioral of REG_NBIT32_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n27, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n105, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n105, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n105, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n105, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n105, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n107, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n105, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n105, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n105, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n105, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n105, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n105, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n105, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n106, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n106, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n106, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n106, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n106, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n106, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n106, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n107, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n107, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n107, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n107, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n107, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n107, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n107, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n27, Z => n104);
   U3 : BUF_X1 port map( A => n27, Z => n103);
   U4 : BUF_X1 port map( A => n104, Z => n98);
   U5 : BUF_X1 port map( A => n104, Z => n96);
   U6 : BUF_X1 port map( A => n104, Z => n99);
   U7 : BUF_X1 port map( A => n103, Z => n100);
   U8 : BUF_X1 port map( A => n103, Z => n101);
   U9 : BUF_X1 port map( A => n108, Z => n106);
   U10 : BUF_X1 port map( A => n108, Z => n105);
   U11 : BUF_X1 port map( A => n108, Z => n107);
   U12 : BUF_X1 port map( A => n103, Z => n102);
   U13 : INV_X1 port map( A => reset, ZN => n108);
   U14 : BUF_X1 port map( A => enable, Z => n27);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n101, A => n204, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n102, A2 => data_in(0), ZN => n204);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n101, A => n203, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n99, ZN => n203);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n101, A => n202, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n99, ZN => n202);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n101, A => n201, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n99, ZN => n201);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n101, A => n200, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n99, ZN => n200);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n100, A => n199, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n98, ZN => n199);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n100, A => n198, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n99, ZN => n198);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n197, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n197);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n99, A => n196, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n98, ZN => n196);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n99, A => n195, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n98, ZN => n195);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n99, A => n194, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n98, ZN => n194);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n193, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n98, ZN => n193);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n99, A => n192, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n98, ZN => n192);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n99, A => n191, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n98, ZN => n191);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n190, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n98, ZN => n190);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n99, A => n189, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n98, ZN => n189);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n100, A => n188, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n98, ZN => n188);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n100, A => n187, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n98, ZN => n187);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n100, A => n186, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n98, ZN => n186);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n100, A => n185, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n96, ZN => n185);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n100, A => n184, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n96, ZN => n184);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n100, A => n183, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n96, ZN => n183);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n100, A => n182, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n96, ZN => n182);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n101, A => n181, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n96, ZN => n181);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n101, A => n180, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n96, ZN => n180);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n101, A => n179, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n96, ZN => n179);
   U67 : OAI21_X1 port map( B1 => n146, B2 => n101, A => n178, ZN => n114);
   U68 : NAND2_X1 port map( A1 => data_in(27), A2 => n96, ZN => n178);
   U69 : OAI21_X1 port map( B1 => n145, B2 => n101, A => n177, ZN => n113);
   U70 : NAND2_X1 port map( A1 => data_in(28), A2 => n96, ZN => n177);
   U71 : OAI21_X1 port map( B1 => n144, B2 => n101, A => n176, ZN => n112);
   U72 : NAND2_X1 port map( A1 => data_in(29), A2 => n96, ZN => n176);
   U73 : OAI21_X1 port map( B1 => n143, B2 => n101, A => n175, ZN => n111);
   U74 : NAND2_X1 port map( A1 => data_in(30), A2 => n96, ZN => n175);
   U75 : OAI21_X1 port map( B1 => n142, B2 => n102, A => n174, ZN => n110);
   U76 : NAND2_X1 port map( A1 => data_in(31), A2 => n96, ZN => n174);
   U77 : INV_X1 port map( A => n147, ZN => n109);
   U78 : MUX2_X1 port map( A => n109, B => data_in(26), S => n102, Z => n115);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_12 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_12;

architecture SYN_Behavioral of REG_NBIT32_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_8_port, 
      data_out_7_port, data_out_6_port, data_out_4_port, data_out_3_port, 
      data_out_2_port, data_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10
      , data_out_1_port, n12, n13, n14, data_out_5_port, n16, n17, n18, 
      data_out_9_port, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n34, 
      n38, n42, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n_1248,
      n_1249, n_1250 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_31_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n5, Q => 
                           data_out_31_port, QN => n135);
   reg_reg_28_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n5, Q => 
                           data_out_28_port, QN => n138);
   reg_reg_27_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n5, Q => 
                           data_out_27_port, QN => n139);
   reg_reg_26_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n5, Q => 
                           data_out_26_port, QN => n140);
   reg_reg_25_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n5, Q => 
                           data_out_25_port, QN => n141);
   reg_reg_24_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n5, Q => 
                           data_out_24_port, QN => n142);
   reg_reg_23_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n5, Q => 
                           data_out_23_port, QN => n143);
   reg_reg_22_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n5, Q => 
                           data_out_22_port, QN => n144);
   reg_reg_21_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n5, Q => 
                           data_out_21_port, QN => n145);
   reg_reg_20_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n5, Q => 
                           data_out_20_port, QN => n146);
   reg_reg_19_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n6, Q => 
                           data_out_19_port, QN => n147);
   reg_reg_18_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n6, Q => 
                           data_out_18_port, QN => n148);
   reg_reg_17_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n6, Q => 
                           data_out_17_port, QN => n149);
   reg_reg_16_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n6, Q => 
                           data_out_16_port, QN => n150);
   reg_reg_15_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n6, Q => 
                           data_out_15_port, QN => n151);
   reg_reg_14_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n6, Q => 
                           data_out_14_port, QN => n152);
   reg_reg_13_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n6, Q => 
                           data_out_13_port, QN => n153);
   reg_reg_12_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n6, Q => 
                           data_out_12_port, QN => n154);
   reg_reg_11_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n6, Q => 
                           data_out_11_port, QN => n155);
   reg_reg_10_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n6, Q => 
                           data_out_10_port, QN => n156);
   reg_reg_9_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n6, Q => 
                           data_out_9_port, QN => n_1248);
   reg_reg_8_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n6, Q => 
                           data_out_8_port, QN => n157);
   reg_reg_7_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n7, Q => 
                           data_out_7_port, QN => n158);
   reg_reg_6_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n7, Q => 
                           data_out_6_port, QN => n159);
   reg_reg_4_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n7, Q => 
                           data_out_4_port, QN => n160);
   reg_reg_3_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n7, Q => 
                           data_out_3_port, QN => n161);
   reg_reg_2_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n7, Q => 
                           data_out_2_port, QN => n162);
   reg_reg_1_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n7, Q => 
                           data_out_1_port, QN => n_1249);
   reg_reg_0_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n7, Q => 
                           data_out_0_port, QN => n163);
   reg_reg_30_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n9, Q => 
                           data_out_30_port, QN => n136);
   reg_reg_29_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n9, Q => 
                           data_out_29_port, QN => n137);
   reg_reg_5_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n9, Q => 
                           data_out_5_port, QN => n_1250);
   U2 : BUF_X1 port map( A => n9, Z => n8);
   U3 : BUF_X1 port map( A => enable, Z => n4);
   U4 : BUF_X1 port map( A => n8, Z => n6);
   U5 : BUF_X1 port map( A => n8, Z => n5);
   U6 : BUF_X1 port map( A => n8, Z => n7);
   U7 : INV_X1 port map( A => reset, ZN => n9);
   U8 : BUF_X1 port map( A => n4, Z => n1);
   U9 : BUF_X1 port map( A => n4, Z => n2);
   U10 : BUF_X1 port map( A => n4, Z => n3);
   U11 : OAI21_X1 port map( B1 => n137, B2 => n1, A => n166, ZN => n105);
   U12 : NAND2_X1 port map( A1 => data_in(29), A2 => n1, ZN => n166);
   U13 : OAI21_X1 port map( B1 => n136, B2 => n1, A => n165, ZN => n104);
   U14 : NAND2_X1 port map( A1 => data_in(30), A2 => n1, ZN => n165);
   U15 : OAI21_X1 port map( B1 => n135, B2 => n1, A => n164, ZN => n103);
   U16 : NAND2_X1 port map( A1 => data_in(31), A2 => n1, ZN => n164);
   U17 : INV_X1 port map( A => n163, ZN => n10);
   U18 : MUX2_X1 port map( A => n10, B => data_in(0), S => n2, Z => n134);
   U19 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n1, Z =>
                           n133);
   U20 : INV_X1 port map( A => n162, ZN => n12);
   U21 : MUX2_X1 port map( A => n12, B => data_in(2), S => n3, Z => n132);
   U22 : INV_X1 port map( A => n161, ZN => n13);
   U23 : MUX2_X1 port map( A => n13, B => data_in(3), S => n3, Z => n131);
   U24 : INV_X1 port map( A => n160, ZN => n14);
   U25 : MUX2_X1 port map( A => n14, B => data_in(4), S => n2, Z => n130);
   U26 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n2, Z =>
                           n129);
   U27 : INV_X1 port map( A => n159, ZN => n16);
   U28 : MUX2_X1 port map( A => n16, B => data_in(6), S => n2, Z => n128);
   U29 : INV_X1 port map( A => n158, ZN => n17);
   U30 : MUX2_X1 port map( A => n17, B => data_in(7), S => n2, Z => n127);
   U31 : INV_X1 port map( A => n157, ZN => n18);
   U32 : MUX2_X1 port map( A => n18, B => data_in(8), S => n2, Z => n126);
   U33 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n2, Z =>
                           n125);
   U34 : INV_X1 port map( A => n156, ZN => n20);
   U35 : MUX2_X1 port map( A => n20, B => data_in(10), S => n2, Z => n124);
   U36 : INV_X1 port map( A => n155, ZN => n21);
   U37 : MUX2_X1 port map( A => n21, B => data_in(11), S => n2, Z => n123);
   U38 : INV_X1 port map( A => n154, ZN => n22);
   U39 : MUX2_X1 port map( A => n22, B => data_in(12), S => n2, Z => n122);
   U40 : INV_X1 port map( A => n153, ZN => n23);
   U41 : MUX2_X1 port map( A => n23, B => data_in(13), S => n2, Z => n121);
   U42 : INV_X1 port map( A => n152, ZN => n24);
   U43 : MUX2_X1 port map( A => n24, B => data_in(14), S => n2, Z => n120);
   U44 : INV_X1 port map( A => n151, ZN => n25);
   U45 : MUX2_X1 port map( A => n25, B => data_in(15), S => n2, Z => n119);
   U46 : INV_X1 port map( A => n150, ZN => n26);
   U47 : MUX2_X1 port map( A => n26, B => data_in(16), S => n2, Z => n118);
   U48 : INV_X1 port map( A => n149, ZN => n27);
   U49 : MUX2_X1 port map( A => n27, B => data_in(17), S => n2, Z => n117);
   U50 : INV_X1 port map( A => n148, ZN => n28);
   U51 : MUX2_X1 port map( A => n28, B => data_in(18), S => n2, Z => n116);
   U52 : INV_X1 port map( A => n147, ZN => n29);
   U53 : MUX2_X1 port map( A => n29, B => data_in(19), S => n2, Z => n115);
   U54 : INV_X1 port map( A => n146, ZN => n34);
   U55 : MUX2_X1 port map( A => n34, B => data_in(20), S => n2, Z => n114);
   U56 : INV_X1 port map( A => n145, ZN => n38);
   U57 : MUX2_X1 port map( A => n38, B => data_in(21), S => n1, Z => n113);
   U58 : INV_X1 port map( A => n144, ZN => n42);
   U59 : MUX2_X1 port map( A => n42, B => data_in(22), S => n1, Z => n112);
   U60 : INV_X1 port map( A => n143, ZN => n96);
   U61 : MUX2_X1 port map( A => n96, B => data_in(23), S => n1, Z => n111);
   U62 : INV_X1 port map( A => n142, ZN => n98);
   U63 : MUX2_X1 port map( A => n98, B => data_in(24), S => n1, Z => n110);
   U64 : INV_X1 port map( A => n141, ZN => n99);
   U65 : MUX2_X1 port map( A => n99, B => data_in(25), S => n1, Z => n109);
   U66 : INV_X1 port map( A => n140, ZN => n100);
   U67 : MUX2_X1 port map( A => n100, B => data_in(26), S => n1, Z => n108);
   U68 : INV_X1 port map( A => n139, ZN => n101);
   U69 : MUX2_X1 port map( A => n101, B => data_in(27), S => n1, Z => n107);
   U70 : INV_X1 port map( A => n138, ZN => n102);
   U71 : MUX2_X1 port map( A => n102, B => data_in(28), S => n1, Z => n106);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_11 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_11;

architecture SYN_Behavioral of REG_NBIT32_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n107, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n107, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n105, Z => n98);
   U5 : BUF_X1 port map( A => n105, Z => n99);
   U6 : BUF_X1 port map( A => n105, Z => n100);
   U7 : BUF_X1 port map( A => n104, Z => n101);
   U8 : BUF_X1 port map( A => n104, Z => n102);
   U9 : BUF_X1 port map( A => n109, Z => n106);
   U10 : BUF_X1 port map( A => n109, Z => n107);
   U11 : BUF_X1 port map( A => n109, Z => n108);
   U12 : BUF_X1 port map( A => n104, Z => n103);
   U13 : INV_X1 port map( A => reset, ZN => n109);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_10 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_10;

architecture SYN_Behavioral of REG_NBIT32_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201 : 
      std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n102, Q => 
                           data_out(31), QN => n141);
   reg_reg_30_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n102, Q => 
                           data_out(30), QN => n142);
   reg_reg_29_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n102, Q => 
                           data_out(29), QN => n143);
   reg_reg_28_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n102, Q => 
                           data_out(28), QN => n144);
   reg_reg_27_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n102, Q => 
                           data_out(27), QN => n145);
   reg_reg_26_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n102, Q => 
                           data_out(26), QN => n146);
   reg_reg_25_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n102, Q => 
                           data_out(25), QN => n147);
   reg_reg_24_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n102, Q => 
                           data_out(24), QN => n148);
   reg_reg_23_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n102, Q => 
                           data_out(23), QN => n149);
   reg_reg_22_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n102, Q => 
                           data_out(22), QN => n150);
   reg_reg_21_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n102, Q => 
                           data_out(21), QN => n151);
   reg_reg_20_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n102, Q => 
                           data_out(20), QN => n152);
   reg_reg_19_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n103, Q => 
                           data_out(19), QN => n153);
   reg_reg_18_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n103, Q => 
                           data_out(18), QN => n154);
   reg_reg_17_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n103, Q => 
                           data_out(17), QN => n155);
   reg_reg_16_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n103, Q => 
                           data_out(16), QN => n156);
   reg_reg_15_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n103, Q => 
                           data_out(15), QN => n157);
   reg_reg_14_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n103, Q => 
                           data_out(14), QN => n158);
   reg_reg_13_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n103, Q => 
                           data_out(13), QN => n159);
   reg_reg_12_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n103, Q => 
                           data_out(12), QN => n160);
   reg_reg_11_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n103, Q => 
                           data_out(11), QN => n161);
   reg_reg_10_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n103, Q => 
                           data_out(10), QN => n162);
   reg_reg_9_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n103, Q => 
                           data_out(9), QN => n163);
   reg_reg_8_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n103, Q => 
                           data_out(8), QN => n164);
   reg_reg_7_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n104, Q => 
                           data_out(7), QN => n165);
   reg_reg_6_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n104, Q => 
                           data_out(6), QN => n166);
   reg_reg_5_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n104, Q => 
                           data_out(5), QN => n167);
   reg_reg_4_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n104, Q => 
                           data_out(4), QN => n168);
   reg_reg_3_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n104, Q => 
                           data_out(3), QN => n169);
   reg_reg_2_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n104, Q => 
                           data_out(2), QN => n170);
   reg_reg_1_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n104, Q => 
                           data_out(1), QN => n171);
   reg_reg_0_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n104, Q => 
                           data_out(0), QN => n172);
   U2 : BUF_X1 port map( A => n1, Z => n100);
   U3 : BUF_X1 port map( A => n101, Z => n3);
   U4 : BUF_X1 port map( A => n101, Z => n2);
   U5 : BUF_X1 port map( A => n100, Z => n96);
   U6 : BUF_X1 port map( A => n100, Z => n98);
   U7 : BUF_X1 port map( A => n100, Z => n99);
   U8 : BUF_X1 port map( A => n105, Z => n103);
   U9 : BUF_X1 port map( A => n105, Z => n102);
   U10 : BUF_X1 port map( A => n105, Z => n104);
   U11 : INV_X1 port map( A => reset, ZN => n105);
   U12 : BUF_X1 port map( A => n1, Z => n101);
   U13 : BUF_X1 port map( A => enable, Z => n1);
   U14 : OAI21_X1 port map( B1 => n169, B2 => n99, A => n201, ZN => n137);
   U15 : NAND2_X1 port map( A1 => data_in(3), A2 => n2, ZN => n201);
   U16 : OAI21_X1 port map( B1 => n168, B2 => n99, A => n200, ZN => n136);
   U17 : NAND2_X1 port map( A1 => data_in(4), A2 => n2, ZN => n200);
   U18 : OAI21_X1 port map( B1 => n167, B2 => n98, A => n199, ZN => n135);
   U19 : NAND2_X1 port map( A1 => data_in(5), A2 => n2, ZN => n199);
   U20 : OAI21_X1 port map( B1 => n166, B2 => n99, A => n198, ZN => n134);
   U21 : NAND2_X1 port map( A1 => data_in(6), A2 => n2, ZN => n198);
   U22 : OAI21_X1 port map( B1 => n165, B2 => n99, A => n197, ZN => n133);
   U23 : NAND2_X1 port map( A1 => data_in(7), A2 => n2, ZN => n197);
   U24 : OAI21_X1 port map( B1 => n164, B2 => n99, A => n196, ZN => n132);
   U25 : NAND2_X1 port map( A1 => data_in(8), A2 => n2, ZN => n196);
   U26 : OAI21_X1 port map( B1 => n163, B2 => n99, A => n195, ZN => n131);
   U27 : NAND2_X1 port map( A1 => data_in(9), A2 => n3, ZN => n195);
   U28 : OAI21_X1 port map( B1 => n162, B2 => n99, A => n194, ZN => n130);
   U29 : NAND2_X1 port map( A1 => data_in(10), A2 => n3, ZN => n194);
   U30 : OAI21_X1 port map( B1 => n161, B2 => n99, A => n193, ZN => n129);
   U31 : NAND2_X1 port map( A1 => data_in(11), A2 => n2, ZN => n193);
   U32 : OAI21_X1 port map( B1 => n160, B2 => n99, A => n192, ZN => n128);
   U33 : NAND2_X1 port map( A1 => data_in(12), A2 => n3, ZN => n192);
   U34 : OAI21_X1 port map( B1 => n159, B2 => n99, A => n191, ZN => n127);
   U35 : NAND2_X1 port map( A1 => data_in(13), A2 => n3, ZN => n191);
   U36 : OAI21_X1 port map( B1 => n158, B2 => n98, A => n190, ZN => n126);
   U37 : NAND2_X1 port map( A1 => data_in(14), A2 => n3, ZN => n190);
   U38 : OAI21_X1 port map( B1 => n157, B2 => n98, A => n189, ZN => n125);
   U39 : NAND2_X1 port map( A1 => data_in(15), A2 => n3, ZN => n189);
   U40 : OAI21_X1 port map( B1 => n156, B2 => n98, A => n188, ZN => n124);
   U41 : NAND2_X1 port map( A1 => data_in(16), A2 => n3, ZN => n188);
   U42 : OAI21_X1 port map( B1 => n155, B2 => n98, A => n187, ZN => n123);
   U43 : NAND2_X1 port map( A1 => data_in(17), A2 => n3, ZN => n187);
   U44 : OAI21_X1 port map( B1 => n154, B2 => n98, A => n186, ZN => n122);
   U45 : NAND2_X1 port map( A1 => data_in(18), A2 => n96, ZN => n186);
   U46 : OAI21_X1 port map( B1 => n153, B2 => n98, A => n185, ZN => n121);
   U47 : NAND2_X1 port map( A1 => data_in(19), A2 => n96, ZN => n185);
   U48 : OAI21_X1 port map( B1 => n152, B2 => n98, A => n184, ZN => n120);
   U49 : NAND2_X1 port map( A1 => data_in(20), A2 => n96, ZN => n184);
   U50 : OAI21_X1 port map( B1 => n151, B2 => n98, A => n183, ZN => n119);
   U51 : NAND2_X1 port map( A1 => data_in(21), A2 => n96, ZN => n183);
   U52 : OAI21_X1 port map( B1 => n150, B2 => n98, A => n182, ZN => n118);
   U53 : NAND2_X1 port map( A1 => data_in(22), A2 => n96, ZN => n182);
   U54 : OAI21_X1 port map( B1 => n149, B2 => n98, A => n181, ZN => n117);
   U55 : NAND2_X1 port map( A1 => data_in(23), A2 => n3, ZN => n181);
   U56 : OAI21_X1 port map( B1 => n148, B2 => n96, A => n180, ZN => n116);
   U57 : NAND2_X1 port map( A1 => data_in(24), A2 => n3, ZN => n180);
   U58 : OAI21_X1 port map( B1 => n147, B2 => n98, A => n179, ZN => n115);
   U59 : NAND2_X1 port map( A1 => data_in(25), A2 => n3, ZN => n179);
   U60 : OAI21_X1 port map( B1 => n146, B2 => n96, A => n178, ZN => n114);
   U61 : NAND2_X1 port map( A1 => data_in(26), A2 => n2, ZN => n178);
   U62 : OAI21_X1 port map( B1 => n145, B2 => n96, A => n177, ZN => n113);
   U63 : NAND2_X1 port map( A1 => data_in(27), A2 => n3, ZN => n177);
   U64 : OAI21_X1 port map( B1 => n144, B2 => n96, A => n176, ZN => n112);
   U65 : NAND2_X1 port map( A1 => data_in(28), A2 => n2, ZN => n176);
   U66 : OAI21_X1 port map( B1 => n143, B2 => n96, A => n175, ZN => n111);
   U67 : NAND2_X1 port map( A1 => data_in(29), A2 => n2, ZN => n175);
   U68 : OAI21_X1 port map( B1 => n142, B2 => n96, A => n174, ZN => n110);
   U69 : NAND2_X1 port map( A1 => data_in(30), A2 => n2, ZN => n174);
   U70 : OAI21_X1 port map( B1 => n141, B2 => n96, A => n173, ZN => n109);
   U71 : NAND2_X1 port map( A1 => data_in(31), A2 => n2, ZN => n173);
   U72 : INV_X1 port map( A => n172, ZN => n106);
   U73 : MUX2_X1 port map( A => n106, B => data_in(0), S => n99, Z => n140);
   U74 : INV_X1 port map( A => n171, ZN => n107);
   U75 : MUX2_X1 port map( A => n107, B => data_in(1), S => n99, Z => n139);
   U76 : INV_X1 port map( A => n170, ZN => n108);
   U77 : MUX2_X1 port map( A => n108, B => data_in(2), S => n99, Z => n138);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_9 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_9;

architecture SYN_Behavioral of REG_NBIT32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n147);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n107, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n174);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n110, Z => n109);
   U5 : BUF_X1 port map( A => n105, Z => n98);
   U6 : BUF_X1 port map( A => n105, Z => n99);
   U7 : BUF_X1 port map( A => n105, Z => n100);
   U8 : BUF_X1 port map( A => n104, Z => n101);
   U9 : BUF_X1 port map( A => n104, Z => n102);
   U10 : BUF_X1 port map( A => n109, Z => n106);
   U11 : BUF_X1 port map( A => n109, Z => n107);
   U12 : BUF_X1 port map( A => n109, Z => n108);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : INV_X1 port map( A => reset, ZN => n110);
   U15 : BUF_X1 port map( A => enable, Z => n96);
   U16 : OAI21_X1 port map( B1 => n174, B2 => n103, A => n206, ZN => n142);
   U17 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n206);
   U18 : OAI21_X1 port map( B1 => n173, B2 => n102, A => n205, ZN => n141);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n205);
   U20 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n204);
   U22 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n203);
   U24 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n202);
   U26 : OAI21_X1 port map( B1 => n169, B2 => n101, A => n201, ZN => n137);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n201);
   U28 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n200);
   U30 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n199);
   U32 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n198, ZN => n134);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n198);
   U34 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n197, ZN => n133);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n197);
   U36 : OAI21_X1 port map( B1 => n164, B2 => n100, A => n196, ZN => n132);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n196);
   U38 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n195);
   U40 : OAI21_X1 port map( B1 => n162, B2 => n101, A => n194, ZN => n130);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n194);
   U42 : OAI21_X1 port map( B1 => n161, B2 => n100, A => n193, ZN => n129);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n193);
   U44 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n192);
   U46 : OAI21_X1 port map( B1 => n159, B2 => n101, A => n191, ZN => n127);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n191);
   U48 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n190);
   U50 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n189);
   U52 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n188);
   U54 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n187);
   U56 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n186);
   U58 : OAI21_X1 port map( B1 => n153, B2 => n102, A => n185, ZN => n121);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n185);
   U60 : OAI21_X1 port map( B1 => n152, B2 => n101, A => n184, ZN => n120);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n184);
   U62 : OAI21_X1 port map( B1 => n151, B2 => n102, A => n183, ZN => n119);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n183);
   U64 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n182);
   U66 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n181);
   U68 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n180);
   U70 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U71 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n179);
   U72 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n178);
   U74 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n177);
   U76 : OAI21_X1 port map( B1 => n144, B2 => n103, A => n176, ZN => n112);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n176);
   U78 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n175);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_8 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_8;

architecture SYN_Behavioral of REG_NBIT32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n147);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n107, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n174);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n110, Z => n109);
   U5 : BUF_X1 port map( A => n105, Z => n98);
   U6 : BUF_X1 port map( A => n105, Z => n99);
   U7 : BUF_X1 port map( A => n105, Z => n100);
   U8 : BUF_X1 port map( A => n104, Z => n101);
   U9 : BUF_X1 port map( A => n104, Z => n102);
   U10 : BUF_X1 port map( A => n109, Z => n106);
   U11 : BUF_X1 port map( A => n109, Z => n107);
   U12 : BUF_X1 port map( A => n109, Z => n108);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : INV_X1 port map( A => reset, ZN => n110);
   U15 : BUF_X1 port map( A => enable, Z => n96);
   U16 : OAI21_X1 port map( B1 => n174, B2 => n103, A => n206, ZN => n142);
   U17 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n206);
   U18 : OAI21_X1 port map( B1 => n173, B2 => n102, A => n205, ZN => n141);
   U19 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n205);
   U20 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U21 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n204);
   U22 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n203);
   U24 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n202);
   U26 : OAI21_X1 port map( B1 => n169, B2 => n101, A => n201, ZN => n137);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n201);
   U28 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n200);
   U30 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n199);
   U32 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n198, ZN => n134);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n198);
   U34 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n197, ZN => n133);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n197);
   U36 : OAI21_X1 port map( B1 => n164, B2 => n100, A => n196, ZN => n132);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n196);
   U38 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n195);
   U40 : OAI21_X1 port map( B1 => n162, B2 => n101, A => n194, ZN => n130);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n194);
   U42 : OAI21_X1 port map( B1 => n161, B2 => n100, A => n193, ZN => n129);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n193);
   U44 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n192);
   U46 : OAI21_X1 port map( B1 => n159, B2 => n101, A => n191, ZN => n127);
   U47 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n191);
   U48 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n190);
   U50 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U51 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n189);
   U52 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U53 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n188);
   U54 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U55 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n187);
   U56 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U57 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n186);
   U58 : OAI21_X1 port map( B1 => n153, B2 => n102, A => n185, ZN => n121);
   U59 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n185);
   U60 : OAI21_X1 port map( B1 => n152, B2 => n101, A => n184, ZN => n120);
   U61 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n184);
   U62 : OAI21_X1 port map( B1 => n151, B2 => n102, A => n183, ZN => n119);
   U63 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n183);
   U64 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U65 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n182);
   U66 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U67 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n181);
   U68 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U69 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n180);
   U70 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U71 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n179);
   U72 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U73 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n178);
   U74 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U75 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n177);
   U76 : OAI21_X1 port map( B1 => n144, B2 => n103, A => n176, ZN => n112);
   U77 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n176);
   U78 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n175);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_7 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_7;

architecture SYN_Behavioral of REG_NBIT32_7 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n69, n70, n71, n72, n73
      , n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270 : 
      std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_31_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n8, Q => 
                           data_out_31_port, QN => n73);
   reg_reg_30_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n8, Q => 
                           data_out_30_port, QN => n74);
   reg_reg_29_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n8, Q => 
                           data_out_29_port, QN => n75);
   reg_reg_27_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n8, Q => 
                           data_out_27_port, QN => n77);
   reg_reg_26_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n8, Q => 
                           data_out_26_port, QN => n78);
   reg_reg_25_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n8, Q => 
                           data_out_25_port, QN => n79);
   reg_reg_24_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n8, Q => 
                           data_out_24_port, QN => n80);
   reg_reg_23_inst : DFFR_X1 port map( D => n33, CK => clk, RN => n8, Q => 
                           data_out_23_port, QN => n81);
   reg_reg_22_inst : DFFR_X1 port map( D => n34, CK => clk, RN => n8, Q => 
                           data_out_22_port, QN => n82);
   reg_reg_21_inst : DFFR_X1 port map( D => n35, CK => clk, RN => n8, Q => 
                           data_out_21_port, QN => n83);
   reg_reg_20_inst : DFFR_X1 port map( D => n36, CK => clk, RN => n8, Q => 
                           data_out_20_port, QN => n84);
   reg_reg_19_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n9, Q => 
                           data_out_19_port, QN => n_1251);
   reg_reg_18_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n9, Q => 
                           data_out_18_port, QN => n_1252);
   reg_reg_17_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n9, Q => 
                           data_out_17_port, QN => n_1253);
   reg_reg_16_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n9, Q => 
                           data_out_16_port, QN => n_1254);
   reg_reg_15_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n9, Q => 
                           data_out_15_port, QN => n_1255);
   reg_reg_14_inst : DFFR_X1 port map( D => n42, CK => clk, RN => n9, Q => 
                           data_out_14_port, QN => n_1256);
   reg_reg_13_inst : DFFR_X1 port map( D => n43, CK => clk, RN => n9, Q => 
                           data_out_13_port, QN => n_1257);
   reg_reg_12_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n9, Q => 
                           data_out_12_port, QN => n_1258);
   reg_reg_11_inst : DFFR_X1 port map( D => n45, CK => clk, RN => n9, Q => 
                           data_out_11_port, QN => n_1259);
   reg_reg_10_inst : DFFR_X1 port map( D => n46, CK => clk, RN => n9, Q => 
                           data_out_10_port, QN => n_1260);
   reg_reg_9_inst : DFFR_X1 port map( D => n47, CK => clk, RN => n9, Q => 
                           data_out_9_port, QN => n_1261);
   reg_reg_8_inst : DFFR_X1 port map( D => n48, CK => clk, RN => n9, Q => 
                           data_out_8_port, QN => n_1262);
   reg_reg_7_inst : DFFR_X1 port map( D => n49, CK => clk, RN => n10, Q => 
                           data_out_7_port, QN => n_1263);
   reg_reg_6_inst : DFFR_X1 port map( D => n50, CK => clk, RN => n10, Q => 
                           data_out_6_port, QN => n_1264);
   reg_reg_5_inst : DFFR_X1 port map( D => n51, CK => clk, RN => n10, Q => 
                           data_out_5_port, QN => n_1265);
   reg_reg_4_inst : DFFR_X1 port map( D => n52, CK => clk, RN => n10, Q => 
                           data_out_4_port, QN => n_1266);
   reg_reg_3_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n10, Q => 
                           data_out_3_port, QN => n_1267);
   reg_reg_2_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n10, Q => 
                           data_out_2_port, QN => n_1268);
   reg_reg_1_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n10, Q => 
                           data_out_1_port, QN => n_1269);
   reg_reg_0_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n10, Q => 
                           data_out_0_port, QN => n_1270);
   reg_reg_28_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n8, Q => 
                           data_out_28_port, QN => n76);
   U2 : BUF_X1 port map( A => n1, Z => n6);
   U3 : BUF_X1 port map( A => n12, Z => n11);
   U4 : BUF_X1 port map( A => n6, Z => n4);
   U5 : BUF_X1 port map( A => n11, Z => n8);
   U6 : BUF_X1 port map( A => n6, Z => n3);
   U7 : BUF_X1 port map( A => n11, Z => n9);
   U8 : BUF_X1 port map( A => n11, Z => n10);
   U9 : BUF_X1 port map( A => n6, Z => n5);
   U10 : INV_X1 port map( A => reset, ZN => n12);
   U11 : BUF_X1 port map( A => n7, Z => n2);
   U12 : BUF_X1 port map( A => n1, Z => n7);
   U13 : BUF_X1 port map( A => enable, Z => n1);
   U14 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => n2, Z =>
                           n72);
   U15 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n2, Z =>
                           n71);
   U16 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => n2, Z =>
                           n70);
   U17 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => n2, Z =>
                           n69);
   U18 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => n2, Z =>
                           n52);
   U19 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n2, Z =>
                           n51);
   U20 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n2, Z =>
                           n50);
   U21 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => n2, Z =>
                           n49);
   U22 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => n2, Z =>
                           n48);
   U23 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n2, Z =>
                           n47);
   U24 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => n2, Z 
                           => n46);
   U25 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => n2, Z 
                           => n45);
   U26 : MUX2_X1 port map( A => data_out_12_port, B => data_in(12), S => n3, Z 
                           => n44);
   U27 : MUX2_X1 port map( A => data_out_13_port, B => data_in(13), S => n3, Z 
                           => n43);
   U28 : MUX2_X1 port map( A => data_out_14_port, B => data_in(14), S => n3, Z 
                           => n42);
   U29 : MUX2_X1 port map( A => data_out_15_port, B => data_in(15), S => n3, Z 
                           => n41);
   U30 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => n3, Z 
                           => n40);
   U31 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => n3, Z 
                           => n39);
   U32 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => n3, Z 
                           => n38);
   U33 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => n3, Z 
                           => n37);
   U34 : NAND2_X1 port map( A1 => data_in(20), A2 => n3, ZN => n13);
   U35 : OAI21_X1 port map( B1 => n84, B2 => n5, A => n13, ZN => n36);
   U36 : NAND2_X1 port map( A1 => data_in(21), A2 => n4, ZN => n14);
   U37 : OAI21_X1 port map( B1 => n83, B2 => n5, A => n14, ZN => n35);
   U38 : NAND2_X1 port map( A1 => data_in(22), A2 => n4, ZN => n15);
   U39 : OAI21_X1 port map( B1 => n82, B2 => n5, A => n15, ZN => n34);
   U40 : NAND2_X1 port map( A1 => data_in(23), A2 => n4, ZN => n16);
   U41 : OAI21_X1 port map( B1 => n81, B2 => n4, A => n16, ZN => n33);
   U42 : NAND2_X1 port map( A1 => data_in(24), A2 => n4, ZN => n17);
   U43 : OAI21_X1 port map( B1 => n80, B2 => n4, A => n17, ZN => n32);
   U44 : NAND2_X1 port map( A1 => data_in(25), A2 => n4, ZN => n18);
   U45 : OAI21_X1 port map( B1 => n79, B2 => n4, A => n18, ZN => n31);
   U46 : NAND2_X1 port map( A1 => data_in(26), A2 => n4, ZN => n19);
   U47 : OAI21_X1 port map( B1 => n78, B2 => n4, A => n19, ZN => n30);
   U48 : NAND2_X1 port map( A1 => data_in(27), A2 => n4, ZN => n20);
   U49 : OAI21_X1 port map( B1 => n77, B2 => n5, A => n20, ZN => n29);
   U50 : NAND2_X1 port map( A1 => data_in(28), A2 => n4, ZN => n21);
   U51 : OAI21_X1 port map( B1 => n76, B2 => n5, A => n21, ZN => n28);
   U52 : NAND2_X1 port map( A1 => data_in(29), A2 => n3, ZN => n22);
   U53 : OAI21_X1 port map( B1 => n75, B2 => n5, A => n22, ZN => n27);
   U54 : NAND2_X1 port map( A1 => data_in(30), A2 => n3, ZN => n23);
   U55 : OAI21_X1 port map( B1 => n74, B2 => n5, A => n23, ZN => n26);
   U56 : NAND2_X1 port map( A1 => data_in(31), A2 => n3, ZN => n24);
   U57 : OAI21_X1 port map( B1 => n73, B2 => n4, A => n24, ZN => n25);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_6 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_6;

architecture SYN_Behavioral of REG_NBIT32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n107, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n107, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n105, Z => n98);
   U5 : BUF_X1 port map( A => n105, Z => n99);
   U6 : BUF_X1 port map( A => n105, Z => n100);
   U7 : BUF_X1 port map( A => n104, Z => n101);
   U8 : BUF_X1 port map( A => n104, Z => n102);
   U9 : BUF_X1 port map( A => n109, Z => n106);
   U10 : BUF_X1 port map( A => n109, Z => n107);
   U11 : BUF_X1 port map( A => n109, Z => n108);
   U12 : BUF_X1 port map( A => n104, Z => n103);
   U13 : INV_X1 port map( A => reset, ZN => n109);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_5 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_5;

architecture SYN_Behavioral of REG_NBIT32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   
   reg_reg_0_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n170);
   reg_reg_8_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n162);
   reg_reg_6_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n164);
   reg_reg_5_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n165);
   reg_reg_4_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n166);
   reg_reg_3_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n167);
   reg_reg_2_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n168);
   reg_reg_1_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n169);
   reg_reg_31_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n106, Q => 
                           data_out(31), QN => n139);
   reg_reg_30_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n106, Q => 
                           data_out(30), QN => n140);
   reg_reg_14_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n106, Q => 
                           data_out(14), QN => n156);
   reg_reg_13_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n106, Q => 
                           data_out(13), QN => n157);
   reg_reg_11_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n159);
   reg_reg_10_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n160);
   reg_reg_29_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n106, Q => 
                           data_out(29), QN => n141);
   reg_reg_28_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n106, Q => 
                           data_out(28), QN => n142);
   reg_reg_27_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n106, Q => 
                           data_out(27), QN => n143);
   reg_reg_26_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n106, Q => 
                           data_out(26), QN => n144);
   reg_reg_25_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n106, Q => 
                           data_out(25), QN => n145);
   reg_reg_24_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n106, Q => 
                           data_out(24), QN => n146);
   reg_reg_23_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n106, Q => 
                           data_out(23), QN => n147);
   reg_reg_22_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n106, Q => 
                           data_out(22), QN => n148);
   reg_reg_21_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n106, Q => 
                           data_out(21), QN => n149);
   reg_reg_20_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n106, Q => 
                           data_out(20), QN => n150);
   reg_reg_19_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n106, Q => 
                           data_out(19), QN => n151);
   reg_reg_18_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n106, Q => 
                           data_out(18), QN => n152);
   reg_reg_17_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n106, Q => 
                           data_out(17), QN => n153);
   reg_reg_16_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n106, Q => 
                           data_out(16), QN => n154);
   reg_reg_15_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n106, Q => 
                           data_out(15), QN => n155);
   reg_reg_12_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n106, Q => 
                           data_out(12), QN => n158);
   reg_reg_9_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n161);
   reg_reg_7_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n163);
   U2 : INV_X2 port map( A => reset, ZN => n106);
   U3 : BUF_X1 port map( A => n96, Z => n105);
   U4 : CLKBUF_X1 port map( A => n96, Z => n104);
   U5 : BUF_X1 port map( A => n105, Z => n98);
   U6 : BUF_X1 port map( A => n105, Z => n99);
   U7 : BUF_X1 port map( A => n105, Z => n100);
   U8 : BUF_X1 port map( A => n104, Z => n103);
   U9 : BUF_X1 port map( A => n104, Z => n101);
   U10 : BUF_X1 port map( A => n104, Z => n102);
   U11 : BUF_X1 port map( A => enable, Z => n96);
   U12 : OAI21_X1 port map( B1 => n163, B2 => n101, A => n195, ZN => n131);
   U13 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n195);
   U14 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U15 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n192);
   U16 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U17 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n191);
   U18 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U19 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n190);
   U20 : OAI21_X1 port map( B1 => n157, B2 => n100, A => n189, ZN => n125);
   U21 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n189);
   U22 : OAI21_X1 port map( B1 => n156, B2 => n100, A => n188, ZN => n124);
   U23 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n188);
   U24 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U25 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n187);
   U26 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U27 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n186);
   U28 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U29 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n185);
   U30 : OAI21_X1 port map( B1 => n152, B2 => n101, A => n184, ZN => n120);
   U31 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n184);
   U32 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U33 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n183);
   U34 : OAI21_X1 port map( B1 => n150, B2 => n101, A => n182, ZN => n118);
   U35 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n182);
   U36 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U37 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n181);
   U38 : OAI21_X1 port map( B1 => n148, B2 => n101, A => n180, ZN => n116);
   U39 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n180);
   U40 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U41 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n179);
   U42 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U43 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n178);
   U44 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U45 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n177);
   U46 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U47 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n176);
   U48 : OAI21_X1 port map( B1 => n143, B2 => n102, A => n175, ZN => n111);
   U49 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n175);
   U50 : OAI21_X1 port map( B1 => n142, B2 => n102, A => n174, ZN => n110);
   U51 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n174);
   U52 : OAI21_X1 port map( B1 => n141, B2 => n102, A => n173, ZN => n109);
   U53 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n173);
   U54 : OAI21_X1 port map( B1 => n140, B2 => n103, A => n172, ZN => n108);
   U55 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n172);
   U56 : OAI21_X1 port map( B1 => n139, B2 => n103, A => n171, ZN => n107);
   U57 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n171);
   U58 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U59 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n193);
   U60 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U61 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n201);
   U62 : OAI21_X1 port map( B1 => n168, B2 => n102, A => n200, ZN => n136);
   U63 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n200);
   U64 : OAI21_X1 port map( B1 => n167, B2 => n102, A => n199, ZN => n135);
   U65 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n199);
   U66 : OAI21_X1 port map( B1 => n166, B2 => n102, A => n198, ZN => n134);
   U67 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n198);
   U68 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n197, ZN => n133);
   U69 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n197);
   U70 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U71 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n196);
   U72 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U73 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n194);
   U74 : OAI21_X1 port map( B1 => n170, B2 => n103, A => n202, ZN => n138);
   U75 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n202);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_4 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_4;

architecture SYN_Behavioral of REG_NBIT32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   
   reg_reg_0_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n170);
   reg_reg_8_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n162);
   reg_reg_6_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n164);
   reg_reg_5_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n165);
   reg_reg_4_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n166);
   reg_reg_3_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n167);
   reg_reg_2_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n168);
   reg_reg_1_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n169);
   reg_reg_31_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n106, Q => 
                           data_out(31), QN => n139);
   reg_reg_30_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n106, Q => 
                           data_out(30), QN => n140);
   reg_reg_14_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n106, Q => 
                           data_out(14), QN => n156);
   reg_reg_13_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n106, Q => 
                           data_out(13), QN => n157);
   reg_reg_11_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n159);
   reg_reg_10_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n160);
   reg_reg_29_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n106, Q => 
                           data_out(29), QN => n141);
   reg_reg_28_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n106, Q => 
                           data_out(28), QN => n142);
   reg_reg_27_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n106, Q => 
                           data_out(27), QN => n143);
   reg_reg_26_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n106, Q => 
                           data_out(26), QN => n144);
   reg_reg_25_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n106, Q => 
                           data_out(25), QN => n145);
   reg_reg_24_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n106, Q => 
                           data_out(24), QN => n146);
   reg_reg_23_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n106, Q => 
                           data_out(23), QN => n147);
   reg_reg_22_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n106, Q => 
                           data_out(22), QN => n148);
   reg_reg_21_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n106, Q => 
                           data_out(21), QN => n149);
   reg_reg_20_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n106, Q => 
                           data_out(20), QN => n150);
   reg_reg_19_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n106, Q => 
                           data_out(19), QN => n151);
   reg_reg_18_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n106, Q => 
                           data_out(18), QN => n152);
   reg_reg_17_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n106, Q => 
                           data_out(17), QN => n153);
   reg_reg_16_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n106, Q => 
                           data_out(16), QN => n154);
   reg_reg_15_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n106, Q => 
                           data_out(15), QN => n155);
   reg_reg_12_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n106, Q => 
                           data_out(12), QN => n158);
   reg_reg_9_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n161);
   reg_reg_7_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n163);
   U2 : INV_X2 port map( A => reset, ZN => n106);
   U3 : BUF_X1 port map( A => n96, Z => n105);
   U4 : CLKBUF_X1 port map( A => n96, Z => n104);
   U5 : BUF_X1 port map( A => n105, Z => n98);
   U6 : BUF_X1 port map( A => n105, Z => n99);
   U7 : BUF_X1 port map( A => n105, Z => n100);
   U8 : BUF_X1 port map( A => n104, Z => n103);
   U9 : BUF_X1 port map( A => n104, Z => n101);
   U10 : BUF_X1 port map( A => n104, Z => n102);
   U11 : BUF_X1 port map( A => enable, Z => n96);
   U12 : OAI21_X1 port map( B1 => n163, B2 => n101, A => n195, ZN => n131);
   U13 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n195);
   U14 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U15 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n193);
   U16 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U17 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n192);
   U18 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U19 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n191);
   U20 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U21 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n190);
   U22 : OAI21_X1 port map( B1 => n157, B2 => n100, A => n189, ZN => n125);
   U23 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n189);
   U24 : OAI21_X1 port map( B1 => n156, B2 => n100, A => n188, ZN => n124);
   U25 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n188);
   U26 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U27 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n187);
   U28 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U29 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n186);
   U30 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U31 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n185);
   U32 : OAI21_X1 port map( B1 => n152, B2 => n101, A => n184, ZN => n120);
   U33 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n184);
   U34 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U35 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n183);
   U36 : OAI21_X1 port map( B1 => n150, B2 => n101, A => n182, ZN => n118);
   U37 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n182);
   U38 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U39 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n181);
   U40 : OAI21_X1 port map( B1 => n148, B2 => n101, A => n180, ZN => n116);
   U41 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n180);
   U42 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U43 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n179);
   U44 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U45 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n178);
   U46 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U47 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n177);
   U48 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U49 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n176);
   U50 : OAI21_X1 port map( B1 => n143, B2 => n102, A => n175, ZN => n111);
   U51 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n175);
   U52 : OAI21_X1 port map( B1 => n142, B2 => n102, A => n174, ZN => n110);
   U53 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n174);
   U54 : OAI21_X1 port map( B1 => n141, B2 => n102, A => n173, ZN => n109);
   U55 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n173);
   U56 : OAI21_X1 port map( B1 => n140, B2 => n103, A => n172, ZN => n108);
   U57 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n172);
   U58 : OAI21_X1 port map( B1 => n139, B2 => n103, A => n171, ZN => n107);
   U59 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n171);
   U60 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U61 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n201);
   U62 : OAI21_X1 port map( B1 => n168, B2 => n102, A => n200, ZN => n136);
   U63 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n200);
   U64 : OAI21_X1 port map( B1 => n167, B2 => n102, A => n199, ZN => n135);
   U65 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n199);
   U66 : OAI21_X1 port map( B1 => n166, B2 => n102, A => n198, ZN => n134);
   U67 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n198);
   U68 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n197, ZN => n133);
   U69 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n197);
   U70 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U71 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n196);
   U72 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U73 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n194);
   U74 : OAI21_X1 port map( B1 => n170, B2 => n103, A => n202, ZN => n138);
   U75 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n202);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_3 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_3;

architecture SYN_Behavioral of REG_NBIT32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n1, Q => 
                           data_out(31), QN => n133);
   reg_reg_30_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n1, Q => 
                           data_out(30), QN => n134);
   reg_reg_29_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n1, Q => 
                           data_out(29), QN => n135);
   reg_reg_28_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n1, Q => 
                           data_out(28), QN => n136);
   reg_reg_27_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n1, Q => 
                           data_out(27), QN => n137);
   reg_reg_26_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n1, Q => 
                           data_out(26), QN => n138);
   reg_reg_25_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n1, Q => 
                           data_out(25), QN => n139);
   reg_reg_24_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n1, Q => 
                           data_out(24), QN => n140);
   reg_reg_23_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n1, Q => 
                           data_out(23), QN => n141);
   reg_reg_22_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n1, Q => 
                           data_out(22), QN => n142);
   reg_reg_21_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n1, Q => 
                           data_out(21), QN => n143);
   reg_reg_20_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n1, Q => 
                           data_out(20), QN => n144);
   reg_reg_19_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n2, Q => 
                           data_out(19), QN => n145);
   reg_reg_18_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n2, Q => 
                           data_out(18), QN => n146);
   reg_reg_17_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n2, Q => 
                           data_out(17), QN => n147);
   reg_reg_16_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n2, Q => 
                           data_out(16), QN => n148);
   reg_reg_15_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n2, Q => 
                           data_out(15), QN => n149);
   reg_reg_14_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n2, Q => 
                           data_out(14), QN => n150);
   reg_reg_13_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n2, Q => 
                           data_out(13), QN => n151);
   reg_reg_12_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n2, Q => 
                           data_out(12), QN => n152);
   reg_reg_11_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n2, Q => 
                           data_out(11), QN => n153);
   reg_reg_10_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n2, Q => 
                           data_out(10), QN => n154);
   reg_reg_9_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n2, Q => 
                           data_out(9), QN => n155);
   reg_reg_8_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n2, Q => 
                           data_out(8), QN => n156);
   reg_reg_7_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n3, Q => 
                           data_out(7), QN => n157);
   reg_reg_6_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n3, Q => 
                           data_out(6), QN => n158);
   reg_reg_5_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n3, Q => 
                           data_out(5), QN => n159);
   reg_reg_4_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n3, Q => 
                           data_out(4), QN => n160);
   reg_reg_3_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n3, Q => 
                           data_out(3), QN => n161);
   reg_reg_2_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n3, Q => 
                           data_out(2), QN => n162);
   reg_reg_1_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n3, Q => 
                           data_out(1), QN => n163);
   reg_reg_0_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n3, Q => 
                           data_out(0), QN => n164);
   U2 : BUF_X1 port map( A => n100, Z => n2);
   U3 : BUF_X1 port map( A => n100, Z => n1);
   U4 : BUF_X1 port map( A => n100, Z => n3);
   U5 : INV_X1 port map( A => n164, ZN => n4);
   U6 : MUX2_X1 port map( A => n4, B => data_in(0), S => enable, Z => n132);
   U7 : INV_X1 port map( A => reset, ZN => n100);
   U8 : INV_X1 port map( A => n163, ZN => n5);
   U9 : MUX2_X1 port map( A => n5, B => data_in(1), S => enable, Z => n131);
   U10 : INV_X1 port map( A => n162, ZN => n6);
   U11 : MUX2_X1 port map( A => n6, B => data_in(2), S => enable, Z => n130);
   U12 : INV_X1 port map( A => n161, ZN => n7);
   U13 : MUX2_X1 port map( A => n7, B => data_in(3), S => enable, Z => n129);
   U14 : INV_X1 port map( A => n160, ZN => n8);
   U15 : MUX2_X1 port map( A => n8, B => data_in(4), S => enable, Z => n128);
   U16 : INV_X1 port map( A => n159, ZN => n9);
   U17 : MUX2_X1 port map( A => n9, B => data_in(5), S => enable, Z => n127);
   U18 : INV_X1 port map( A => n158, ZN => n10);
   U19 : MUX2_X1 port map( A => n10, B => data_in(6), S => enable, Z => n126);
   U20 : INV_X1 port map( A => n157, ZN => n11);
   U21 : MUX2_X1 port map( A => n11, B => data_in(7), S => enable, Z => n125);
   U22 : INV_X1 port map( A => n156, ZN => n12);
   U23 : MUX2_X1 port map( A => n12, B => data_in(8), S => enable, Z => n124);
   U24 : INV_X1 port map( A => n155, ZN => n13);
   U25 : MUX2_X1 port map( A => n13, B => data_in(9), S => enable, Z => n123);
   U26 : INV_X1 port map( A => n154, ZN => n14);
   U27 : MUX2_X1 port map( A => n14, B => data_in(10), S => enable, Z => n122);
   U28 : INV_X1 port map( A => n153, ZN => n15);
   U29 : MUX2_X1 port map( A => n15, B => data_in(11), S => enable, Z => n121);
   U30 : INV_X1 port map( A => n152, ZN => n16);
   U31 : MUX2_X1 port map( A => n16, B => data_in(12), S => enable, Z => n120);
   U32 : INV_X1 port map( A => n151, ZN => n17);
   U33 : MUX2_X1 port map( A => n17, B => data_in(13), S => enable, Z => n119);
   U34 : INV_X1 port map( A => n150, ZN => n18);
   U35 : MUX2_X1 port map( A => n18, B => data_in(14), S => enable, Z => n118);
   U36 : INV_X1 port map( A => n149, ZN => n19);
   U37 : MUX2_X1 port map( A => n19, B => data_in(15), S => enable, Z => n117);
   U38 : INV_X1 port map( A => n148, ZN => n20);
   U39 : MUX2_X1 port map( A => n20, B => data_in(16), S => enable, Z => n116);
   U40 : INV_X1 port map( A => n147, ZN => n21);
   U41 : MUX2_X1 port map( A => n21, B => data_in(17), S => enable, Z => n115);
   U42 : INV_X1 port map( A => n146, ZN => n22);
   U43 : MUX2_X1 port map( A => n22, B => data_in(18), S => enable, Z => n114);
   U44 : INV_X1 port map( A => n145, ZN => n23);
   U45 : MUX2_X1 port map( A => n23, B => data_in(19), S => enable, Z => n113);
   U46 : INV_X1 port map( A => n144, ZN => n24);
   U47 : MUX2_X1 port map( A => n24, B => data_in(20), S => enable, Z => n112);
   U48 : INV_X1 port map( A => n143, ZN => n25);
   U49 : MUX2_X1 port map( A => n25, B => data_in(21), S => enable, Z => n111);
   U50 : INV_X1 port map( A => n142, ZN => n26);
   U51 : MUX2_X1 port map( A => n26, B => data_in(22), S => enable, Z => n110);
   U52 : INV_X1 port map( A => n141, ZN => n27);
   U53 : MUX2_X1 port map( A => n27, B => data_in(23), S => enable, Z => n109);
   U54 : INV_X1 port map( A => n140, ZN => n28);
   U55 : MUX2_X1 port map( A => n28, B => data_in(24), S => enable, Z => n108);
   U56 : INV_X1 port map( A => n139, ZN => n29);
   U57 : MUX2_X1 port map( A => n29, B => data_in(25), S => enable, Z => n107);
   U58 : INV_X1 port map( A => n138, ZN => n30);
   U59 : MUX2_X1 port map( A => n30, B => data_in(26), S => enable, Z => n106);
   U60 : INV_X1 port map( A => n137, ZN => n31);
   U61 : MUX2_X1 port map( A => n31, B => data_in(27), S => enable, Z => n105);
   U62 : INV_X1 port map( A => n136, ZN => n32);
   U63 : MUX2_X1 port map( A => n32, B => data_in(28), S => enable, Z => n104);
   U64 : INV_X1 port map( A => n135, ZN => n96);
   U65 : MUX2_X1 port map( A => n96, B => data_in(29), S => enable, Z => n103);
   U66 : INV_X1 port map( A => n134, ZN => n98);
   U67 : MUX2_X1 port map( A => n98, B => data_in(30), S => enable, Z => n102);
   U68 : INV_X1 port map( A => n133, ZN => n99);
   U69 : MUX2_X1 port map( A => n99, B => data_in(31), S => enable, Z => n101);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_2 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_2;

architecture SYN_Behavioral of REG_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      data_out_16_port, data_out_17_port, data_out_18_port, data_out_19_port, 
      data_out_20_port, data_out_21_port, data_out_22_port, data_out_23_port, 
      data_out_24_port, data_out_25_port, data_out_26_port, data_out_27_port, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n23, Q => 
                           data_out_15_port, QN => n147);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n23, Q => 
                           data_out_14_port, QN => n148);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n23, Q => 
                           data_out_13_port, QN => n149);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n23, Q => 
                           data_out_12_port, QN => n150);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n23, Q => 
                           data_out_11_port, QN => n151);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n23, Q => 
                           data_out_10_port, QN => n152);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n23, Q => 
                           data_out_9_port, QN => n153);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n23, Q => 
                           data_out_8_port, QN => n154);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n24, Q => 
                           data_out_7_port, QN => n155);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n24, Q => 
                           data_out_6_port, QN => n156);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n24, Q => 
                           data_out_5_port, QN => n157);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n24, Q => 
                           data_out_4_port, QN => n158);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n24, Q => 
                           data_out_3_port, QN => n159);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n24, Q => 
                           data_out_2_port, QN => n160);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n24, Q => 
                           data_out_1_port, QN => n161);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n24, Q => 
                           data_out_0_port, QN => n162);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n110, Q => 
                           data_out_19_port, QN => n_1271);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n110, Q => 
                           data_out_18_port, QN => n_1272);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n110, Q => 
                           data_out_17_port, QN => n_1273);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n110, Q => 
                           data_out_16_port, QN => n_1274);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n110, Q => 
                           data_out_21_port, QN => n_1275);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n110, Q => 
                           data_out_20_port, QN => n_1276);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n110, Q => 
                           data_out_26_port, QN => n_1277);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n110, Q => 
                           data_out_24_port, QN => n_1278);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n110, Q => 
                           data_out_25_port, QN => n_1279);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n110, Q => 
                           data_out_30_port, QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n110, Q => 
                           data_out_29_port, QN => n145);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n110, Q => 
                           data_out_28_port, QN => n146);
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n110, Q => 
                           data_out_31_port, QN => n143);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n110, Q => 
                           data_out_23_port, QN => n_1280);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n110, Q => 
                           data_out_22_port, QN => n_1281);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n110, Q => 
                           data_out_27_port, QN => n_1282);
   U2 : OR2_X2 port map( A1 => n144, A2 => enable, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n108, A2 => n1, ZN => n112);
   U4 : OR2_X2 port map( A1 => n146, A2 => enable, ZN => n2);
   U5 : NAND2_X1 port map( A1 => n106, A2 => n2, ZN => n114);
   U6 : INV_X1 port map( A => enable, ZN => n21);
   U7 : OR2_X1 port map( A1 => n143, A2 => enable, ZN => n4);
   U8 : OR2_X1 port map( A1 => n145, A2 => enable, ZN => n3);
   U9 : INV_X1 port map( A => enable, ZN => n18);
   U10 : INV_X1 port map( A => enable, ZN => n17);
   U11 : NAND2_X1 port map( A1 => n107, A2 => n3, ZN => n113);
   U12 : NAND2_X1 port map( A1 => n109, A2 => n4, ZN => n111);
   U13 : NAND2_X1 port map( A1 => data_in(26), A2 => n5, ZN => n6);
   U14 : NAND2_X1 port map( A1 => data_out_26_port, A2 => n22, ZN => n7);
   U15 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => n116);
   U16 : INV_X1 port map( A => n22, ZN => n5);
   U17 : INV_X1 port map( A => enable, ZN => n22);
   U18 : NAND2_X1 port map( A1 => data_in(21), A2 => n8, ZN => n9);
   U19 : NAND2_X1 port map( A1 => data_out_21_port, A2 => n19, ZN => n10);
   U20 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n121);
   U21 : INV_X1 port map( A => n19, ZN => n8);
   U22 : INV_X1 port map( A => enable, ZN => n19);
   U23 : NAND2_X1 port map( A1 => data_in(20), A2 => n5, ZN => n11);
   U24 : NAND2_X1 port map( A1 => data_out_20_port, A2 => n20, ZN => n12);
   U25 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n122);
   U26 : INV_X1 port map( A => enable, ZN => n20);
   U27 : NAND2_X1 port map( A1 => data_in(25), A2 => n8, ZN => n13);
   U28 : NAND2_X1 port map( A1 => data_out_25_port, A2 => n18, ZN => n14);
   U29 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n117);
   U30 : NAND2_X1 port map( A1 => data_in(24), A2 => n5, ZN => n15);
   U31 : NAND2_X1 port map( A1 => data_out_24_port, A2 => n17, ZN => n16);
   U32 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => n118);
   U33 : MUX2_X1 port map( A => data_in(23), B => data_out_23_port, S => n17, Z
                           => n119);
   U34 : MUX2_X1 port map( A => data_in(22), B => data_out_22_port, S => n18, Z
                           => n120);
   U35 : MUX2_X1 port map( A => data_in(27), B => data_out_27_port, S => n21, Z
                           => n115);
   U36 : BUF_X1 port map( A => n110, Z => n25);
   U37 : BUF_X1 port map( A => n25, Z => n23);
   U38 : BUF_X1 port map( A => n25, Z => n24);
   U39 : INV_X1 port map( A => n162, ZN => n26);
   U40 : MUX2_X1 port map( A => n26, B => data_in(0), S => enable, Z => n142);
   U41 : INV_X1 port map( A => reset, ZN => n110);
   U42 : INV_X1 port map( A => n161, ZN => n27);
   U43 : MUX2_X1 port map( A => n27, B => data_in(1), S => enable, Z => n141);
   U44 : INV_X1 port map( A => n160, ZN => n28);
   U45 : MUX2_X1 port map( A => n28, B => data_in(2), S => enable, Z => n140);
   U46 : INV_X1 port map( A => n159, ZN => n29);
   U47 : MUX2_X1 port map( A => n29, B => data_in(3), S => enable, Z => n139);
   U48 : INV_X1 port map( A => n158, ZN => n30);
   U49 : MUX2_X1 port map( A => n30, B => data_in(4), S => enable, Z => n138);
   U50 : INV_X1 port map( A => n157, ZN => n31);
   U51 : MUX2_X1 port map( A => n31, B => data_in(5), S => enable, Z => n137);
   U52 : INV_X1 port map( A => n156, ZN => n32);
   U53 : MUX2_X1 port map( A => n32, B => data_in(6), S => enable, Z => n136);
   U54 : INV_X1 port map( A => n155, ZN => n49);
   U55 : MUX2_X1 port map( A => n49, B => data_in(7), S => enable, Z => n135);
   U56 : INV_X1 port map( A => n154, ZN => n50);
   U57 : MUX2_X1 port map( A => n50, B => data_in(8), S => enable, Z => n134);
   U58 : INV_X1 port map( A => n153, ZN => n51);
   U59 : MUX2_X1 port map( A => n51, B => data_in(9), S => enable, Z => n133);
   U60 : INV_X1 port map( A => n152, ZN => n52);
   U61 : MUX2_X1 port map( A => n52, B => data_in(10), S => enable, Z => n132);
   U62 : INV_X1 port map( A => n151, ZN => n53);
   U63 : MUX2_X1 port map( A => n53, B => data_in(11), S => enable, Z => n131);
   U64 : INV_X1 port map( A => n150, ZN => n54);
   U65 : MUX2_X1 port map( A => n54, B => data_in(12), S => enable, Z => n130);
   U66 : INV_X1 port map( A => n149, ZN => n55);
   U67 : MUX2_X1 port map( A => n55, B => data_in(13), S => enable, Z => n129);
   U68 : INV_X1 port map( A => n148, ZN => n56);
   U69 : MUX2_X1 port map( A => n56, B => data_in(14), S => enable, Z => n128);
   U70 : INV_X1 port map( A => n147, ZN => n57);
   U71 : MUX2_X1 port map( A => n57, B => data_in(15), S => enable, Z => n127);
   U72 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => enable
                           , Z => n126);
   U73 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => enable
                           , Z => n125);
   U74 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => enable
                           , Z => n124);
   U75 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => enable
                           , Z => n123);
   U76 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n106);
   U77 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n107);
   U78 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n108);
   U79 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n109);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_1 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_1;

architecture SYN_Behavioral of REG_NBIT32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_20_port, n1, n2, n3, n4, data_out_0_port, data_out_1_port, 
      data_out_2_port, data_out_3_port, data_out_4_port, data_out_5_port, 
      data_out_6_port, data_out_7_port, data_out_8_port, data_out_9_port, 
      data_out_10_port, data_out_11_port, data_out_12_port, data_out_13_port, 
      data_out_14_port, data_out_15_port, data_out_16_port, data_out_17_port, 
      data_out_18_port, data_out_19_port, data_out_21_port, data_out_22_port, 
      data_out_23_port, data_out_24_port, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_1_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n3, Q => 
                           data_out_1_port, QN => n_1283);
   reg_reg_0_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n3, Q => 
                           data_out_0_port, QN => n_1284);
   reg_reg_2_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n33, Q => 
                           data_out_2_port, QN => n_1285);
   reg_reg_3_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n33, Q => 
                           data_out_3_port, QN => n_1286);
   reg_reg_6_inst : DFFR_X1 port map( D => n59, CK => clk, RN => n33, Q => 
                           data_out_6_port, QN => n_1287);
   reg_reg_5_inst : DFFR_X1 port map( D => n60, CK => clk, RN => n33, Q => 
                           data_out_5_port, QN => n_1288);
   reg_reg_4_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n33, Q => 
                           data_out_4_port, QN => n_1289);
   reg_reg_7_inst : DFFR_X1 port map( D => n58, CK => clk, RN => n33, Q => 
                           data_out_7_port, QN => n_1290);
   reg_reg_10_inst : DFFR_X1 port map( D => n55, CK => clk, RN => n33, Q => 
                           data_out_10_port, QN => n_1291);
   reg_reg_9_inst : DFFR_X1 port map( D => n56, CK => clk, RN => n33, Q => 
                           data_out_9_port, QN => n_1292);
   reg_reg_8_inst : DFFR_X1 port map( D => n57, CK => clk, RN => n33, Q => 
                           data_out_8_port, QN => n_1293);
   reg_reg_11_inst : DFFR_X1 port map( D => n54, CK => clk, RN => n33, Q => 
                           data_out_11_port, QN => n_1294);
   reg_reg_15_inst : DFFR_X1 port map( D => n50, CK => clk, RN => n33, Q => 
                           data_out_15_port, QN => n_1295);
   reg_reg_14_inst : DFFR_X1 port map( D => n51, CK => clk, RN => n33, Q => 
                           data_out_14_port, QN => n_1296);
   reg_reg_13_inst : DFFR_X1 port map( D => n52, CK => clk, RN => n33, Q => 
                           data_out_13_port, QN => n_1297);
   reg_reg_12_inst : DFFR_X1 port map( D => n53, CK => clk, RN => n33, Q => 
                           data_out_12_port, QN => n_1298);
   reg_reg_19_inst : DFFR_X1 port map( D => n46, CK => clk, RN => n33, Q => 
                           data_out_19_port, QN => n_1299);
   reg_reg_18_inst : DFFR_X1 port map( D => n47, CK => clk, RN => n33, Q => 
                           data_out_18_port, QN => n_1300);
   reg_reg_17_inst : DFFR_X1 port map( D => n48, CK => clk, RN => n33, Q => 
                           data_out_17_port, QN => n_1301);
   reg_reg_16_inst : DFFR_X1 port map( D => n49, CK => clk, RN => n33, Q => 
                           data_out_16_port, QN => n_1302);
   reg_reg_31_inst : DFFR_X1 port map( D => n34, CK => clk, RN => n33, Q => 
                           data_out_31_port, QN => n75);
   reg_reg_30_inst : DFFR_X1 port map( D => n35, CK => clk, RN => n33, Q => 
                           data_out_30_port, QN => n76);
   reg_reg_29_inst : DFFR_X1 port map( D => n36, CK => clk, RN => n33, Q => 
                           data_out_29_port, QN => n77);
   reg_reg_28_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n33, Q => 
                           data_out_28_port, QN => n78);
   reg_reg_24_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n33, Q => 
                           data_out_24_port, QN => n_1303);
   reg_reg_23_inst : DFFR_X1 port map( D => n42, CK => clk, RN => n33, Q => 
                           data_out_23_port, QN => n_1304);
   reg_reg_22_inst : DFFR_X1 port map( D => n43, CK => clk, RN => n33, Q => 
                           data_out_22_port, QN => n_1305);
   reg_reg_21_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n33, Q => 
                           data_out_21_port, QN => n_1306);
   reg_reg_20_inst : DFFR_X1 port map( D => n45, CK => clk, RN => n33, Q => 
                           data_out_20_port, QN => n_1307);
   reg_reg_27_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n33, Q => 
                           data_out_27_port, QN => n_1308);
   reg_reg_26_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n33, Q => 
                           data_out_26_port, QN => n_1309);
   reg_reg_25_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n33, Q => 
                           data_out_25_port, QN => n_1310);
   U2 : INV_X1 port map( A => enable, ZN => n1);
   U3 : INV_X2 port map( A => reset, ZN => n33);
   U4 : MUX2_X1 port map( A => data_out_20_port, B => data_in(20), S => enable,
                           Z => n45);
   U5 : MUX2_X1 port map( A => data_out_27_port, B => data_in(27), S => enable,
                           Z => n38);
   U6 : MUX2_X1 port map( A => data_out_26_port, B => data_in(26), S => enable,
                           Z => n39);
   U7 : MUX2_X1 port map( A => data_out_25_port, B => data_in(25), S => enable,
                           Z => n40);
   U8 : MUX2_X1 port map( A => data_in(24), B => data_out_24_port, S => n1, Z 
                           => n41);
   U9 : OR2_X2 port map( A1 => n75, A2 => enable, ZN => n2);
   U10 : NAND2_X1 port map( A1 => n32, A2 => n2, ZN => n34);
   U11 : BUF_X1 port map( A => n33, Z => n4);
   U12 : BUF_X1 port map( A => n4, Z => n3);
   U13 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => enable, 
                           Z => n74);
   U14 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => enable, 
                           Z => n73);
   U15 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => enable, 
                           Z => n72);
   U16 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => enable, 
                           Z => n71);
   U17 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => enable, 
                           Z => n70);
   U18 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => enable, 
                           Z => n60);
   U19 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => enable, 
                           Z => n59);
   U20 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => enable, 
                           Z => n58);
   U21 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => enable, 
                           Z => n57);
   U22 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => enable, 
                           Z => n56);
   U23 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => enable
                           , Z => n55);
   U24 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => enable
                           , Z => n54);
   U25 : MUX2_X1 port map( A => data_out_12_port, B => data_in(12), S => enable
                           , Z => n53);
   U26 : MUX2_X1 port map( A => data_out_13_port, B => data_in(13), S => enable
                           , Z => n52);
   U27 : MUX2_X1 port map( A => data_out_14_port, B => data_in(14), S => enable
                           , Z => n51);
   U28 : MUX2_X1 port map( A => data_out_15_port, B => data_in(15), S => enable
                           , Z => n50);
   U29 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => enable
                           , Z => n49);
   U30 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => enable
                           , Z => n48);
   U31 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => enable
                           , Z => n47);
   U32 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => enable
                           , Z => n46);
   U33 : MUX2_X1 port map( A => data_out_21_port, B => data_in(21), S => enable
                           , Z => n44);
   U34 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => enable
                           , Z => n43);
   U35 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => enable
                           , Z => n42);
   U36 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n29);
   U37 : OAI21_X1 port map( B1 => n78, B2 => enable, A => n29, ZN => n37);
   U38 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n30);
   U39 : OAI21_X1 port map( B1 => n77, B2 => enable, A => n30, ZN => n36);
   U40 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n31);
   U41 : OAI21_X1 port map( B1 => n76, B2 => enable, A => n31, ZN => n35);
   U42 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n32);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_0;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : AOI22_X1 port map( A1 => B(3), A2 => SEL, B1 => A(3), B2 => n1, ZN => 
                           n2);
   U6 : INV_X1 port map( A => n2, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_0;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n18, A2 => n17, ZN => n19);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n15);
   U3 : NAND2_X1 port map( A1 => n16, A2 => n15, ZN => n17);
   U4 : XNOR2_X1 port map( A => n20, B => n19, ZN => S(2));
   U5 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n20);
   U6 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U7 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => Ci, ZN => n2);
   U8 : INV_X1 port map( A => A(3), ZN => n10);
   U9 : INV_X1 port map( A => B(3), ZN => n9);
   U10 : INV_X1 port map( A => A(2), ZN => n7);
   U11 : INV_X1 port map( A => B(2), ZN => n6);
   U12 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n18);
   U13 : INV_X1 port map( A => n18, ZN => n4);
   U14 : INV_X1 port map( A => A(1), ZN => n12);
   U15 : INV_X1 port map( A => B(1), ZN => n3);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n3, ZN => n16);
   U17 : OAI221_X1 port map( B1 => B(2), B2 => A(2), C1 => n4, C2 => n15, A => 
                           n16, ZN => n5);
   U18 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n5, ZN => n21);
   U19 : OAI21_X1 port map( B1 => B(3), B2 => A(3), A => n21, ZN => n8);
   U20 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => Co);
   U21 : XOR2_X1 port map( A => B(0), B => A(0), Z => n11);
   U22 : XOR2_X1 port map( A => Ci, B => n11, Z => S(0));
   U23 : XOR2_X1 port map( A => n12, B => B(1), Z => n14);
   U24 : INV_X1 port map( A => n15, ZN => n13);
   U25 : XOR2_X1 port map( A => n14, B => n13, Z => S(1));
   U26 : XOR2_X1 port map( A => n21, B => A(3), Z => n22);
   U27 : XOR2_X1 port map( A => n22, B => B(3), Z => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_0;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_0 is

   component MUX2to1_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_127
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1311, n_1312 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1311);
   RCA0 : RCAN_NBIT4_127 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1312);
   MUX21 : MUX2to1_NBIT4_0 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_0 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_0;

architecture SYN_BEHAVIORAL of PG_block_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_0 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_0;

architecture SYN_BEHAVIORAL of G_block_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B, A => A(0), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_0;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => A(7), A2 => B(7), ZN => Gout(7));
   U2 : AND2_X1 port map( A1 => A(6), A2 => B(6), ZN => Gout(6));
   U3 : AND2_X1 port map( A1 => A(29), A2 => B(29), ZN => Gout(29));
   U4 : AND2_X1 port map( A1 => A(28), A2 => B(28), ZN => Gout(28));
   U5 : INV_X1 port map( A => B(0), ZN => n2);
   U6 : INV_X1 port map( A => A(0), ZN => n1);
   U7 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Gout(0));
   U8 : INV_X1 port map( A => A(1), ZN => n4);
   U9 : INV_X1 port map( A => B(1), ZN => n3);
   U10 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Gout(1));
   U11 : INV_X1 port map( A => A(2), ZN => n6);
   U12 : INV_X1 port map( A => B(2), ZN => n5);
   U13 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Gout(2));
   U14 : INV_X1 port map( A => A(3), ZN => n8);
   U15 : INV_X1 port map( A => B(3), ZN => n7);
   U16 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => Gout(3));
   U17 : INV_X1 port map( A => A(4), ZN => n10);
   U18 : INV_X1 port map( A => B(4), ZN => n9);
   U19 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => Gout(4));
   U20 : INV_X1 port map( A => A(5), ZN => n12);
   U21 : INV_X1 port map( A => B(5), ZN => n11);
   U22 : NOR2_X1 port map( A1 => n12, A2 => n11, ZN => Gout(5));
   U23 : INV_X1 port map( A => A(8), ZN => n14);
   U24 : INV_X1 port map( A => B(8), ZN => n13);
   U25 : NOR2_X1 port map( A1 => n14, A2 => n13, ZN => Gout(8));
   U26 : INV_X1 port map( A => A(9), ZN => n16);
   U27 : INV_X1 port map( A => B(9), ZN => n15);
   U28 : NOR2_X1 port map( A1 => n16, A2 => n15, ZN => Gout(9));
   U29 : INV_X1 port map( A => A(10), ZN => n18);
   U30 : INV_X1 port map( A => B(10), ZN => n17);
   U31 : NOR2_X1 port map( A1 => n18, A2 => n17, ZN => Gout(10));
   U32 : INV_X1 port map( A => A(11), ZN => n20);
   U33 : INV_X1 port map( A => B(11), ZN => n19);
   U34 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => Gout(11));
   U35 : INV_X1 port map( A => A(12), ZN => n22);
   U36 : INV_X1 port map( A => B(12), ZN => n21);
   U37 : NOR2_X1 port map( A1 => n22, A2 => n21, ZN => Gout(12));
   U38 : INV_X1 port map( A => A(13), ZN => n24);
   U39 : INV_X1 port map( A => B(13), ZN => n23);
   U40 : NOR2_X1 port map( A1 => n24, A2 => n23, ZN => Gout(13));
   U41 : INV_X1 port map( A => A(14), ZN => n26);
   U42 : INV_X1 port map( A => B(14), ZN => n25);
   U43 : NOR2_X1 port map( A1 => n26, A2 => n25, ZN => Gout(14));
   U44 : INV_X1 port map( A => A(15), ZN => n28);
   U45 : INV_X1 port map( A => B(15), ZN => n27);
   U46 : NOR2_X1 port map( A1 => n28, A2 => n27, ZN => Gout(15));
   U47 : INV_X1 port map( A => A(16), ZN => n30);
   U48 : INV_X1 port map( A => B(16), ZN => n29);
   U49 : NOR2_X1 port map( A1 => n30, A2 => n29, ZN => Gout(16));
   U50 : INV_X1 port map( A => A(17), ZN => n32);
   U51 : INV_X1 port map( A => B(17), ZN => n31);
   U52 : NOR2_X1 port map( A1 => n32, A2 => n31, ZN => Gout(17));
   U53 : INV_X1 port map( A => A(18), ZN => n34);
   U54 : INV_X1 port map( A => B(18), ZN => n33);
   U55 : NOR2_X1 port map( A1 => n34, A2 => n33, ZN => Gout(18));
   U56 : INV_X1 port map( A => A(19), ZN => n36);
   U57 : INV_X1 port map( A => B(19), ZN => n35);
   U58 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => Gout(19));
   U59 : INV_X1 port map( A => A(20), ZN => n38);
   U60 : INV_X1 port map( A => B(20), ZN => n37);
   U61 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => Gout(20));
   U62 : INV_X1 port map( A => A(21), ZN => n40);
   U63 : INV_X1 port map( A => B(21), ZN => n39);
   U65 : NOR2_X1 port map( A1 => n40, A2 => n39, ZN => Gout(21));
   U66 : INV_X1 port map( A => A(22), ZN => n42);
   U67 : INV_X1 port map( A => B(22), ZN => n41);
   U68 : NOR2_X1 port map( A1 => n42, A2 => n41, ZN => Gout(22));
   U69 : INV_X1 port map( A => A(23), ZN => n44);
   U70 : INV_X1 port map( A => B(23), ZN => n43);
   U71 : NOR2_X1 port map( A1 => n44, A2 => n43, ZN => Gout(23));
   U72 : INV_X1 port map( A => A(24), ZN => n46);
   U73 : INV_X1 port map( A => B(24), ZN => n45);
   U74 : NOR2_X1 port map( A1 => n46, A2 => n45, ZN => Gout(24));
   U75 : INV_X1 port map( A => A(25), ZN => n48);
   U76 : INV_X1 port map( A => B(25), ZN => n47);
   U77 : NOR2_X1 port map( A1 => n48, A2 => n47, ZN => Gout(25));
   U78 : INV_X1 port map( A => A(26), ZN => n50);
   U79 : INV_X1 port map( A => B(26), ZN => n49);
   U80 : NOR2_X1 port map( A1 => n50, A2 => n49, ZN => Gout(26));
   U81 : INV_X1 port map( A => A(27), ZN => n52);
   U82 : INV_X1 port map( A => B(27), ZN => n51);
   U83 : NOR2_X1 port map( A1 => n52, A2 => n51, ZN => Gout(27));
   U84 : INV_X1 port map( A => A(30), ZN => n54);
   U85 : INV_X1 port map( A => B(30), ZN => n53);
   U86 : NOR2_X1 port map( A1 => n54, A2 => n53, ZN => Gout(30));
   U87 : INV_X1 port map( A => A(31), ZN => n56);
   U88 : INV_X1 port map( A => B(31), ZN => n55);
   U89 : NOR2_X1 port map( A1 => n56, A2 => n55, ZN => Gout(31));
   U90 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U91 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U92 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U93 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U94 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U95 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U96 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U97 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U98 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U99 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U100 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U101 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U102 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U103 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U104 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U105 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U106 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U107 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U108 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U109 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U110 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U111 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U112 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U113 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U114 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U115 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U116 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U117 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U118 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U119 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U120 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_0 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_0;

architecture SYN_BEHAVIORAL of ENCODER_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n1, n2 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n4);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n3, A3 => n4, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n5, ZN => OUTPUT(0));
   U3 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n5, ZN => OUTPUT(1));
   U4 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => n5);
   U6 : INV_X1 port map( A => n4, ZN => n2);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_0 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_0;

architecture SYN_ARCH1 of ND4_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_0 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_0;

architecture SYN_ARCH1 of ND3_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 is

   component CARRY_SEL_N_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_63 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_62 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_61 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_60 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_59 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_58 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_57 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_64
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_65
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_66
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_67
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_190
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_191
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_68
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_69
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_192
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_193
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_194
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_70
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_195
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_196
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_197
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_198
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_199
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_200
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_201
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_71
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_202
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_203
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_204
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_205
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_206
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_207
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_208
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_209
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_210
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_211
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_212
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_213
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_214
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_215
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_0
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_0
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, n9,
      Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, 
      P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, 
      P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, 
      P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, 
      P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, 
      P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, Co_2_port, n2, n3, n4, n5, n6, n8, n_1313 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_0 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1313, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n8);
   gblock1_1_1 : G_block_0 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B 
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_0 port map( A(1) => P_4_4_port, A(0) => G_4_4_port, 
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_215 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_214 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_213 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_212 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_211 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_210 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_209 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_208 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_207 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_206 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_205 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_204 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_203 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_202 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_71 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_201 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_200 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_199 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_198 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_197 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_196 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_195 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_70 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => n9);
   pgblock1_3_2 : PG_block_194 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_193 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_192 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_69 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => n9, Gout => Co_3_port);
   gblock2_4_4 : G_block_68 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_191 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_190 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_67 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_66 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_65 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_64 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : BUF_X1 port map( A => n9, Z => Co_2_port);
   U2 : INV_X1 port map( A => A(0), ZN => n4);
   U3 : INV_X1 port map( A => Cin, ZN => n3);
   U4 : INV_X1 port map( A => B(0), ZN => n2);
   U5 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => n5);
   U6 : OAI211_X1 port map( C1 => Cin, C2 => A(0), A => n5, B => n8, ZN => n6);
   U7 : INV_X1 port map( A => n6, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUL is

   port( CLOCK : in std_logic;  A, B : in std_logic_vector (15 downto 0);  Y : 
         out std_logic_vector (31 downto 0));

end MUL;

architecture SYN_BEHAVIORAL of MUL is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_1
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_4
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_2
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_5
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_6
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_3
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_7
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component MUX5to1_NBIT32_1
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_2
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_3
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_4
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_5
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_6
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_7
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_8
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component ENCODER_1
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_2
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_3
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_4
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_5
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_6
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_7
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_0
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, A_neg_15_30_port, A_neg_15_29_port, 
      A_neg_15_28_port, A_neg_15_27_port, A_neg_15_26_port, A_neg_15_25_port, 
      A_neg_15_24_port, A_neg_15_23_port, A_neg_15_22_port, A_neg_15_21_port, 
      A_neg_15_20_port, A_neg_15_19_port, A_neg_15_18_port, A_neg_15_17_port, 
      A_neg_15_16_port, A_neg_14_29_port, A_neg_14_28_port, A_neg_14_27_port, 
      A_neg_14_26_port, A_neg_14_25_port, A_neg_14_24_port, A_neg_14_23_port, 
      A_neg_14_22_port, A_neg_14_21_port, A_neg_14_20_port, A_neg_14_19_port, 
      A_neg_14_18_port, A_neg_14_17_port, A_neg_14_16_port, A_neg_14_15_port, 
      A_neg_13_28_port, A_neg_13_27_port, A_neg_13_26_port, A_neg_13_25_port, 
      A_neg_13_24_port, A_neg_13_23_port, A_neg_13_22_port, A_neg_13_21_port, 
      A_neg_13_20_port, A_neg_13_19_port, A_neg_13_18_port, A_neg_13_17_port, 
      A_neg_13_16_port, A_neg_13_15_port, A_neg_13_14_port, A_neg_12_27_port, 
      A_neg_12_26_port, A_neg_12_25_port, A_neg_12_24_port, A_neg_12_23_port, 
      A_neg_12_22_port, A_neg_12_21_port, A_neg_12_20_port, A_neg_12_19_port, 
      A_neg_12_18_port, A_neg_12_17_port, A_neg_12_16_port, A_neg_12_15_port, 
      A_neg_12_14_port, A_neg_12_13_port, A_neg_11_26_port, A_neg_11_25_port, 
      A_neg_11_24_port, A_neg_11_23_port, A_neg_11_22_port, A_neg_11_21_port, 
      A_neg_11_20_port, A_neg_11_19_port, A_neg_11_18_port, A_neg_11_17_port, 
      A_neg_11_16_port, A_neg_11_15_port, A_neg_11_14_port, A_neg_11_13_port, 
      A_neg_11_12_port, A_neg_10_25_port, A_neg_10_24_port, A_neg_10_23_port, 
      A_neg_10_22_port, A_neg_10_21_port, A_neg_10_20_port, A_neg_10_19_port, 
      A_neg_10_18_port, A_neg_10_17_port, A_neg_10_16_port, A_neg_10_15_port, 
      A_neg_10_14_port, A_neg_10_13_port, A_neg_10_12_port, A_neg_10_11_port, 
      A_neg_9_24_port, A_neg_9_23_port, A_neg_9_22_port, A_neg_9_21_port, 
      A_neg_9_20_port, A_neg_9_19_port, A_neg_9_18_port, A_neg_9_17_port, 
      A_neg_9_16_port, A_neg_9_15_port, A_neg_9_14_port, A_neg_9_13_port, 
      A_neg_9_12_port, A_neg_9_11_port, A_neg_9_10_port, A_neg_8_23_port, 
      A_neg_8_22_port, A_neg_8_21_port, A_neg_8_20_port, A_neg_8_19_port, 
      A_neg_8_18_port, A_neg_8_17_port, A_neg_8_16_port, A_neg_8_15_port, 
      A_neg_8_14_port, A_neg_8_13_port, A_neg_8_12_port, A_neg_8_11_port, 
      A_neg_8_10_port, A_neg_8_9_port, A_neg_7_22_port, A_neg_7_21_port, 
      A_neg_7_20_port, A_neg_7_19_port, A_neg_7_18_port, A_neg_7_17_port, 
      A_neg_7_16_port, A_neg_7_15_port, A_neg_7_14_port, A_neg_7_13_port, 
      A_neg_7_12_port, A_neg_7_11_port, A_neg_7_10_port, A_neg_7_9_port, 
      A_neg_7_8_port, A_neg_6_21_port, A_neg_6_20_port, A_neg_6_19_port, 
      A_neg_6_18_port, A_neg_6_17_port, A_neg_6_16_port, A_neg_6_15_port, 
      A_neg_6_14_port, A_neg_6_13_port, A_neg_6_12_port, A_neg_6_11_port, 
      A_neg_6_10_port, A_neg_6_9_port, A_neg_6_8_port, A_neg_6_7_port, 
      A_neg_5_20_port, A_neg_5_19_port, A_neg_5_18_port, A_neg_5_17_port, 
      A_neg_5_16_port, A_neg_5_15_port, A_neg_5_14_port, A_neg_5_13_port, 
      A_neg_5_12_port, A_neg_5_11_port, A_neg_5_10_port, A_neg_5_9_port, 
      A_neg_5_8_port, A_neg_5_7_port, A_neg_5_6_port, A_neg_4_19_port, 
      A_neg_4_18_port, A_neg_4_17_port, A_neg_4_16_port, A_neg_4_15_port, 
      A_neg_4_14_port, A_neg_4_13_port, A_neg_4_12_port, A_neg_4_11_port, 
      A_neg_4_10_port, A_neg_4_9_port, A_neg_4_8_port, A_neg_4_7_port, 
      A_neg_4_6_port, A_neg_4_5_port, A_neg_3_18_port, A_neg_3_17_port, 
      A_neg_3_16_port, A_neg_3_15_port, A_neg_3_14_port, A_neg_3_13_port, 
      A_neg_3_12_port, A_neg_3_11_port, A_neg_3_10_port, A_neg_3_9_port, 
      A_neg_3_8_port, A_neg_3_7_port, A_neg_3_6_port, A_neg_3_5_port, 
      A_neg_3_4_port, A_neg_2_17_port, A_neg_2_16_port, A_neg_2_15_port, 
      A_neg_2_14_port, A_neg_2_13_port, A_neg_2_12_port, A_neg_2_11_port, 
      A_neg_2_10_port, A_neg_2_9_port, A_neg_2_8_port, A_neg_2_7_port, 
      A_neg_2_6_port, A_neg_2_5_port, A_neg_2_4_port, A_neg_2_3_port, 
      A_neg_1_16_port, A_neg_1_15_port, A_neg_1_14_port, A_neg_1_13_port, 
      A_neg_1_12_port, A_neg_1_11_port, A_neg_1_10_port, A_neg_1_9_port, 
      A_neg_1_8_port, A_neg_1_7_port, A_neg_1_6_port, A_neg_1_5_port, 
      A_neg_1_4_port, A_neg_1_3_port, A_neg_1_2_port, A_neg_0_15_port, 
      A_neg_0_14_port, A_neg_0_13_port, A_neg_0_12_port, A_neg_0_11_port, 
      A_neg_0_10_port, A_neg_0_9_port, A_neg_0_8_port, A_neg_0_7_port, 
      A_neg_0_6_port, A_neg_0_5_port, A_neg_0_4_port, A_neg_0_3_port, 
      A_neg_0_2_port, A_neg_0_1_port, mux_out_7_31_port, mux_out_7_30_port, 
      mux_out_7_29_port, mux_out_7_28_port, mux_out_7_27_port, 
      mux_out_7_26_port, mux_out_7_25_port, mux_out_7_24_port, 
      mux_out_7_23_port, mux_out_7_22_port, mux_out_7_21_port, 
      mux_out_7_20_port, mux_out_7_19_port, mux_out_7_18_port, 
      mux_out_7_17_port, mux_out_7_16_port, mux_out_7_15_port, 
      mux_out_7_14_port, mux_out_7_13_port, mux_out_7_12_port, 
      mux_out_7_11_port, mux_out_7_10_port, mux_out_7_9_port, mux_out_7_8_port,
      mux_out_7_7_port, mux_out_7_6_port, mux_out_7_5_port, mux_out_7_4_port, 
      mux_out_7_3_port, mux_out_7_2_port, mux_out_7_1_port, mux_out_7_0_port, 
      mux_out_6_31_port, mux_out_6_30_port, mux_out_6_29_port, 
      mux_out_6_28_port, mux_out_6_27_port, mux_out_6_26_port, 
      mux_out_6_25_port, mux_out_6_24_port, mux_out_6_23_port, 
      mux_out_6_22_port, mux_out_6_21_port, mux_out_6_20_port, 
      mux_out_6_19_port, mux_out_6_18_port, mux_out_6_17_port, 
      mux_out_6_16_port, mux_out_6_15_port, mux_out_6_14_port, 
      mux_out_6_13_port, mux_out_6_12_port, mux_out_6_11_port, 
      mux_out_6_10_port, mux_out_6_9_port, mux_out_6_8_port, mux_out_6_7_port, 
      mux_out_6_6_port, mux_out_6_5_port, mux_out_6_4_port, mux_out_6_3_port, 
      mux_out_6_2_port, mux_out_6_1_port, mux_out_6_0_port, mux_out_5_31_port, 
      mux_out_5_30_port, mux_out_5_29_port, mux_out_5_28_port, 
      mux_out_5_27_port, mux_out_5_26_port, mux_out_5_25_port, 
      mux_out_5_24_port, mux_out_5_23_port, mux_out_5_22_port, 
      mux_out_5_21_port, mux_out_5_20_port, mux_out_5_19_port, 
      mux_out_5_18_port, mux_out_5_17_port, mux_out_5_16_port, 
      mux_out_5_15_port, mux_out_5_14_port, mux_out_5_13_port, 
      mux_out_5_12_port, mux_out_5_11_port, mux_out_5_10_port, mux_out_5_9_port
      , mux_out_5_8_port, mux_out_5_7_port, mux_out_5_6_port, mux_out_5_5_port,
      mux_out_5_4_port, mux_out_5_3_port, mux_out_5_2_port, mux_out_5_1_port, 
      mux_out_5_0_port, mux_out_4_31_port, mux_out_4_30_port, mux_out_4_29_port
      , mux_out_4_28_port, mux_out_4_27_port, mux_out_4_26_port, 
      mux_out_4_25_port, mux_out_4_24_port, mux_out_4_23_port, 
      mux_out_4_22_port, mux_out_4_21_port, mux_out_4_20_port, 
      mux_out_4_19_port, mux_out_4_18_port, mux_out_4_17_port, 
      mux_out_4_16_port, mux_out_4_15_port, mux_out_4_14_port, 
      mux_out_4_13_port, mux_out_4_12_port, mux_out_4_11_port, 
      mux_out_4_10_port, mux_out_4_9_port, mux_out_4_8_port, mux_out_4_7_port, 
      mux_out_4_6_port, mux_out_4_5_port, mux_out_4_4_port, mux_out_4_3_port, 
      mux_out_4_2_port, mux_out_4_1_port, mux_out_4_0_port, mux_out_3_31_port, 
      mux_out_3_30_port, mux_out_3_29_port, mux_out_3_28_port, 
      mux_out_3_27_port, mux_out_3_26_port, mux_out_3_25_port, 
      mux_out_3_24_port, mux_out_3_23_port, mux_out_3_22_port, 
      mux_out_3_21_port, mux_out_3_20_port, mux_out_3_19_port, 
      mux_out_3_18_port, mux_out_3_17_port, mux_out_3_16_port, 
      mux_out_3_15_port, mux_out_3_14_port, mux_out_3_13_port, 
      mux_out_3_12_port, mux_out_3_11_port, mux_out_3_10_port, mux_out_3_9_port
      , mux_out_3_8_port, mux_out_3_7_port, mux_out_3_6_port, mux_out_3_5_port,
      mux_out_3_4_port, mux_out_3_3_port, mux_out_3_2_port, mux_out_3_1_port, 
      mux_out_3_0_port, mux_out_2_31_port, mux_out_2_30_port, mux_out_2_29_port
      , mux_out_2_28_port, mux_out_2_27_port, mux_out_2_26_port, 
      mux_out_2_25_port, mux_out_2_24_port, mux_out_2_23_port, 
      mux_out_2_22_port, mux_out_2_21_port, mux_out_2_20_port, 
      mux_out_2_19_port, mux_out_2_18_port, mux_out_2_17_port, 
      mux_out_2_16_port, mux_out_2_15_port, mux_out_2_14_port, 
      mux_out_2_13_port, mux_out_2_12_port, mux_out_2_11_port, 
      mux_out_2_10_port, mux_out_2_9_port, mux_out_2_8_port, mux_out_2_7_port, 
      mux_out_2_6_port, mux_out_2_5_port, mux_out_2_4_port, mux_out_2_3_port, 
      mux_out_2_2_port, mux_out_2_1_port, mux_out_2_0_port, addends_7_31_port, 
      addends_7_30_port, addends_7_29_port, addends_7_28_port, 
      addends_7_27_port, addends_7_26_port, addends_7_25_port, 
      addends_7_24_port, addends_7_23_port, addends_7_22_port, 
      addends_7_21_port, addends_7_20_port, addends_7_19_port, 
      addends_7_18_port, addends_7_17_port, addends_7_16_port, 
      addends_7_15_port, addends_7_14_port, addends_7_13_port, 
      addends_7_12_port, addends_7_11_port, addends_7_10_port, addends_7_9_port
      , addends_7_8_port, addends_7_7_port, addends_7_6_port, addends_7_5_port,
      addends_7_4_port, addends_7_3_port, addends_7_2_port, addends_7_1_port, 
      addends_7_0_port, addends_6_31_port, addends_6_30_port, addends_6_29_port
      , addends_6_28_port, addends_6_27_port, addends_6_26_port, 
      addends_6_25_port, addends_6_24_port, addends_6_23_port, 
      addends_6_22_port, addends_6_21_port, addends_6_20_port, 
      addends_6_19_port, addends_6_18_port, addends_6_17_port, 
      addends_6_16_port, addends_6_15_port, addends_6_14_port, 
      addends_6_13_port, addends_6_12_port, addends_6_11_port, 
      addends_6_10_port, addends_6_9_port, addends_6_8_port, addends_6_7_port, 
      addends_6_6_port, addends_6_5_port, addends_6_4_port, addends_6_3_port, 
      addends_6_2_port, addends_6_1_port, addends_6_0_port, addends_5_31_port, 
      addends_5_30_port, addends_5_29_port, addends_5_28_port, 
      addends_5_27_port, addends_5_26_port, addends_5_25_port, 
      addends_5_24_port, addends_5_23_port, addends_5_22_port, 
      addends_5_21_port, addends_5_20_port, addends_5_19_port, 
      addends_5_18_port, addends_5_17_port, addends_5_16_port, 
      addends_5_15_port, addends_5_14_port, addends_5_13_port, 
      addends_5_12_port, addends_5_11_port, addends_5_10_port, addends_5_9_port
      , addends_5_8_port, addends_5_7_port, addends_5_6_port, addends_5_5_port,
      addends_5_4_port, addends_5_3_port, addends_5_2_port, addends_5_1_port, 
      addends_5_0_port, addends_4_31_port, addends_4_30_port, addends_4_29_port
      , addends_4_28_port, addends_4_27_port, addends_4_26_port, 
      addends_4_25_port, addends_4_24_port, addends_4_23_port, 
      addends_4_22_port, addends_4_21_port, addends_4_20_port, 
      addends_4_19_port, addends_4_18_port, addends_4_17_port, 
      addends_4_16_port, addends_4_15_port, addends_4_14_port, 
      addends_4_13_port, addends_4_12_port, addends_4_11_port, 
      addends_4_10_port, addends_4_9_port, addends_4_8_port, addends_4_7_port, 
      addends_4_6_port, addends_4_5_port, addends_4_4_port, addends_4_3_port, 
      addends_4_2_port, addends_4_1_port, addends_4_0_port, addends_3_31_port, 
      addends_3_30_port, addends_3_29_port, addends_3_28_port, 
      addends_3_27_port, addends_3_26_port, addends_3_25_port, 
      addends_3_24_port, addends_3_23_port, addends_3_22_port, 
      addends_3_21_port, addends_3_20_port, addends_3_19_port, 
      addends_3_18_port, addends_3_17_port, addends_3_16_port, 
      addends_3_15_port, addends_3_14_port, addends_3_13_port, 
      addends_3_12_port, addends_3_11_port, addends_3_10_port, addends_3_9_port
      , addends_3_8_port, addends_3_7_port, addends_3_6_port, addends_3_5_port,
      addends_3_4_port, addends_3_3_port, addends_3_2_port, addends_3_1_port, 
      addends_3_0_port, addends_2_31_port, addends_2_30_port, addends_2_29_port
      , addends_2_28_port, addends_2_27_port, addends_2_26_port, 
      addends_2_25_port, addends_2_24_port, addends_2_23_port, 
      addends_2_22_port, addends_2_21_port, addends_2_20_port, 
      addends_2_19_port, addends_2_18_port, addends_2_17_port, 
      addends_2_16_port, addends_2_15_port, addends_2_14_port, 
      addends_2_13_port, addends_2_12_port, addends_2_11_port, 
      addends_2_10_port, addends_2_9_port, addends_2_8_port, addends_2_7_port, 
      addends_2_6_port, addends_2_5_port, addends_2_4_port, addends_2_3_port, 
      addends_2_2_port, addends_2_1_port, addends_2_0_port, addends_1_31_port, 
      addends_1_30_port, addends_1_29_port, addends_1_28_port, 
      addends_1_27_port, addends_1_26_port, addends_1_25_port, 
      addends_1_24_port, addends_1_23_port, addends_1_22_port, 
      addends_1_21_port, addends_1_20_port, addends_1_19_port, 
      addends_1_18_port, addends_1_17_port, addends_1_16_port, 
      addends_1_15_port, addends_1_14_port, addends_1_13_port, 
      addends_1_12_port, addends_1_11_port, addends_1_10_port, addends_1_9_port
      , addends_1_8_port, addends_1_7_port, addends_1_6_port, addends_1_5_port,
      addends_1_4_port, addends_1_3_port, addends_1_2_port, addends_1_1_port, 
      addends_1_0_port, addends_0_31_port, addends_0_30_port, addends_0_29_port
      , addends_0_28_port, addends_0_27_port, addends_0_26_port, 
      addends_0_25_port, addends_0_24_port, addends_0_23_port, 
      addends_0_22_port, addends_0_21_port, addends_0_20_port, 
      addends_0_19_port, addends_0_18_port, addends_0_17_port, 
      addends_0_16_port, addends_0_15_port, addends_0_14_port, 
      addends_0_13_port, addends_0_12_port, addends_0_11_port, 
      addends_0_10_port, addends_0_9_port, addends_0_8_port, addends_0_7_port, 
      addends_0_6_port, addends_0_5_port, addends_0_4_port, addends_0_3_port, 
      addends_0_2_port, addends_0_1_port, addends_0_0_port, pipe1_3_31_port, 
      pipe1_3_30_port, pipe1_3_29_port, pipe1_3_28_port, pipe1_3_27_port, 
      pipe1_3_26_port, pipe1_3_25_port, pipe1_3_24_port, pipe1_3_23_port, 
      pipe1_3_22_port, pipe1_3_21_port, pipe1_3_20_port, pipe1_3_19_port, 
      pipe1_3_18_port, pipe1_3_17_port, pipe1_3_16_port, pipe1_3_15_port, 
      pipe1_3_14_port, pipe1_3_13_port, pipe1_3_12_port, pipe1_3_11_port, 
      pipe1_3_10_port, pipe1_3_9_port, pipe1_3_8_port, pipe1_3_7_port, 
      pipe1_3_6_port, pipe1_3_5_port, pipe1_3_4_port, pipe1_3_3_port, 
      pipe1_3_2_port, pipe1_3_1_port, pipe1_3_0_port, pipe1_2_31_port, 
      pipe1_2_30_port, pipe1_2_29_port, pipe1_2_28_port, pipe1_2_27_port, 
      pipe1_2_26_port, pipe1_2_25_port, pipe1_2_24_port, pipe1_2_23_port, 
      pipe1_2_22_port, pipe1_2_21_port, pipe1_2_20_port, pipe1_2_19_port, 
      pipe1_2_18_port, pipe1_2_17_port, pipe1_2_16_port, pipe1_2_15_port, 
      pipe1_2_14_port, pipe1_2_13_port, pipe1_2_12_port, pipe1_2_11_port, 
      pipe1_2_10_port, pipe1_2_9_port, pipe1_2_8_port, pipe1_2_7_port, 
      pipe1_2_6_port, pipe1_2_5_port, pipe1_2_4_port, pipe1_2_3_port, 
      pipe1_2_2_port, pipe1_2_1_port, pipe1_2_0_port, pipe1_1_31_port, 
      pipe1_1_30_port, pipe1_1_29_port, pipe1_1_28_port, pipe1_1_27_port, 
      pipe1_1_26_port, pipe1_1_25_port, pipe1_1_24_port, pipe1_1_23_port, 
      pipe1_1_22_port, pipe1_1_21_port, pipe1_1_20_port, pipe1_1_19_port, 
      pipe1_1_18_port, pipe1_1_17_port, pipe1_1_16_port, pipe1_1_15_port, 
      pipe1_1_14_port, pipe1_1_13_port, pipe1_1_12_port, pipe1_1_11_port, 
      pipe1_1_10_port, pipe1_1_9_port, pipe1_1_8_port, pipe1_1_7_port, 
      pipe1_1_6_port, pipe1_1_5_port, pipe1_1_4_port, pipe1_1_3_port, 
      pipe1_1_2_port, pipe1_1_1_port, pipe1_1_0_port, pipe1_0_31_port, 
      pipe1_0_30_port, pipe1_0_29_port, pipe1_0_28_port, pipe1_0_27_port, 
      pipe1_0_26_port, pipe1_0_25_port, pipe1_0_24_port, pipe1_0_23_port, 
      pipe1_0_22_port, pipe1_0_21_port, pipe1_0_20_port, pipe1_0_19_port, 
      pipe1_0_18_port, pipe1_0_17_port, pipe1_0_16_port, pipe1_0_15_port, 
      pipe1_0_14_port, pipe1_0_13_port, pipe1_0_12_port, pipe1_0_11_port, 
      pipe1_0_10_port, pipe1_0_9_port, pipe1_0_8_port, pipe1_0_7_port, 
      pipe1_0_6_port, pipe1_0_5_port, pipe1_0_4_port, pipe1_0_3_port, 
      pipe1_0_2_port, pipe1_0_1_port, pipe1_0_0_port, pipe2_1_31_port, 
      pipe2_1_30_port, pipe2_1_29_port, pipe2_1_28_port, pipe2_1_27_port, 
      pipe2_1_26_port, pipe2_1_25_port, pipe2_1_24_port, pipe2_1_23_port, 
      pipe2_1_22_port, pipe2_1_21_port, pipe2_1_20_port, pipe2_1_19_port, 
      pipe2_1_18_port, pipe2_1_17_port, pipe2_1_16_port, pipe2_1_15_port, 
      pipe2_1_14_port, pipe2_1_13_port, pipe2_1_12_port, pipe2_1_11_port, 
      pipe2_1_10_port, pipe2_1_9_port, pipe2_1_8_port, pipe2_1_7_port, 
      pipe2_1_6_port, pipe2_1_5_port, pipe2_1_4_port, pipe2_1_3_port, 
      pipe2_1_2_port, pipe2_1_1_port, pipe2_1_0_port, pipe2_0_31_port, 
      pipe2_0_30_port, pipe2_0_29_port, pipe2_0_28_port, pipe2_0_27_port, 
      pipe2_0_26_port, pipe2_0_25_port, pipe2_0_24_port, pipe2_0_23_port, 
      pipe2_0_22_port, pipe2_0_21_port, pipe2_0_20_port, pipe2_0_19_port, 
      pipe2_0_18_port, pipe2_0_17_port, pipe2_0_16_port, pipe2_0_15_port, 
      pipe2_0_14_port, pipe2_0_13_port, pipe2_0_12_port, pipe2_0_11_port, 
      pipe2_0_10_port, pipe2_0_9_port, pipe2_0_8_port, pipe2_0_7_port, 
      pipe2_0_6_port, pipe2_0_5_port, pipe2_0_4_port, pipe2_0_3_port, 
      pipe2_0_2_port, pipe2_0_1_port, pipe2_0_0_port, selector_23_port, 
      selector_22_port, selector_21_port, selector_20_port, selector_19_port, 
      selector_18_port, selector_17_port, selector_16_port, selector_15_port, 
      selector_14_port, selector_13_port, selector_12_port, selector_11_port, 
      selector_10_port, selector_9_port, selector_8_port, selector_7_port, 
      selector_6_port, selector_5_port, selector_4_port, selector_3_port, 
      selector_2_port, selector_1_port, selector_0_port, reg_in_2_31_port, 
      reg_in_2_30_port, reg_in_2_29_port, reg_in_2_28_port, reg_in_2_27_port, 
      reg_in_2_26_port, reg_in_2_25_port, reg_in_2_24_port, reg_in_2_23_port, 
      reg_in_2_22_port, reg_in_2_21_port, reg_in_2_20_port, reg_in_2_19_port, 
      reg_in_2_18_port, reg_in_2_17_port, reg_in_2_16_port, reg_in_2_15_port, 
      reg_in_2_14_port, reg_in_2_13_port, reg_in_2_12_port, reg_in_2_11_port, 
      reg_in_2_10_port, reg_in_2_9_port, reg_in_2_8_port, reg_in_2_7_port, 
      reg_in_2_6_port, reg_in_2_5_port, reg_in_2_4_port, reg_in_2_3_port, 
      reg_in_2_2_port, reg_in_2_1_port, reg_in_2_0_port, reg_in_1_31_port, 
      reg_in_1_30_port, reg_in_1_29_port, reg_in_1_28_port, reg_in_1_27_port, 
      reg_in_1_26_port, reg_in_1_25_port, reg_in_1_24_port, reg_in_1_23_port, 
      reg_in_1_22_port, reg_in_1_21_port, reg_in_1_20_port, reg_in_1_19_port, 
      reg_in_1_18_port, reg_in_1_17_port, reg_in_1_16_port, reg_in_1_15_port, 
      reg_in_1_14_port, reg_in_1_13_port, reg_in_1_12_port, reg_in_1_11_port, 
      reg_in_1_10_port, reg_in_1_9_port, reg_in_1_8_port, reg_in_1_7_port, 
      reg_in_1_6_port, reg_in_1_5_port, reg_in_1_4_port, reg_in_1_3_port, 
      reg_in_1_2_port, reg_in_1_1_port, reg_in_1_0_port, reg_in_0_31_port, 
      reg_in_0_30_port, reg_in_0_29_port, reg_in_0_28_port, reg_in_0_27_port, 
      reg_in_0_26_port, reg_in_0_25_port, reg_in_0_24_port, reg_in_0_23_port, 
      reg_in_0_22_port, reg_in_0_21_port, reg_in_0_20_port, reg_in_0_19_port, 
      reg_in_0_18_port, reg_in_0_17_port, reg_in_0_16_port, reg_in_0_15_port, 
      reg_in_0_14_port, reg_in_0_13_port, reg_in_0_12_port, reg_in_0_11_port, 
      reg_in_0_10_port, reg_in_0_9_port, reg_in_0_8_port, reg_in_0_7_port, 
      reg_in_0_6_port, reg_in_0_5_port, reg_in_0_4_port, reg_in_0_3_port, 
      reg_in_0_2_port, reg_in_0_1_port, reg_in_0_0_port, reg_out_2_31_port, 
      reg_out_2_30_port, reg_out_2_29_port, reg_out_2_28_port, 
      reg_out_2_27_port, reg_out_2_26_port, reg_out_2_25_port, 
      reg_out_2_24_port, reg_out_2_23_port, reg_out_2_22_port, 
      reg_out_2_21_port, reg_out_2_20_port, reg_out_2_19_port, 
      reg_out_2_18_port, reg_out_2_17_port, reg_out_2_16_port, 
      reg_out_2_15_port, reg_out_2_14_port, reg_out_2_13_port, 
      reg_out_2_12_port, reg_out_2_11_port, reg_out_2_10_port, reg_out_2_9_port
      , reg_out_2_8_port, reg_out_2_7_port, reg_out_2_6_port, reg_out_2_5_port,
      reg_out_2_4_port, reg_out_2_3_port, reg_out_2_2_port, reg_out_2_1_port, 
      reg_out_2_0_port, reg_out_1_31_port, reg_out_1_30_port, reg_out_1_29_port
      , reg_out_1_28_port, reg_out_1_27_port, reg_out_1_26_port, 
      reg_out_1_25_port, reg_out_1_24_port, reg_out_1_23_port, 
      reg_out_1_22_port, reg_out_1_21_port, reg_out_1_20_port, 
      reg_out_1_19_port, reg_out_1_18_port, reg_out_1_17_port, 
      reg_out_1_16_port, reg_out_1_15_port, reg_out_1_14_port, 
      reg_out_1_13_port, reg_out_1_12_port, reg_out_1_11_port, 
      reg_out_1_10_port, reg_out_1_9_port, reg_out_1_8_port, reg_out_1_7_port, 
      reg_out_1_6_port, reg_out_1_5_port, reg_out_1_4_port, reg_out_1_3_port, 
      reg_out_1_2_port, reg_out_1_1_port, reg_out_1_0_port, reg_out_0_31_port, 
      reg_out_0_30_port, reg_out_0_29_port, reg_out_0_28_port, 
      reg_out_0_27_port, reg_out_0_26_port, reg_out_0_25_port, 
      reg_out_0_24_port, reg_out_0_23_port, reg_out_0_22_port, 
      reg_out_0_21_port, reg_out_0_20_port, reg_out_0_19_port, 
      reg_out_0_18_port, reg_out_0_17_port, reg_out_0_16_port, 
      reg_out_0_15_port, reg_out_0_14_port, reg_out_0_13_port, 
      reg_out_0_12_port, reg_out_0_11_port, reg_out_0_10_port, reg_out_0_9_port
      , reg_out_0_8_port, reg_out_0_7_port, reg_out_0_6_port, reg_out_0_5_port,
      reg_out_0_4_port, reg_out_0_3_port, reg_out_0_2_port, reg_out_0_1_port, 
      reg_out_0_0_port, add_out_2_31_port, add_out_2_30_port, add_out_2_29_port
      , add_out_2_28_port, add_out_2_27_port, add_out_2_26_port, 
      add_out_2_25_port, add_out_2_24_port, add_out_2_23_port, 
      add_out_2_22_port, add_out_2_21_port, add_out_2_20_port, 
      add_out_2_19_port, add_out_2_18_port, add_out_2_17_port, 
      add_out_2_16_port, add_out_2_15_port, add_out_2_14_port, 
      add_out_2_13_port, add_out_2_12_port, add_out_2_11_port, 
      add_out_2_10_port, add_out_2_9_port, add_out_2_8_port, add_out_2_7_port, 
      add_out_2_6_port, add_out_2_5_port, add_out_2_4_port, add_out_2_3_port, 
      add_out_2_2_port, add_out_2_1_port, add_out_2_0_port, add_out_1_31_port, 
      add_out_1_30_port, add_out_1_29_port, add_out_1_28_port, 
      add_out_1_27_port, add_out_1_26_port, add_out_1_25_port, 
      add_out_1_24_port, add_out_1_23_port, add_out_1_22_port, 
      add_out_1_21_port, add_out_1_20_port, add_out_1_19_port, 
      add_out_1_18_port, add_out_1_17_port, add_out_1_16_port, 
      add_out_1_15_port, add_out_1_14_port, add_out_1_13_port, 
      add_out_1_12_port, add_out_1_11_port, add_out_1_10_port, add_out_1_9_port
      , add_out_1_8_port, add_out_1_7_port, add_out_1_6_port, add_out_1_5_port,
      add_out_1_4_port, add_out_1_3_port, add_out_1_2_port, add_out_1_1_port, 
      add_out_1_0_port, add_out_0_31_port, add_out_0_30_port, add_out_0_29_port
      , add_out_0_28_port, add_out_0_27_port, add_out_0_26_port, 
      add_out_0_25_port, add_out_0_24_port, add_out_0_23_port, 
      add_out_0_22_port, add_out_0_21_port, add_out_0_20_port, 
      add_out_0_19_port, add_out_0_18_port, add_out_0_17_port, 
      add_out_0_16_port, add_out_0_15_port, add_out_0_14_port, 
      add_out_0_13_port, add_out_0_12_port, add_out_0_11_port, 
      add_out_0_10_port, add_out_0_9_port, add_out_0_8_port, add_out_0_7_port, 
      add_out_0_6_port, add_out_0_5_port, add_out_0_4_port, add_out_0_3_port, 
      add_out_0_2_port, add_out_0_1_port, add_out_0_0_port, 
      sub_126_G16_carry_17_port, sub_126_G16_carry_18_port, 
      sub_126_G16_carry_19_port, sub_126_G16_carry_20_port, 
      sub_126_G16_carry_21_port, sub_126_G16_carry_22_port, 
      sub_126_G16_carry_23_port, sub_126_G16_carry_24_port, 
      sub_126_G16_carry_25_port, sub_126_G16_carry_26_port, 
      sub_126_G16_carry_27_port, sub_126_G16_carry_28_port, 
      sub_126_G16_carry_29_port, sub_126_G16_carry_30_port, 
      sub_126_G15_carry_16_port, sub_126_G15_carry_17_port, 
      sub_126_G15_carry_18_port, sub_126_G15_carry_19_port, 
      sub_126_G15_carry_20_port, sub_126_G15_carry_21_port, 
      sub_126_G15_carry_22_port, sub_126_G15_carry_23_port, 
      sub_126_G15_carry_24_port, sub_126_G15_carry_25_port, 
      sub_126_G15_carry_26_port, sub_126_G15_carry_27_port, 
      sub_126_G15_carry_28_port, sub_126_G15_carry_29_port, 
      sub_126_G14_carry_15_port, sub_126_G14_carry_16_port, 
      sub_126_G14_carry_17_port, sub_126_G14_carry_18_port, 
      sub_126_G14_carry_19_port, sub_126_G14_carry_20_port, 
      sub_126_G14_carry_21_port, sub_126_G14_carry_22_port, 
      sub_126_G14_carry_23_port, sub_126_G14_carry_24_port, 
      sub_126_G14_carry_25_port, sub_126_G14_carry_26_port, 
      sub_126_G14_carry_27_port, sub_126_G14_carry_28_port, 
      sub_126_G13_carry_14_port, sub_126_G13_carry_15_port, 
      sub_126_G13_carry_16_port, sub_126_G13_carry_17_port, 
      sub_126_G13_carry_18_port, sub_126_G13_carry_19_port, 
      sub_126_G13_carry_20_port, sub_126_G13_carry_21_port, 
      sub_126_G13_carry_22_port, sub_126_G13_carry_23_port, 
      sub_126_G13_carry_24_port, sub_126_G13_carry_25_port, 
      sub_126_G13_carry_26_port, sub_126_G13_carry_27_port, 
      sub_126_G12_carry_13_port, sub_126_G12_carry_14_port, 
      sub_126_G12_carry_15_port, sub_126_G12_carry_16_port, 
      sub_126_G12_carry_17_port, sub_126_G12_carry_18_port, 
      sub_126_G12_carry_19_port, sub_126_G12_carry_20_port, 
      sub_126_G12_carry_21_port, sub_126_G12_carry_22_port, 
      sub_126_G12_carry_23_port, sub_126_G12_carry_24_port, 
      sub_126_G12_carry_25_port, sub_126_G12_carry_26_port, 
      sub_126_G11_carry_12_port, sub_126_G11_carry_13_port, 
      sub_126_G11_carry_14_port, sub_126_G11_carry_15_port, 
      sub_126_G11_carry_16_port, sub_126_G11_carry_17_port, 
      sub_126_G11_carry_18_port, sub_126_G11_carry_19_port, 
      sub_126_G11_carry_20_port, sub_126_G11_carry_21_port, 
      sub_126_G11_carry_22_port, sub_126_G11_carry_23_port, 
      sub_126_G11_carry_24_port, sub_126_G11_carry_25_port, 
      sub_126_G10_carry_11_port, sub_126_G10_carry_12_port, 
      sub_126_G10_carry_13_port, sub_126_G10_carry_14_port, 
      sub_126_G10_carry_15_port, sub_126_G10_carry_16_port, 
      sub_126_G10_carry_17_port, sub_126_G10_carry_18_port, 
      sub_126_G10_carry_19_port, sub_126_G10_carry_20_port, 
      sub_126_G10_carry_21_port, sub_126_G10_carry_22_port, 
      sub_126_G10_carry_23_port, sub_126_G10_carry_24_port, 
      sub_126_G9_carry_10_port, sub_126_G9_carry_11_port, 
      sub_126_G9_carry_12_port, sub_126_G9_carry_13_port, 
      sub_126_G9_carry_14_port, sub_126_G9_carry_15_port, 
      sub_126_G9_carry_16_port, sub_126_G9_carry_17_port, 
      sub_126_G9_carry_18_port, sub_126_G9_carry_19_port, 
      sub_126_G9_carry_20_port, sub_126_G9_carry_21_port, 
      sub_126_G9_carry_22_port, sub_126_G9_carry_23_port, 
      sub_126_G8_carry_9_port, sub_126_G8_carry_10_port, 
      sub_126_G8_carry_11_port, sub_126_G8_carry_12_port, 
      sub_126_G8_carry_13_port, sub_126_G8_carry_14_port, 
      sub_126_G8_carry_15_port, sub_126_G8_carry_16_port, 
      sub_126_G8_carry_17_port, sub_126_G8_carry_18_port, 
      sub_126_G8_carry_19_port, sub_126_G8_carry_20_port, 
      sub_126_G8_carry_21_port, sub_126_G8_carry_22_port, 
      sub_126_G7_carry_8_port, sub_126_G7_carry_9_port, 
      sub_126_G7_carry_10_port, sub_126_G7_carry_11_port, 
      sub_126_G7_carry_12_port, sub_126_G7_carry_13_port, 
      sub_126_G7_carry_14_port, sub_126_G7_carry_15_port, 
      sub_126_G7_carry_16_port, sub_126_G7_carry_17_port, 
      sub_126_G7_carry_18_port, sub_126_G7_carry_19_port, 
      sub_126_G7_carry_20_port, sub_126_G7_carry_21_port, 
      sub_126_G6_carry_7_port, sub_126_G6_carry_8_port, sub_126_G6_carry_9_port
      , sub_126_G6_carry_10_port, sub_126_G6_carry_11_port, 
      sub_126_G6_carry_12_port, sub_126_G6_carry_13_port, 
      sub_126_G6_carry_14_port, sub_126_G6_carry_15_port, 
      sub_126_G6_carry_16_port, sub_126_G6_carry_17_port, 
      sub_126_G6_carry_18_port, sub_126_G6_carry_19_port, 
      sub_126_G6_carry_20_port, sub_126_G5_carry_6_port, 
      sub_126_G5_carry_7_port, sub_126_G5_carry_8_port, sub_126_G5_carry_9_port
      , sub_126_G5_carry_10_port, sub_126_G5_carry_11_port, 
      sub_126_G5_carry_12_port, sub_126_G5_carry_13_port, 
      sub_126_G5_carry_14_port, sub_126_G5_carry_15_port, 
      sub_126_G5_carry_16_port, sub_126_G5_carry_17_port, 
      sub_126_G5_carry_18_port, sub_126_G5_carry_19_port, 
      sub_126_G4_carry_5_port, sub_126_G4_carry_6_port, sub_126_G4_carry_7_port
      , sub_126_G4_carry_8_port, sub_126_G4_carry_9_port, 
      sub_126_G4_carry_10_port, sub_126_G4_carry_11_port, 
      sub_126_G4_carry_12_port, sub_126_G4_carry_13_port, 
      sub_126_G4_carry_14_port, sub_126_G4_carry_15_port, 
      sub_126_G4_carry_16_port, sub_126_G4_carry_17_port, 
      sub_126_G4_carry_18_port, sub_126_G3_carry_4_port, 
      sub_126_G3_carry_5_port, sub_126_G3_carry_6_port, sub_126_G3_carry_7_port
      , sub_126_G3_carry_8_port, sub_126_G3_carry_9_port, 
      sub_126_G3_carry_10_port, sub_126_G3_carry_11_port, 
      sub_126_G3_carry_12_port, sub_126_G3_carry_13_port, 
      sub_126_G3_carry_14_port, sub_126_G3_carry_15_port, 
      sub_126_G3_carry_16_port, sub_126_G3_carry_17_port, 
      sub_126_G2_carry_3_port, sub_126_G2_carry_4_port, sub_126_G2_carry_5_port
      , sub_126_G2_carry_6_port, sub_126_G2_carry_7_port, 
      sub_126_G2_carry_8_port, sub_126_G2_carry_9_port, 
      sub_126_G2_carry_10_port, sub_126_G2_carry_11_port, 
      sub_126_G2_carry_12_port, sub_126_G2_carry_13_port, 
      sub_126_G2_carry_14_port, sub_126_G2_carry_15_port, 
      sub_126_G2_carry_16_port, sub_126_carry_2_port, sub_126_carry_3_port, 
      sub_126_carry_4_port, sub_126_carry_5_port, sub_126_carry_6_port, 
      sub_126_carry_7_port, sub_126_carry_8_port, sub_126_carry_9_port, 
      sub_126_carry_10_port, sub_126_carry_11_port, sub_126_carry_12_port, 
      sub_126_carry_13_port, sub_126_carry_14_port, sub_126_carry_15_port, n1, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   addends_reg_3_31_inst : DFF_X1 port map( D => mux_out_3_31_port, CK => CLOCK
                           , Q => addends_3_31_port, QN => n_1314);
   addends_reg_3_30_inst : DFF_X1 port map( D => mux_out_3_30_port, CK => CLOCK
                           , Q => addends_3_30_port, QN => n_1315);
   addends_reg_3_29_inst : DFF_X1 port map( D => mux_out_3_29_port, CK => CLOCK
                           , Q => addends_3_29_port, QN => n_1316);
   addends_reg_3_28_inst : DFF_X1 port map( D => mux_out_3_28_port, CK => CLOCK
                           , Q => addends_3_28_port, QN => n_1317);
   addends_reg_3_27_inst : DFF_X1 port map( D => mux_out_3_27_port, CK => CLOCK
                           , Q => addends_3_27_port, QN => n_1318);
   addends_reg_3_26_inst : DFF_X1 port map( D => mux_out_3_26_port, CK => CLOCK
                           , Q => addends_3_26_port, QN => n_1319);
   addends_reg_3_25_inst : DFF_X1 port map( D => mux_out_3_25_port, CK => CLOCK
                           , Q => addends_3_25_port, QN => n_1320);
   addends_reg_3_24_inst : DFF_X1 port map( D => mux_out_3_24_port, CK => CLOCK
                           , Q => addends_3_24_port, QN => n_1321);
   addends_reg_3_23_inst : DFF_X1 port map( D => mux_out_3_23_port, CK => CLOCK
                           , Q => addends_3_23_port, QN => n_1322);
   addends_reg_3_22_inst : DFF_X1 port map( D => mux_out_3_22_port, CK => CLOCK
                           , Q => addends_3_22_port, QN => n_1323);
   addends_reg_3_21_inst : DFF_X1 port map( D => mux_out_3_21_port, CK => CLOCK
                           , Q => addends_3_21_port, QN => n_1324);
   addends_reg_3_20_inst : DFF_X1 port map( D => mux_out_3_20_port, CK => CLOCK
                           , Q => addends_3_20_port, QN => n_1325);
   addends_reg_3_19_inst : DFF_X1 port map( D => mux_out_3_19_port, CK => CLOCK
                           , Q => addends_3_19_port, QN => n_1326);
   addends_reg_3_18_inst : DFF_X1 port map( D => mux_out_3_18_port, CK => CLOCK
                           , Q => addends_3_18_port, QN => n_1327);
   addends_reg_3_17_inst : DFF_X1 port map( D => mux_out_3_17_port, CK => CLOCK
                           , Q => addends_3_17_port, QN => n_1328);
   addends_reg_3_16_inst : DFF_X1 port map( D => mux_out_3_16_port, CK => CLOCK
                           , Q => addends_3_16_port, QN => n_1329);
   addends_reg_3_15_inst : DFF_X1 port map( D => mux_out_3_15_port, CK => CLOCK
                           , Q => addends_3_15_port, QN => n_1330);
   addends_reg_3_14_inst : DFF_X1 port map( D => mux_out_3_14_port, CK => CLOCK
                           , Q => addends_3_14_port, QN => n_1331);
   addends_reg_3_13_inst : DFF_X1 port map( D => mux_out_3_13_port, CK => CLOCK
                           , Q => addends_3_13_port, QN => n_1332);
   addends_reg_3_12_inst : DFF_X1 port map( D => mux_out_3_12_port, CK => CLOCK
                           , Q => addends_3_12_port, QN => n_1333);
   addends_reg_3_11_inst : DFF_X1 port map( D => mux_out_3_11_port, CK => CLOCK
                           , Q => addends_3_11_port, QN => n_1334);
   addends_reg_3_10_inst : DFF_X1 port map( D => mux_out_3_10_port, CK => CLOCK
                           , Q => addends_3_10_port, QN => n_1335);
   addends_reg_3_9_inst : DFF_X1 port map( D => mux_out_3_9_port, CK => CLOCK, 
                           Q => addends_3_9_port, QN => n_1336);
   addends_reg_3_8_inst : DFF_X1 port map( D => mux_out_3_8_port, CK => CLOCK, 
                           Q => addends_3_8_port, QN => n_1337);
   addends_reg_3_7_inst : DFF_X1 port map( D => mux_out_3_7_port, CK => CLOCK, 
                           Q => addends_3_7_port, QN => n_1338);
   addends_reg_3_6_inst : DFF_X1 port map( D => mux_out_3_6_port, CK => CLOCK, 
                           Q => addends_3_6_port, QN => n_1339);
   addends_reg_3_5_inst : DFF_X1 port map( D => mux_out_3_5_port, CK => CLOCK, 
                           Q => addends_3_5_port, QN => n_1340);
   addends_reg_3_4_inst : DFF_X1 port map( D => mux_out_3_4_port, CK => CLOCK, 
                           Q => addends_3_4_port, QN => n_1341);
   addends_reg_3_3_inst : DFF_X1 port map( D => mux_out_3_3_port, CK => CLOCK, 
                           Q => addends_3_3_port, QN => n_1342);
   addends_reg_3_2_inst : DFF_X1 port map( D => mux_out_3_2_port, CK => CLOCK, 
                           Q => addends_3_2_port, QN => n_1343);
   addends_reg_3_1_inst : DFF_X1 port map( D => mux_out_3_1_port, CK => CLOCK, 
                           Q => addends_3_1_port, QN => n_1344);
   addends_reg_3_0_inst : DFF_X1 port map( D => mux_out_3_0_port, CK => CLOCK, 
                           Q => addends_3_0_port, QN => n_1345);
   addends_reg_2_31_inst : DFF_X1 port map( D => mux_out_2_31_port, CK => CLOCK
                           , Q => addends_2_31_port, QN => n_1346);
   addends_reg_2_30_inst : DFF_X1 port map( D => mux_out_2_30_port, CK => CLOCK
                           , Q => addends_2_30_port, QN => n_1347);
   addends_reg_2_29_inst : DFF_X1 port map( D => mux_out_2_29_port, CK => CLOCK
                           , Q => addends_2_29_port, QN => n_1348);
   addends_reg_2_28_inst : DFF_X1 port map( D => mux_out_2_28_port, CK => CLOCK
                           , Q => addends_2_28_port, QN => n_1349);
   addends_reg_2_27_inst : DFF_X1 port map( D => mux_out_2_27_port, CK => CLOCK
                           , Q => addends_2_27_port, QN => n_1350);
   addends_reg_2_26_inst : DFF_X1 port map( D => mux_out_2_26_port, CK => CLOCK
                           , Q => addends_2_26_port, QN => n_1351);
   addends_reg_2_25_inst : DFF_X1 port map( D => mux_out_2_25_port, CK => CLOCK
                           , Q => addends_2_25_port, QN => n_1352);
   addends_reg_2_24_inst : DFF_X1 port map( D => mux_out_2_24_port, CK => CLOCK
                           , Q => addends_2_24_port, QN => n_1353);
   addends_reg_2_23_inst : DFF_X1 port map( D => mux_out_2_23_port, CK => CLOCK
                           , Q => addends_2_23_port, QN => n_1354);
   addends_reg_2_22_inst : DFF_X1 port map( D => mux_out_2_22_port, CK => CLOCK
                           , Q => addends_2_22_port, QN => n_1355);
   addends_reg_2_21_inst : DFF_X1 port map( D => mux_out_2_21_port, CK => CLOCK
                           , Q => addends_2_21_port, QN => n_1356);
   addends_reg_2_20_inst : DFF_X1 port map( D => mux_out_2_20_port, CK => CLOCK
                           , Q => addends_2_20_port, QN => n_1357);
   addends_reg_2_19_inst : DFF_X1 port map( D => mux_out_2_19_port, CK => CLOCK
                           , Q => addends_2_19_port, QN => n_1358);
   addends_reg_2_18_inst : DFF_X1 port map( D => mux_out_2_18_port, CK => CLOCK
                           , Q => addends_2_18_port, QN => n_1359);
   addends_reg_2_17_inst : DFF_X1 port map( D => mux_out_2_17_port, CK => CLOCK
                           , Q => addends_2_17_port, QN => n_1360);
   addends_reg_2_16_inst : DFF_X1 port map( D => mux_out_2_16_port, CK => CLOCK
                           , Q => addends_2_16_port, QN => n_1361);
   addends_reg_2_15_inst : DFF_X1 port map( D => mux_out_2_15_port, CK => CLOCK
                           , Q => addends_2_15_port, QN => n_1362);
   addends_reg_2_14_inst : DFF_X1 port map( D => mux_out_2_14_port, CK => CLOCK
                           , Q => addends_2_14_port, QN => n_1363);
   addends_reg_2_13_inst : DFF_X1 port map( D => mux_out_2_13_port, CK => CLOCK
                           , Q => addends_2_13_port, QN => n_1364);
   addends_reg_2_12_inst : DFF_X1 port map( D => mux_out_2_12_port, CK => CLOCK
                           , Q => addends_2_12_port, QN => n_1365);
   addends_reg_2_11_inst : DFF_X1 port map( D => mux_out_2_11_port, CK => CLOCK
                           , Q => addends_2_11_port, QN => n_1366);
   addends_reg_2_10_inst : DFF_X1 port map( D => mux_out_2_10_port, CK => CLOCK
                           , Q => addends_2_10_port, QN => n_1367);
   addends_reg_2_9_inst : DFF_X1 port map( D => mux_out_2_9_port, CK => CLOCK, 
                           Q => addends_2_9_port, QN => n_1368);
   addends_reg_2_8_inst : DFF_X1 port map( D => mux_out_2_8_port, CK => CLOCK, 
                           Q => addends_2_8_port, QN => n_1369);
   addends_reg_2_7_inst : DFF_X1 port map( D => mux_out_2_7_port, CK => CLOCK, 
                           Q => addends_2_7_port, QN => n_1370);
   addends_reg_2_6_inst : DFF_X1 port map( D => mux_out_2_6_port, CK => CLOCK, 
                           Q => addends_2_6_port, QN => n_1371);
   addends_reg_2_5_inst : DFF_X1 port map( D => mux_out_2_5_port, CK => CLOCK, 
                           Q => addends_2_5_port, QN => n_1372);
   addends_reg_2_4_inst : DFF_X1 port map( D => mux_out_2_4_port, CK => CLOCK, 
                           Q => addends_2_4_port, QN => n_1373);
   addends_reg_2_3_inst : DFF_X1 port map( D => mux_out_2_3_port, CK => CLOCK, 
                           Q => addends_2_3_port, QN => n_1374);
   addends_reg_2_2_inst : DFF_X1 port map( D => mux_out_2_2_port, CK => CLOCK, 
                           Q => addends_2_2_port, QN => n_1375);
   addends_reg_2_1_inst : DFF_X1 port map( D => mux_out_2_1_port, CK => CLOCK, 
                           Q => addends_2_1_port, QN => n_1376);
   addends_reg_2_0_inst : DFF_X1 port map( D => mux_out_2_0_port, CK => CLOCK, 
                           Q => addends_2_0_port, QN => n_1377);
   pipe1_reg_3_31_inst : DFF_X1 port map( D => mux_out_7_31_port, CK => CLOCK, 
                           Q => pipe1_3_31_port, QN => n_1378);
   pipe1_reg_3_30_inst : DFF_X1 port map( D => mux_out_7_30_port, CK => CLOCK, 
                           Q => pipe1_3_30_port, QN => n_1379);
   pipe1_reg_3_29_inst : DFF_X1 port map( D => mux_out_7_29_port, CK => CLOCK, 
                           Q => pipe1_3_29_port, QN => n_1380);
   pipe1_reg_3_28_inst : DFF_X1 port map( D => mux_out_7_28_port, CK => CLOCK, 
                           Q => pipe1_3_28_port, QN => n_1381);
   pipe1_reg_3_27_inst : DFF_X1 port map( D => mux_out_7_27_port, CK => CLOCK, 
                           Q => pipe1_3_27_port, QN => n_1382);
   pipe1_reg_3_26_inst : DFF_X1 port map( D => mux_out_7_26_port, CK => CLOCK, 
                           Q => pipe1_3_26_port, QN => n_1383);
   pipe1_reg_3_25_inst : DFF_X1 port map( D => mux_out_7_25_port, CK => CLOCK, 
                           Q => pipe1_3_25_port, QN => n_1384);
   pipe1_reg_3_24_inst : DFF_X1 port map( D => mux_out_7_24_port, CK => CLOCK, 
                           Q => pipe1_3_24_port, QN => n_1385);
   pipe1_reg_3_23_inst : DFF_X1 port map( D => mux_out_7_23_port, CK => CLOCK, 
                           Q => pipe1_3_23_port, QN => n_1386);
   pipe1_reg_3_22_inst : DFF_X1 port map( D => mux_out_7_22_port, CK => CLOCK, 
                           Q => pipe1_3_22_port, QN => n_1387);
   pipe1_reg_3_21_inst : DFF_X1 port map( D => mux_out_7_21_port, CK => CLOCK, 
                           Q => pipe1_3_21_port, QN => n_1388);
   pipe1_reg_3_20_inst : DFF_X1 port map( D => mux_out_7_20_port, CK => CLOCK, 
                           Q => pipe1_3_20_port, QN => n_1389);
   pipe1_reg_3_19_inst : DFF_X1 port map( D => mux_out_7_19_port, CK => CLOCK, 
                           Q => pipe1_3_19_port, QN => n_1390);
   pipe1_reg_3_18_inst : DFF_X1 port map( D => mux_out_7_18_port, CK => CLOCK, 
                           Q => pipe1_3_18_port, QN => n_1391);
   pipe1_reg_3_17_inst : DFF_X1 port map( D => mux_out_7_17_port, CK => CLOCK, 
                           Q => pipe1_3_17_port, QN => n_1392);
   pipe1_reg_3_16_inst : DFF_X1 port map( D => mux_out_7_16_port, CK => CLOCK, 
                           Q => pipe1_3_16_port, QN => n_1393);
   pipe1_reg_3_15_inst : DFF_X1 port map( D => mux_out_7_15_port, CK => CLOCK, 
                           Q => pipe1_3_15_port, QN => n_1394);
   pipe1_reg_3_14_inst : DFF_X1 port map( D => mux_out_7_14_port, CK => CLOCK, 
                           Q => pipe1_3_14_port, QN => n_1395);
   pipe1_reg_3_13_inst : DFF_X1 port map( D => mux_out_7_13_port, CK => CLOCK, 
                           Q => pipe1_3_13_port, QN => n_1396);
   pipe1_reg_3_12_inst : DFF_X1 port map( D => mux_out_7_12_port, CK => CLOCK, 
                           Q => pipe1_3_12_port, QN => n_1397);
   pipe1_reg_3_11_inst : DFF_X1 port map( D => mux_out_7_11_port, CK => CLOCK, 
                           Q => pipe1_3_11_port, QN => n_1398);
   pipe1_reg_3_10_inst : DFF_X1 port map( D => mux_out_7_10_port, CK => CLOCK, 
                           Q => pipe1_3_10_port, QN => n_1399);
   pipe1_reg_3_9_inst : DFF_X1 port map( D => mux_out_7_9_port, CK => CLOCK, Q 
                           => pipe1_3_9_port, QN => n_1400);
   pipe1_reg_3_8_inst : DFF_X1 port map( D => mux_out_7_8_port, CK => CLOCK, Q 
                           => pipe1_3_8_port, QN => n_1401);
   pipe1_reg_3_7_inst : DFF_X1 port map( D => mux_out_7_7_port, CK => CLOCK, Q 
                           => pipe1_3_7_port, QN => n_1402);
   pipe1_reg_3_6_inst : DFF_X1 port map( D => mux_out_7_6_port, CK => CLOCK, Q 
                           => pipe1_3_6_port, QN => n_1403);
   pipe1_reg_3_5_inst : DFF_X1 port map( D => mux_out_7_5_port, CK => CLOCK, Q 
                           => pipe1_3_5_port, QN => n_1404);
   pipe1_reg_3_4_inst : DFF_X1 port map( D => mux_out_7_4_port, CK => CLOCK, Q 
                           => pipe1_3_4_port, QN => n_1405);
   pipe1_reg_3_3_inst : DFF_X1 port map( D => mux_out_7_3_port, CK => CLOCK, Q 
                           => pipe1_3_3_port, QN => n_1406);
   pipe1_reg_3_2_inst : DFF_X1 port map( D => mux_out_7_2_port, CK => CLOCK, Q 
                           => pipe1_3_2_port, QN => n_1407);
   pipe1_reg_3_1_inst : DFF_X1 port map( D => mux_out_7_1_port, CK => CLOCK, Q 
                           => pipe1_3_1_port, QN => n_1408);
   pipe1_reg_3_0_inst : DFF_X1 port map( D => mux_out_7_0_port, CK => CLOCK, Q 
                           => pipe1_3_0_port, QN => n_1409);
   pipe1_reg_2_31_inst : DFF_X1 port map( D => mux_out_6_31_port, CK => CLOCK, 
                           Q => pipe1_2_31_port, QN => n_1410);
   pipe1_reg_2_30_inst : DFF_X1 port map( D => mux_out_6_30_port, CK => CLOCK, 
                           Q => pipe1_2_30_port, QN => n_1411);
   pipe1_reg_2_29_inst : DFF_X1 port map( D => mux_out_6_29_port, CK => CLOCK, 
                           Q => pipe1_2_29_port, QN => n_1412);
   pipe1_reg_2_28_inst : DFF_X1 port map( D => mux_out_6_28_port, CK => CLOCK, 
                           Q => pipe1_2_28_port, QN => n_1413);
   pipe1_reg_2_27_inst : DFF_X1 port map( D => mux_out_6_27_port, CK => CLOCK, 
                           Q => pipe1_2_27_port, QN => n_1414);
   pipe1_reg_2_26_inst : DFF_X1 port map( D => mux_out_6_26_port, CK => CLOCK, 
                           Q => pipe1_2_26_port, QN => n_1415);
   pipe1_reg_2_25_inst : DFF_X1 port map( D => mux_out_6_25_port, CK => CLOCK, 
                           Q => pipe1_2_25_port, QN => n_1416);
   pipe1_reg_2_24_inst : DFF_X1 port map( D => mux_out_6_24_port, CK => CLOCK, 
                           Q => pipe1_2_24_port, QN => n_1417);
   pipe1_reg_2_23_inst : DFF_X1 port map( D => mux_out_6_23_port, CK => CLOCK, 
                           Q => pipe1_2_23_port, QN => n_1418);
   pipe1_reg_2_22_inst : DFF_X1 port map( D => mux_out_6_22_port, CK => CLOCK, 
                           Q => pipe1_2_22_port, QN => n_1419);
   pipe1_reg_2_21_inst : DFF_X1 port map( D => mux_out_6_21_port, CK => CLOCK, 
                           Q => pipe1_2_21_port, QN => n_1420);
   pipe1_reg_2_20_inst : DFF_X1 port map( D => mux_out_6_20_port, CK => CLOCK, 
                           Q => pipe1_2_20_port, QN => n_1421);
   pipe1_reg_2_19_inst : DFF_X1 port map( D => mux_out_6_19_port, CK => CLOCK, 
                           Q => pipe1_2_19_port, QN => n_1422);
   pipe1_reg_2_18_inst : DFF_X1 port map( D => mux_out_6_18_port, CK => CLOCK, 
                           Q => pipe1_2_18_port, QN => n_1423);
   pipe1_reg_2_17_inst : DFF_X1 port map( D => mux_out_6_17_port, CK => CLOCK, 
                           Q => pipe1_2_17_port, QN => n_1424);
   pipe1_reg_2_16_inst : DFF_X1 port map( D => mux_out_6_16_port, CK => CLOCK, 
                           Q => pipe1_2_16_port, QN => n_1425);
   pipe1_reg_2_15_inst : DFF_X1 port map( D => mux_out_6_15_port, CK => CLOCK, 
                           Q => pipe1_2_15_port, QN => n_1426);
   pipe1_reg_2_14_inst : DFF_X1 port map( D => mux_out_6_14_port, CK => CLOCK, 
                           Q => pipe1_2_14_port, QN => n_1427);
   pipe1_reg_2_13_inst : DFF_X1 port map( D => mux_out_6_13_port, CK => CLOCK, 
                           Q => pipe1_2_13_port, QN => n_1428);
   pipe1_reg_2_12_inst : DFF_X1 port map( D => mux_out_6_12_port, CK => CLOCK, 
                           Q => pipe1_2_12_port, QN => n_1429);
   pipe1_reg_2_11_inst : DFF_X1 port map( D => mux_out_6_11_port, CK => CLOCK, 
                           Q => pipe1_2_11_port, QN => n_1430);
   pipe1_reg_2_10_inst : DFF_X1 port map( D => mux_out_6_10_port, CK => CLOCK, 
                           Q => pipe1_2_10_port, QN => n_1431);
   pipe1_reg_2_9_inst : DFF_X1 port map( D => mux_out_6_9_port, CK => CLOCK, Q 
                           => pipe1_2_9_port, QN => n_1432);
   pipe1_reg_2_8_inst : DFF_X1 port map( D => mux_out_6_8_port, CK => CLOCK, Q 
                           => pipe1_2_8_port, QN => n_1433);
   pipe1_reg_2_7_inst : DFF_X1 port map( D => mux_out_6_7_port, CK => CLOCK, Q 
                           => pipe1_2_7_port, QN => n_1434);
   pipe1_reg_2_6_inst : DFF_X1 port map( D => mux_out_6_6_port, CK => CLOCK, Q 
                           => pipe1_2_6_port, QN => n_1435);
   pipe1_reg_2_5_inst : DFF_X1 port map( D => mux_out_6_5_port, CK => CLOCK, Q 
                           => pipe1_2_5_port, QN => n_1436);
   pipe1_reg_2_4_inst : DFF_X1 port map( D => mux_out_6_4_port, CK => CLOCK, Q 
                           => pipe1_2_4_port, QN => n_1437);
   pipe1_reg_2_3_inst : DFF_X1 port map( D => mux_out_6_3_port, CK => CLOCK, Q 
                           => pipe1_2_3_port, QN => n_1438);
   pipe1_reg_2_2_inst : DFF_X1 port map( D => mux_out_6_2_port, CK => CLOCK, Q 
                           => pipe1_2_2_port, QN => n_1439);
   pipe1_reg_2_1_inst : DFF_X1 port map( D => mux_out_6_1_port, CK => CLOCK, Q 
                           => pipe1_2_1_port, QN => n_1440);
   pipe1_reg_2_0_inst : DFF_X1 port map( D => mux_out_6_0_port, CK => CLOCK, Q 
                           => pipe1_2_0_port, QN => n_1441);
   pipe1_reg_1_31_inst : DFF_X1 port map( D => mux_out_5_31_port, CK => CLOCK, 
                           Q => pipe1_1_31_port, QN => n_1442);
   pipe1_reg_1_30_inst : DFF_X1 port map( D => mux_out_5_30_port, CK => CLOCK, 
                           Q => pipe1_1_30_port, QN => n_1443);
   pipe1_reg_1_29_inst : DFF_X1 port map( D => mux_out_5_29_port, CK => CLOCK, 
                           Q => pipe1_1_29_port, QN => n_1444);
   pipe1_reg_1_28_inst : DFF_X1 port map( D => mux_out_5_28_port, CK => CLOCK, 
                           Q => pipe1_1_28_port, QN => n_1445);
   addends_reg_5_28_inst : DFF_X1 port map( D => pipe1_1_28_port, CK => CLOCK, 
                           Q => addends_5_28_port, QN => n_1446);
   pipe1_reg_1_27_inst : DFF_X1 port map( D => mux_out_5_27_port, CK => CLOCK, 
                           Q => pipe1_1_27_port, QN => n_1447);
   addends_reg_5_27_inst : DFF_X1 port map( D => pipe1_1_27_port, CK => CLOCK, 
                           Q => addends_5_27_port, QN => n_1448);
   pipe1_reg_1_26_inst : DFF_X1 port map( D => mux_out_5_26_port, CK => CLOCK, 
                           Q => pipe1_1_26_port, QN => n_1449);
   addends_reg_5_26_inst : DFF_X1 port map( D => pipe1_1_26_port, CK => CLOCK, 
                           Q => addends_5_26_port, QN => n_1450);
   pipe1_reg_1_25_inst : DFF_X1 port map( D => mux_out_5_25_port, CK => CLOCK, 
                           Q => pipe1_1_25_port, QN => n_1451);
   addends_reg_5_25_inst : DFF_X1 port map( D => pipe1_1_25_port, CK => CLOCK, 
                           Q => addends_5_25_port, QN => n_1452);
   pipe1_reg_1_24_inst : DFF_X1 port map( D => mux_out_5_24_port, CK => CLOCK, 
                           Q => pipe1_1_24_port, QN => n_1453);
   addends_reg_5_24_inst : DFF_X1 port map( D => pipe1_1_24_port, CK => CLOCK, 
                           Q => addends_5_24_port, QN => n_1454);
   pipe1_reg_1_23_inst : DFF_X1 port map( D => mux_out_5_23_port, CK => CLOCK, 
                           Q => pipe1_1_23_port, QN => n_1455);
   addends_reg_5_23_inst : DFF_X1 port map( D => pipe1_1_23_port, CK => CLOCK, 
                           Q => addends_5_23_port, QN => n_1456);
   pipe1_reg_1_22_inst : DFF_X1 port map( D => mux_out_5_22_port, CK => CLOCK, 
                           Q => pipe1_1_22_port, QN => n_1457);
   addends_reg_5_22_inst : DFF_X1 port map( D => pipe1_1_22_port, CK => CLOCK, 
                           Q => addends_5_22_port, QN => n_1458);
   pipe1_reg_1_21_inst : DFF_X1 port map( D => mux_out_5_21_port, CK => CLOCK, 
                           Q => pipe1_1_21_port, QN => n_1459);
   addends_reg_5_21_inst : DFF_X1 port map( D => pipe1_1_21_port, CK => CLOCK, 
                           Q => addends_5_21_port, QN => n_1460);
   pipe1_reg_1_20_inst : DFF_X1 port map( D => mux_out_5_20_port, CK => CLOCK, 
                           Q => pipe1_1_20_port, QN => n_1461);
   addends_reg_5_20_inst : DFF_X1 port map( D => pipe1_1_20_port, CK => CLOCK, 
                           Q => addends_5_20_port, QN => n_1462);
   pipe1_reg_1_19_inst : DFF_X1 port map( D => mux_out_5_19_port, CK => CLOCK, 
                           Q => pipe1_1_19_port, QN => n_1463);
   addends_reg_5_19_inst : DFF_X1 port map( D => pipe1_1_19_port, CK => CLOCK, 
                           Q => addends_5_19_port, QN => n_1464);
   pipe1_reg_1_18_inst : DFF_X1 port map( D => mux_out_5_18_port, CK => CLOCK, 
                           Q => pipe1_1_18_port, QN => n_1465);
   addends_reg_5_18_inst : DFF_X1 port map( D => pipe1_1_18_port, CK => CLOCK, 
                           Q => addends_5_18_port, QN => n_1466);
   pipe1_reg_1_17_inst : DFF_X1 port map( D => mux_out_5_17_port, CK => CLOCK, 
                           Q => pipe1_1_17_port, QN => n_1467);
   addends_reg_5_17_inst : DFF_X1 port map( D => pipe1_1_17_port, CK => CLOCK, 
                           Q => addends_5_17_port, QN => n_1468);
   pipe1_reg_1_16_inst : DFF_X1 port map( D => mux_out_5_16_port, CK => CLOCK, 
                           Q => pipe1_1_16_port, QN => n_1469);
   addends_reg_5_16_inst : DFF_X1 port map( D => pipe1_1_16_port, CK => CLOCK, 
                           Q => addends_5_16_port, QN => n_1470);
   pipe1_reg_1_15_inst : DFF_X1 port map( D => mux_out_5_15_port, CK => CLOCK, 
                           Q => pipe1_1_15_port, QN => n_1471);
   addends_reg_5_15_inst : DFF_X1 port map( D => pipe1_1_15_port, CK => CLOCK, 
                           Q => addends_5_15_port, QN => n_1472);
   pipe1_reg_1_14_inst : DFF_X1 port map( D => mux_out_5_14_port, CK => CLOCK, 
                           Q => pipe1_1_14_port, QN => n_1473);
   addends_reg_5_14_inst : DFF_X1 port map( D => pipe1_1_14_port, CK => CLOCK, 
                           Q => addends_5_14_port, QN => n_1474);
   pipe1_reg_1_13_inst : DFF_X1 port map( D => mux_out_5_13_port, CK => CLOCK, 
                           Q => pipe1_1_13_port, QN => n_1475);
   addends_reg_5_13_inst : DFF_X1 port map( D => pipe1_1_13_port, CK => CLOCK, 
                           Q => addends_5_13_port, QN => n_1476);
   pipe1_reg_1_12_inst : DFF_X1 port map( D => mux_out_5_12_port, CK => CLOCK, 
                           Q => pipe1_1_12_port, QN => n_1477);
   addends_reg_5_12_inst : DFF_X1 port map( D => pipe1_1_12_port, CK => CLOCK, 
                           Q => addends_5_12_port, QN => n_1478);
   pipe1_reg_1_11_inst : DFF_X1 port map( D => mux_out_5_11_port, CK => CLOCK, 
                           Q => pipe1_1_11_port, QN => n_1479);
   addends_reg_5_11_inst : DFF_X1 port map( D => pipe1_1_11_port, CK => CLOCK, 
                           Q => addends_5_11_port, QN => n_1480);
   pipe1_reg_1_10_inst : DFF_X1 port map( D => mux_out_5_10_port, CK => CLOCK, 
                           Q => pipe1_1_10_port, QN => n_1481);
   addends_reg_5_10_inst : DFF_X1 port map( D => pipe1_1_10_port, CK => CLOCK, 
                           Q => addends_5_10_port, QN => n_1482);
   pipe1_reg_1_9_inst : DFF_X1 port map( D => mux_out_5_9_port, CK => CLOCK, Q 
                           => pipe1_1_9_port, QN => n_1483);
   addends_reg_5_9_inst : DFF_X1 port map( D => pipe1_1_9_port, CK => CLOCK, Q 
                           => addends_5_9_port, QN => n_1484);
   pipe1_reg_1_8_inst : DFF_X1 port map( D => mux_out_5_8_port, CK => CLOCK, Q 
                           => pipe1_1_8_port, QN => n_1485);
   addends_reg_5_8_inst : DFF_X1 port map( D => pipe1_1_8_port, CK => CLOCK, Q 
                           => addends_5_8_port, QN => n_1486);
   pipe1_reg_1_7_inst : DFF_X1 port map( D => mux_out_5_7_port, CK => CLOCK, Q 
                           => pipe1_1_7_port, QN => n_1487);
   addends_reg_5_7_inst : DFF_X1 port map( D => pipe1_1_7_port, CK => CLOCK, Q 
                           => addends_5_7_port, QN => n_1488);
   pipe1_reg_1_6_inst : DFF_X1 port map( D => mux_out_5_6_port, CK => CLOCK, Q 
                           => pipe1_1_6_port, QN => n_1489);
   addends_reg_5_6_inst : DFF_X1 port map( D => pipe1_1_6_port, CK => CLOCK, Q 
                           => addends_5_6_port, QN => n_1490);
   pipe1_reg_1_5_inst : DFF_X1 port map( D => mux_out_5_5_port, CK => CLOCK, Q 
                           => pipe1_1_5_port, QN => n_1491);
   addends_reg_5_5_inst : DFF_X1 port map( D => pipe1_1_5_port, CK => CLOCK, Q 
                           => addends_5_5_port, QN => n_1492);
   pipe1_reg_1_4_inst : DFF_X1 port map( D => mux_out_5_4_port, CK => CLOCK, Q 
                           => pipe1_1_4_port, QN => n_1493);
   pipe1_reg_1_3_inst : DFF_X1 port map( D => mux_out_5_3_port, CK => CLOCK, Q 
                           => pipe1_1_3_port, QN => n_1494);
   addends_reg_5_3_inst : DFF_X1 port map( D => pipe1_1_3_port, CK => CLOCK, Q 
                           => addends_5_3_port, QN => n_1495);
   pipe1_reg_1_2_inst : DFF_X1 port map( D => mux_out_5_2_port, CK => CLOCK, Q 
                           => pipe1_1_2_port, QN => n_1496);
   addends_reg_5_2_inst : DFF_X1 port map( D => pipe1_1_2_port, CK => CLOCK, Q 
                           => addends_5_2_port, QN => n_1497);
   pipe1_reg_1_1_inst : DFF_X1 port map( D => mux_out_5_1_port, CK => CLOCK, Q 
                           => pipe1_1_1_port, QN => n_1498);
   addends_reg_5_1_inst : DFF_X1 port map( D => pipe1_1_1_port, CK => CLOCK, Q 
                           => addends_5_1_port, QN => n_1499);
   pipe1_reg_1_0_inst : DFF_X1 port map( D => mux_out_5_0_port, CK => CLOCK, Q 
                           => pipe1_1_0_port, QN => n_1500);
   addends_reg_5_0_inst : DFF_X1 port map( D => pipe1_1_0_port, CK => CLOCK, Q 
                           => addends_5_0_port, QN => n_1501);
   pipe1_reg_0_31_inst : DFF_X1 port map( D => mux_out_4_31_port, CK => CLOCK, 
                           Q => pipe1_0_31_port, QN => n_1502);
   addends_reg_4_31_inst : DFF_X1 port map( D => pipe1_0_31_port, CK => CLOCK, 
                           Q => addends_4_31_port, QN => n_1503);
   pipe1_reg_0_30_inst : DFF_X1 port map( D => mux_out_4_30_port, CK => CLOCK, 
                           Q => pipe1_0_30_port, QN => n_1504);
   pipe1_reg_0_29_inst : DFF_X1 port map( D => mux_out_4_29_port, CK => CLOCK, 
                           Q => pipe1_0_29_port, QN => n_1505);
   addends_reg_4_29_inst : DFF_X1 port map( D => pipe1_0_29_port, CK => CLOCK, 
                           Q => addends_4_29_port, QN => n_1506);
   pipe1_reg_0_28_inst : DFF_X1 port map( D => mux_out_4_28_port, CK => CLOCK, 
                           Q => pipe1_0_28_port, QN => n_1507);
   addends_reg_4_28_inst : DFF_X1 port map( D => pipe1_0_28_port, CK => CLOCK, 
                           Q => addends_4_28_port, QN => n_1508);
   pipe1_reg_0_27_inst : DFF_X1 port map( D => mux_out_4_27_port, CK => CLOCK, 
                           Q => pipe1_0_27_port, QN => n_1509);
   addends_reg_4_27_inst : DFF_X1 port map( D => pipe1_0_27_port, CK => CLOCK, 
                           Q => addends_4_27_port, QN => n_1510);
   pipe1_reg_0_26_inst : DFF_X1 port map( D => mux_out_4_26_port, CK => CLOCK, 
                           Q => pipe1_0_26_port, QN => n_1511);
   addends_reg_4_26_inst : DFF_X1 port map( D => pipe1_0_26_port, CK => CLOCK, 
                           Q => addends_4_26_port, QN => n_1512);
   pipe1_reg_0_25_inst : DFF_X1 port map( D => mux_out_4_25_port, CK => CLOCK, 
                           Q => pipe1_0_25_port, QN => n_1513);
   addends_reg_4_25_inst : DFF_X1 port map( D => pipe1_0_25_port, CK => CLOCK, 
                           Q => addends_4_25_port, QN => n_1514);
   pipe1_reg_0_24_inst : DFF_X1 port map( D => mux_out_4_24_port, CK => CLOCK, 
                           Q => pipe1_0_24_port, QN => n_1515);
   addends_reg_4_24_inst : DFF_X1 port map( D => pipe1_0_24_port, CK => CLOCK, 
                           Q => addends_4_24_port, QN => n_1516);
   pipe1_reg_0_23_inst : DFF_X1 port map( D => mux_out_4_23_port, CK => CLOCK, 
                           Q => pipe1_0_23_port, QN => n_1517);
   addends_reg_4_23_inst : DFF_X1 port map( D => pipe1_0_23_port, CK => CLOCK, 
                           Q => addends_4_23_port, QN => n_1518);
   pipe1_reg_0_22_inst : DFF_X1 port map( D => mux_out_4_22_port, CK => CLOCK, 
                           Q => pipe1_0_22_port, QN => n_1519);
   addends_reg_4_22_inst : DFF_X1 port map( D => pipe1_0_22_port, CK => CLOCK, 
                           Q => addends_4_22_port, QN => n_1520);
   pipe1_reg_0_21_inst : DFF_X1 port map( D => mux_out_4_21_port, CK => CLOCK, 
                           Q => pipe1_0_21_port, QN => n_1521);
   addends_reg_4_21_inst : DFF_X1 port map( D => pipe1_0_21_port, CK => CLOCK, 
                           Q => addends_4_21_port, QN => n_1522);
   pipe1_reg_0_20_inst : DFF_X1 port map( D => mux_out_4_20_port, CK => CLOCK, 
                           Q => pipe1_0_20_port, QN => n_1523);
   addends_reg_4_20_inst : DFF_X1 port map( D => pipe1_0_20_port, CK => CLOCK, 
                           Q => addends_4_20_port, QN => n_1524);
   pipe1_reg_0_19_inst : DFF_X1 port map( D => mux_out_4_19_port, CK => CLOCK, 
                           Q => pipe1_0_19_port, QN => n_1525);
   addends_reg_4_19_inst : DFF_X1 port map( D => pipe1_0_19_port, CK => CLOCK, 
                           Q => addends_4_19_port, QN => n_1526);
   pipe1_reg_0_18_inst : DFF_X1 port map( D => mux_out_4_18_port, CK => CLOCK, 
                           Q => pipe1_0_18_port, QN => n_1527);
   addends_reg_4_18_inst : DFF_X1 port map( D => pipe1_0_18_port, CK => CLOCK, 
                           Q => addends_4_18_port, QN => n_1528);
   pipe1_reg_0_17_inst : DFF_X1 port map( D => mux_out_4_17_port, CK => CLOCK, 
                           Q => pipe1_0_17_port, QN => n_1529);
   addends_reg_4_17_inst : DFF_X1 port map( D => pipe1_0_17_port, CK => CLOCK, 
                           Q => addends_4_17_port, QN => n_1530);
   pipe1_reg_0_16_inst : DFF_X1 port map( D => mux_out_4_16_port, CK => CLOCK, 
                           Q => pipe1_0_16_port, QN => n_1531);
   addends_reg_4_16_inst : DFF_X1 port map( D => pipe1_0_16_port, CK => CLOCK, 
                           Q => addends_4_16_port, QN => n_1532);
   pipe1_reg_0_15_inst : DFF_X1 port map( D => mux_out_4_15_port, CK => CLOCK, 
                           Q => pipe1_0_15_port, QN => n_1533);
   addends_reg_4_15_inst : DFF_X1 port map( D => pipe1_0_15_port, CK => CLOCK, 
                           Q => addends_4_15_port, QN => n_1534);
   pipe1_reg_0_14_inst : DFF_X1 port map( D => mux_out_4_14_port, CK => CLOCK, 
                           Q => pipe1_0_14_port, QN => n_1535);
   addends_reg_4_14_inst : DFF_X1 port map( D => pipe1_0_14_port, CK => CLOCK, 
                           Q => addends_4_14_port, QN => n_1536);
   pipe1_reg_0_13_inst : DFF_X1 port map( D => mux_out_4_13_port, CK => CLOCK, 
                           Q => pipe1_0_13_port, QN => n_1537);
   addends_reg_4_13_inst : DFF_X1 port map( D => pipe1_0_13_port, CK => CLOCK, 
                           Q => addends_4_13_port, QN => n_1538);
   pipe1_reg_0_12_inst : DFF_X1 port map( D => mux_out_4_12_port, CK => CLOCK, 
                           Q => pipe1_0_12_port, QN => n_1539);
   addends_reg_4_12_inst : DFF_X1 port map( D => pipe1_0_12_port, CK => CLOCK, 
                           Q => addends_4_12_port, QN => n_1540);
   pipe1_reg_0_11_inst : DFF_X1 port map( D => mux_out_4_11_port, CK => CLOCK, 
                           Q => pipe1_0_11_port, QN => n_1541);
   addends_reg_4_11_inst : DFF_X1 port map( D => pipe1_0_11_port, CK => CLOCK, 
                           Q => addends_4_11_port, QN => n_1542);
   pipe1_reg_0_10_inst : DFF_X1 port map( D => mux_out_4_10_port, CK => CLOCK, 
                           Q => pipe1_0_10_port, QN => n_1543);
   addends_reg_4_10_inst : DFF_X1 port map( D => pipe1_0_10_port, CK => CLOCK, 
                           Q => addends_4_10_port, QN => n_1544);
   pipe1_reg_0_9_inst : DFF_X1 port map( D => mux_out_4_9_port, CK => CLOCK, Q 
                           => pipe1_0_9_port, QN => n_1545);
   addends_reg_4_9_inst : DFF_X1 port map( D => pipe1_0_9_port, CK => CLOCK, Q 
                           => addends_4_9_port, QN => n_1546);
   pipe1_reg_0_8_inst : DFF_X1 port map( D => mux_out_4_8_port, CK => CLOCK, Q 
                           => pipe1_0_8_port, QN => n_1547);
   addends_reg_4_8_inst : DFF_X1 port map( D => pipe1_0_8_port, CK => CLOCK, Q 
                           => addends_4_8_port, QN => n_1548);
   pipe1_reg_0_7_inst : DFF_X1 port map( D => mux_out_4_7_port, CK => CLOCK, Q 
                           => pipe1_0_7_port, QN => n_1549);
   addends_reg_4_7_inst : DFF_X1 port map( D => pipe1_0_7_port, CK => CLOCK, Q 
                           => addends_4_7_port, QN => n_1550);
   pipe1_reg_0_6_inst : DFF_X1 port map( D => mux_out_4_6_port, CK => CLOCK, Q 
                           => pipe1_0_6_port, QN => n_1551);
   addends_reg_4_6_inst : DFF_X1 port map( D => pipe1_0_6_port, CK => CLOCK, Q 
                           => addends_4_6_port, QN => n_1552);
   pipe1_reg_0_5_inst : DFF_X1 port map( D => mux_out_4_5_port, CK => CLOCK, Q 
                           => pipe1_0_5_port, QN => n_1553);
   addends_reg_4_5_inst : DFF_X1 port map( D => pipe1_0_5_port, CK => CLOCK, Q 
                           => addends_4_5_port, QN => n_1554);
   pipe1_reg_0_4_inst : DFF_X1 port map( D => mux_out_4_4_port, CK => CLOCK, Q 
                           => pipe1_0_4_port, QN => n_1555);
   addends_reg_4_4_inst : DFF_X1 port map( D => pipe1_0_4_port, CK => CLOCK, Q 
                           => addends_4_4_port, QN => n_1556);
   pipe1_reg_0_3_inst : DFF_X1 port map( D => mux_out_4_3_port, CK => CLOCK, Q 
                           => pipe1_0_3_port, QN => n_1557);
   addends_reg_4_3_inst : DFF_X1 port map( D => pipe1_0_3_port, CK => CLOCK, Q 
                           => addends_4_3_port, QN => n_1558);
   pipe1_reg_0_2_inst : DFF_X1 port map( D => mux_out_4_2_port, CK => CLOCK, Q 
                           => pipe1_0_2_port, QN => n_1559);
   addends_reg_4_2_inst : DFF_X1 port map( D => pipe1_0_2_port, CK => CLOCK, Q 
                           => addends_4_2_port, QN => n_1560);
   pipe1_reg_0_1_inst : DFF_X1 port map( D => mux_out_4_1_port, CK => CLOCK, Q 
                           => pipe1_0_1_port, QN => n_1561);
   addends_reg_4_1_inst : DFF_X1 port map( D => pipe1_0_1_port, CK => CLOCK, Q 
                           => addends_4_1_port, QN => n_1562);
   pipe1_reg_0_0_inst : DFF_X1 port map( D => mux_out_4_0_port, CK => CLOCK, Q 
                           => pipe1_0_0_port, QN => n_1563);
   pipe2_reg_1_31_inst : DFF_X1 port map( D => pipe1_3_31_port, CK => CLOCK, Q 
                           => pipe2_1_31_port, QN => n_1564);
   addends_reg_7_31_inst : DFF_X1 port map( D => pipe2_1_31_port, CK => CLOCK, 
                           Q => addends_7_31_port, QN => n_1565);
   pipe2_reg_1_30_inst : DFF_X1 port map( D => pipe1_3_30_port, CK => CLOCK, Q 
                           => pipe2_1_30_port, QN => n_1566);
   addends_reg_7_30_inst : DFF_X1 port map( D => pipe2_1_30_port, CK => CLOCK, 
                           Q => addends_7_30_port, QN => n_1567);
   pipe2_reg_1_29_inst : DFF_X1 port map( D => pipe1_3_29_port, CK => CLOCK, Q 
                           => pipe2_1_29_port, QN => n_1568);
   addends_reg_7_29_inst : DFF_X1 port map( D => pipe2_1_29_port, CK => CLOCK, 
                           Q => addends_7_29_port, QN => n_1569);
   pipe2_reg_1_28_inst : DFF_X1 port map( D => pipe1_3_28_port, CK => CLOCK, Q 
                           => pipe2_1_28_port, QN => n_1570);
   addends_reg_7_28_inst : DFF_X1 port map( D => pipe2_1_28_port, CK => CLOCK, 
                           Q => addends_7_28_port, QN => n_1571);
   pipe2_reg_1_27_inst : DFF_X1 port map( D => pipe1_3_27_port, CK => CLOCK, Q 
                           => pipe2_1_27_port, QN => n_1572);
   addends_reg_7_27_inst : DFF_X1 port map( D => pipe2_1_27_port, CK => CLOCK, 
                           Q => addends_7_27_port, QN => n_1573);
   pipe2_reg_1_26_inst : DFF_X1 port map( D => pipe1_3_26_port, CK => CLOCK, Q 
                           => pipe2_1_26_port, QN => n_1574);
   addends_reg_7_26_inst : DFF_X1 port map( D => pipe2_1_26_port, CK => CLOCK, 
                           Q => addends_7_26_port, QN => n_1575);
   pipe2_reg_1_25_inst : DFF_X1 port map( D => pipe1_3_25_port, CK => CLOCK, Q 
                           => pipe2_1_25_port, QN => n_1576);
   addends_reg_7_25_inst : DFF_X1 port map( D => pipe2_1_25_port, CK => CLOCK, 
                           Q => addends_7_25_port, QN => n_1577);
   pipe2_reg_1_24_inst : DFF_X1 port map( D => pipe1_3_24_port, CK => CLOCK, Q 
                           => pipe2_1_24_port, QN => n_1578);
   addends_reg_7_24_inst : DFF_X1 port map( D => pipe2_1_24_port, CK => CLOCK, 
                           Q => addends_7_24_port, QN => n_1579);
   pipe2_reg_1_23_inst : DFF_X1 port map( D => pipe1_3_23_port, CK => CLOCK, Q 
                           => pipe2_1_23_port, QN => n_1580);
   addends_reg_7_23_inst : DFF_X1 port map( D => pipe2_1_23_port, CK => CLOCK, 
                           Q => addends_7_23_port, QN => n_1581);
   pipe2_reg_1_22_inst : DFF_X1 port map( D => pipe1_3_22_port, CK => CLOCK, Q 
                           => pipe2_1_22_port, QN => n_1582);
   addends_reg_7_22_inst : DFF_X1 port map( D => pipe2_1_22_port, CK => CLOCK, 
                           Q => addends_7_22_port, QN => n_1583);
   pipe2_reg_1_21_inst : DFF_X1 port map( D => pipe1_3_21_port, CK => CLOCK, Q 
                           => pipe2_1_21_port, QN => n_1584);
   addends_reg_7_21_inst : DFF_X1 port map( D => pipe2_1_21_port, CK => CLOCK, 
                           Q => addends_7_21_port, QN => n_1585);
   pipe2_reg_1_20_inst : DFF_X1 port map( D => pipe1_3_20_port, CK => CLOCK, Q 
                           => pipe2_1_20_port, QN => n_1586);
   addends_reg_7_20_inst : DFF_X1 port map( D => pipe2_1_20_port, CK => CLOCK, 
                           Q => addends_7_20_port, QN => n_1587);
   pipe2_reg_1_19_inst : DFF_X1 port map( D => pipe1_3_19_port, CK => CLOCK, Q 
                           => pipe2_1_19_port, QN => n_1588);
   addends_reg_7_19_inst : DFF_X1 port map( D => pipe2_1_19_port, CK => CLOCK, 
                           Q => addends_7_19_port, QN => n_1589);
   pipe2_reg_1_18_inst : DFF_X1 port map( D => pipe1_3_18_port, CK => CLOCK, Q 
                           => pipe2_1_18_port, QN => n_1590);
   addends_reg_7_18_inst : DFF_X1 port map( D => pipe2_1_18_port, CK => CLOCK, 
                           Q => addends_7_18_port, QN => n_1591);
   pipe2_reg_1_17_inst : DFF_X1 port map( D => pipe1_3_17_port, CK => CLOCK, Q 
                           => pipe2_1_17_port, QN => n_1592);
   addends_reg_7_17_inst : DFF_X1 port map( D => pipe2_1_17_port, CK => CLOCK, 
                           Q => addends_7_17_port, QN => n_1593);
   pipe2_reg_1_16_inst : DFF_X1 port map( D => pipe1_3_16_port, CK => CLOCK, Q 
                           => pipe2_1_16_port, QN => n_1594);
   addends_reg_7_16_inst : DFF_X1 port map( D => pipe2_1_16_port, CK => CLOCK, 
                           Q => addends_7_16_port, QN => n_1595);
   pipe2_reg_1_15_inst : DFF_X1 port map( D => pipe1_3_15_port, CK => CLOCK, Q 
                           => pipe2_1_15_port, QN => n_1596);
   addends_reg_7_15_inst : DFF_X1 port map( D => pipe2_1_15_port, CK => CLOCK, 
                           Q => addends_7_15_port, QN => n_1597);
   pipe2_reg_1_14_inst : DFF_X1 port map( D => pipe1_3_14_port, CK => CLOCK, Q 
                           => pipe2_1_14_port, QN => n_1598);
   addends_reg_7_14_inst : DFF_X1 port map( D => pipe2_1_14_port, CK => CLOCK, 
                           Q => addends_7_14_port, QN => n_1599);
   pipe2_reg_1_13_inst : DFF_X1 port map( D => pipe1_3_13_port, CK => CLOCK, Q 
                           => pipe2_1_13_port, QN => n_1600);
   addends_reg_7_13_inst : DFF_X1 port map( D => pipe2_1_13_port, CK => CLOCK, 
                           Q => addends_7_13_port, QN => n_1601);
   pipe2_reg_1_12_inst : DFF_X1 port map( D => pipe1_3_12_port, CK => CLOCK, Q 
                           => pipe2_1_12_port, QN => n_1602);
   addends_reg_7_12_inst : DFF_X1 port map( D => pipe2_1_12_port, CK => CLOCK, 
                           Q => addends_7_12_port, QN => n_1603);
   pipe2_reg_1_11_inst : DFF_X1 port map( D => pipe1_3_11_port, CK => CLOCK, Q 
                           => pipe2_1_11_port, QN => n_1604);
   addends_reg_7_11_inst : DFF_X1 port map( D => pipe2_1_11_port, CK => CLOCK, 
                           Q => addends_7_11_port, QN => n_1605);
   pipe2_reg_1_10_inst : DFF_X1 port map( D => pipe1_3_10_port, CK => CLOCK, Q 
                           => pipe2_1_10_port, QN => n_1606);
   addends_reg_7_10_inst : DFF_X1 port map( D => pipe2_1_10_port, CK => CLOCK, 
                           Q => addends_7_10_port, QN => n_1607);
   pipe2_reg_1_9_inst : DFF_X1 port map( D => pipe1_3_9_port, CK => CLOCK, Q =>
                           pipe2_1_9_port, QN => n_1608);
   addends_reg_7_9_inst : DFF_X1 port map( D => pipe2_1_9_port, CK => CLOCK, Q 
                           => addends_7_9_port, QN => n_1609);
   pipe2_reg_1_8_inst : DFF_X1 port map( D => pipe1_3_8_port, CK => CLOCK, Q =>
                           pipe2_1_8_port, QN => n_1610);
   addends_reg_7_8_inst : DFF_X1 port map( D => pipe2_1_8_port, CK => CLOCK, Q 
                           => addends_7_8_port, QN => n_1611);
   pipe2_reg_1_7_inst : DFF_X1 port map( D => pipe1_3_7_port, CK => CLOCK, Q =>
                           pipe2_1_7_port, QN => n_1612);
   addends_reg_7_7_inst : DFF_X1 port map( D => pipe2_1_7_port, CK => CLOCK, Q 
                           => addends_7_7_port, QN => n_1613);
   pipe2_reg_1_6_inst : DFF_X1 port map( D => pipe1_3_6_port, CK => CLOCK, Q =>
                           pipe2_1_6_port, QN => n_1614);
   addends_reg_7_6_inst : DFF_X1 port map( D => pipe2_1_6_port, CK => CLOCK, Q 
                           => addends_7_6_port, QN => n_1615);
   pipe2_reg_1_5_inst : DFF_X1 port map( D => pipe1_3_5_port, CK => CLOCK, Q =>
                           pipe2_1_5_port, QN => n_1616);
   addends_reg_7_5_inst : DFF_X1 port map( D => pipe2_1_5_port, CK => CLOCK, Q 
                           => addends_7_5_port, QN => n_1617);
   pipe2_reg_1_4_inst : DFF_X1 port map( D => pipe1_3_4_port, CK => CLOCK, Q =>
                           pipe2_1_4_port, QN => n_1618);
   addends_reg_7_4_inst : DFF_X1 port map( D => pipe2_1_4_port, CK => CLOCK, Q 
                           => addends_7_4_port, QN => n_1619);
   pipe2_reg_1_3_inst : DFF_X1 port map( D => pipe1_3_3_port, CK => CLOCK, Q =>
                           pipe2_1_3_port, QN => n_1620);
   addends_reg_7_3_inst : DFF_X1 port map( D => pipe2_1_3_port, CK => CLOCK, Q 
                           => addends_7_3_port, QN => n_1621);
   pipe2_reg_1_2_inst : DFF_X1 port map( D => pipe1_3_2_port, CK => CLOCK, Q =>
                           pipe2_1_2_port, QN => n_1622);
   addends_reg_7_2_inst : DFF_X1 port map( D => pipe2_1_2_port, CK => CLOCK, Q 
                           => addends_7_2_port, QN => n_1623);
   pipe2_reg_1_1_inst : DFF_X1 port map( D => pipe1_3_1_port, CK => CLOCK, Q =>
                           pipe2_1_1_port, QN => n_1624);
   addends_reg_7_1_inst : DFF_X1 port map( D => pipe2_1_1_port, CK => CLOCK, Q 
                           => addends_7_1_port, QN => n_1625);
   pipe2_reg_1_0_inst : DFF_X1 port map( D => pipe1_3_0_port, CK => CLOCK, Q =>
                           pipe2_1_0_port, QN => n_1626);
   addends_reg_7_0_inst : DFF_X1 port map( D => pipe2_1_0_port, CK => CLOCK, Q 
                           => addends_7_0_port, QN => n_1627);
   pipe2_reg_0_31_inst : DFF_X1 port map( D => pipe1_2_31_port, CK => CLOCK, Q 
                           => pipe2_0_31_port, QN => n_1628);
   addends_reg_6_31_inst : DFF_X1 port map( D => pipe2_0_31_port, CK => CLOCK, 
                           Q => addends_6_31_port, QN => n_1629);
   pipe2_reg_0_30_inst : DFF_X1 port map( D => pipe1_2_30_port, CK => CLOCK, Q 
                           => pipe2_0_30_port, QN => n_1630);
   addends_reg_6_30_inst : DFF_X1 port map( D => pipe2_0_30_port, CK => CLOCK, 
                           Q => addends_6_30_port, QN => n_1631);
   pipe2_reg_0_29_inst : DFF_X1 port map( D => pipe1_2_29_port, CK => CLOCK, Q 
                           => pipe2_0_29_port, QN => n_1632);
   addends_reg_6_29_inst : DFF_X1 port map( D => pipe2_0_29_port, CK => CLOCK, 
                           Q => addends_6_29_port, QN => n_1633);
   pipe2_reg_0_28_inst : DFF_X1 port map( D => pipe1_2_28_port, CK => CLOCK, Q 
                           => pipe2_0_28_port, QN => n_1634);
   addends_reg_6_28_inst : DFF_X1 port map( D => pipe2_0_28_port, CK => CLOCK, 
                           Q => addends_6_28_port, QN => n_1635);
   pipe2_reg_0_27_inst : DFF_X1 port map( D => pipe1_2_27_port, CK => CLOCK, Q 
                           => pipe2_0_27_port, QN => n_1636);
   addends_reg_6_27_inst : DFF_X1 port map( D => pipe2_0_27_port, CK => CLOCK, 
                           Q => addends_6_27_port, QN => n_1637);
   pipe2_reg_0_26_inst : DFF_X1 port map( D => pipe1_2_26_port, CK => CLOCK, Q 
                           => pipe2_0_26_port, QN => n_1638);
   addends_reg_6_26_inst : DFF_X1 port map( D => pipe2_0_26_port, CK => CLOCK, 
                           Q => addends_6_26_port, QN => n_1639);
   pipe2_reg_0_25_inst : DFF_X1 port map( D => pipe1_2_25_port, CK => CLOCK, Q 
                           => pipe2_0_25_port, QN => n_1640);
   addends_reg_6_25_inst : DFF_X1 port map( D => pipe2_0_25_port, CK => CLOCK, 
                           Q => addends_6_25_port, QN => n_1641);
   pipe2_reg_0_24_inst : DFF_X1 port map( D => pipe1_2_24_port, CK => CLOCK, Q 
                           => pipe2_0_24_port, QN => n_1642);
   addends_reg_6_24_inst : DFF_X1 port map( D => pipe2_0_24_port, CK => CLOCK, 
                           Q => addends_6_24_port, QN => n_1643);
   pipe2_reg_0_23_inst : DFF_X1 port map( D => pipe1_2_23_port, CK => CLOCK, Q 
                           => pipe2_0_23_port, QN => n_1644);
   addends_reg_6_23_inst : DFF_X1 port map( D => pipe2_0_23_port, CK => CLOCK, 
                           Q => addends_6_23_port, QN => n_1645);
   pipe2_reg_0_22_inst : DFF_X1 port map( D => pipe1_2_22_port, CK => CLOCK, Q 
                           => pipe2_0_22_port, QN => n_1646);
   addends_reg_6_22_inst : DFF_X1 port map( D => pipe2_0_22_port, CK => CLOCK, 
                           Q => addends_6_22_port, QN => n_1647);
   pipe2_reg_0_21_inst : DFF_X1 port map( D => pipe1_2_21_port, CK => CLOCK, Q 
                           => pipe2_0_21_port, QN => n_1648);
   addends_reg_6_21_inst : DFF_X1 port map( D => pipe2_0_21_port, CK => CLOCK, 
                           Q => addends_6_21_port, QN => n_1649);
   pipe2_reg_0_20_inst : DFF_X1 port map( D => pipe1_2_20_port, CK => CLOCK, Q 
                           => pipe2_0_20_port, QN => n_1650);
   addends_reg_6_20_inst : DFF_X1 port map( D => pipe2_0_20_port, CK => CLOCK, 
                           Q => addends_6_20_port, QN => n_1651);
   pipe2_reg_0_19_inst : DFF_X1 port map( D => pipe1_2_19_port, CK => CLOCK, Q 
                           => pipe2_0_19_port, QN => n_1652);
   addends_reg_6_19_inst : DFF_X1 port map( D => pipe2_0_19_port, CK => CLOCK, 
                           Q => addends_6_19_port, QN => n_1653);
   pipe2_reg_0_18_inst : DFF_X1 port map( D => pipe1_2_18_port, CK => CLOCK, Q 
                           => pipe2_0_18_port, QN => n_1654);
   addends_reg_6_18_inst : DFF_X1 port map( D => pipe2_0_18_port, CK => CLOCK, 
                           Q => addends_6_18_port, QN => n_1655);
   pipe2_reg_0_17_inst : DFF_X1 port map( D => pipe1_2_17_port, CK => CLOCK, Q 
                           => pipe2_0_17_port, QN => n_1656);
   addends_reg_6_17_inst : DFF_X1 port map( D => pipe2_0_17_port, CK => CLOCK, 
                           Q => addends_6_17_port, QN => n_1657);
   pipe2_reg_0_16_inst : DFF_X1 port map( D => pipe1_2_16_port, CK => CLOCK, Q 
                           => pipe2_0_16_port, QN => n_1658);
   addends_reg_6_16_inst : DFF_X1 port map( D => pipe2_0_16_port, CK => CLOCK, 
                           Q => addends_6_16_port, QN => n_1659);
   pipe2_reg_0_15_inst : DFF_X1 port map( D => pipe1_2_15_port, CK => CLOCK, Q 
                           => pipe2_0_15_port, QN => n_1660);
   pipe2_reg_0_14_inst : DFF_X1 port map( D => pipe1_2_14_port, CK => CLOCK, Q 
                           => pipe2_0_14_port, QN => n_1661);
   addends_reg_6_14_inst : DFF_X1 port map( D => pipe2_0_14_port, CK => CLOCK, 
                           Q => addends_6_14_port, QN => n_1662);
   pipe2_reg_0_13_inst : DFF_X1 port map( D => pipe1_2_13_port, CK => CLOCK, Q 
                           => pipe2_0_13_port, QN => n_1663);
   addends_reg_6_13_inst : DFF_X1 port map( D => pipe2_0_13_port, CK => CLOCK, 
                           Q => addends_6_13_port, QN => n_1664);
   pipe2_reg_0_12_inst : DFF_X1 port map( D => pipe1_2_12_port, CK => CLOCK, Q 
                           => pipe2_0_12_port, QN => n_1665);
   addends_reg_6_12_inst : DFF_X1 port map( D => pipe2_0_12_port, CK => CLOCK, 
                           Q => addends_6_12_port, QN => n_1666);
   pipe2_reg_0_11_inst : DFF_X1 port map( D => pipe1_2_11_port, CK => CLOCK, Q 
                           => pipe2_0_11_port, QN => n_1667);
   addends_reg_6_11_inst : DFF_X1 port map( D => pipe2_0_11_port, CK => CLOCK, 
                           Q => addends_6_11_port, QN => n_1668);
   pipe2_reg_0_10_inst : DFF_X1 port map( D => pipe1_2_10_port, CK => CLOCK, Q 
                           => pipe2_0_10_port, QN => n_1669);
   addends_reg_6_10_inst : DFF_X1 port map( D => pipe2_0_10_port, CK => CLOCK, 
                           Q => addends_6_10_port, QN => n_1670);
   pipe2_reg_0_9_inst : DFF_X1 port map( D => pipe1_2_9_port, CK => CLOCK, Q =>
                           pipe2_0_9_port, QN => n_1671);
   addends_reg_6_9_inst : DFF_X1 port map( D => pipe2_0_9_port, CK => CLOCK, Q 
                           => addends_6_9_port, QN => n_1672);
   pipe2_reg_0_8_inst : DFF_X1 port map( D => pipe1_2_8_port, CK => CLOCK, Q =>
                           pipe2_0_8_port, QN => n_1673);
   addends_reg_6_8_inst : DFF_X1 port map( D => pipe2_0_8_port, CK => CLOCK, Q 
                           => addends_6_8_port, QN => n_1674);
   pipe2_reg_0_7_inst : DFF_X1 port map( D => pipe1_2_7_port, CK => CLOCK, Q =>
                           pipe2_0_7_port, QN => n_1675);
   addends_reg_6_7_inst : DFF_X1 port map( D => pipe2_0_7_port, CK => CLOCK, Q 
                           => addends_6_7_port, QN => n_1676);
   pipe2_reg_0_6_inst : DFF_X1 port map( D => pipe1_2_6_port, CK => CLOCK, Q =>
                           pipe2_0_6_port, QN => n_1677);
   pipe2_reg_0_5_inst : DFF_X1 port map( D => pipe1_2_5_port, CK => CLOCK, Q =>
                           pipe2_0_5_port, QN => n_1678);
   addends_reg_6_5_inst : DFF_X1 port map( D => pipe2_0_5_port, CK => CLOCK, Q 
                           => addends_6_5_port, QN => n_1679);
   pipe2_reg_0_4_inst : DFF_X1 port map( D => pipe1_2_4_port, CK => CLOCK, Q =>
                           pipe2_0_4_port, QN => n_1680);
   pipe2_reg_0_3_inst : DFF_X1 port map( D => pipe1_2_3_port, CK => CLOCK, Q =>
                           pipe2_0_3_port, QN => n_1681);
   addends_reg_6_3_inst : DFF_X1 port map( D => pipe2_0_3_port, CK => CLOCK, Q 
                           => addends_6_3_port, QN => n_1682);
   pipe2_reg_0_2_inst : DFF_X1 port map( D => pipe1_2_2_port, CK => CLOCK, Q =>
                           pipe2_0_2_port, QN => n_1683);
   addends_reg_6_2_inst : DFF_X1 port map( D => pipe2_0_2_port, CK => CLOCK, Q 
                           => addends_6_2_port, QN => n_1684);
   pipe2_reg_0_1_inst : DFF_X1 port map( D => pipe1_2_1_port, CK => CLOCK, Q =>
                           pipe2_0_1_port, QN => n_1685);
   pipe2_reg_0_0_inst : DFF_X1 port map( D => pipe1_2_0_port, CK => CLOCK, Q =>
                           pipe2_0_0_port, QN => n_1686);
   enc_1 : ENCODER_0 port map( INPUT(2) => B(1), INPUT(1) => B(0), INPUT(0) => 
                           X_Logic0_port, OUTPUT(2) => selector_2_port, 
                           OUTPUT(1) => selector_1_port, OUTPUT(0) => 
                           selector_0_port);
   enc_2 : ENCODER_7 port map( INPUT(2) => B(3), INPUT(1) => B(2), INPUT(0) => 
                           B(1), OUTPUT(2) => selector_5_port, OUTPUT(1) => 
                           selector_4_port, OUTPUT(0) => selector_3_port);
   enc_3 : ENCODER_6 port map( INPUT(2) => B(5), INPUT(1) => B(4), INPUT(0) => 
                           B(3), OUTPUT(2) => selector_8_port, OUTPUT(1) => 
                           selector_7_port, OUTPUT(0) => selector_6_port);
   enc_4 : ENCODER_5 port map( INPUT(2) => B(7), INPUT(1) => B(6), INPUT(0) => 
                           B(5), OUTPUT(2) => selector_11_port, OUTPUT(1) => 
                           selector_10_port, OUTPUT(0) => selector_9_port);
   enc_5 : ENCODER_4 port map( INPUT(2) => B(9), INPUT(1) => B(8), INPUT(0) => 
                           B(7), OUTPUT(2) => selector_14_port, OUTPUT(1) => 
                           selector_13_port, OUTPUT(0) => selector_12_port);
   enc_6 : ENCODER_3 port map( INPUT(2) => B(11), INPUT(1) => B(10), INPUT(0) 
                           => B(9), OUTPUT(2) => selector_17_port, OUTPUT(1) =>
                           selector_16_port, OUTPUT(0) => selector_15_port);
   enc_7 : ENCODER_2 port map( INPUT(2) => B(13), INPUT(1) => B(12), INPUT(0) 
                           => B(11), OUTPUT(2) => selector_20_port, OUTPUT(1) 
                           => selector_19_port, OUTPUT(0) => selector_18_port);
   enc_8 : ENCODER_1 port map( INPUT(2) => B(15), INPUT(1) => B(14), INPUT(0) 
                           => B(13), OUTPUT(2) => selector_23_port, OUTPUT(1) 
                           => selector_22_port, OUTPUT(0) => selector_21_port);
   MUX_I_0 : MUX5to1_NBIT32_8 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => A(15), B(14) => A(14), B(13)
                           => A(13), B(12) => A(12), B(11) => A(11), B(10) => 
                           A(10), B(9) => A(9), B(8) => A(8), B(7) => A(7), 
                           B(6) => A(6), B(5) => A(5), B(4) => A(4), B(3) => 
                           A(3), B(2) => A(2), B(1) => A(1), B(0) => n21, C(31)
                           => n6, C(30) => n6, C(29) => n6, C(28) => n6, C(27) 
                           => n6, C(26) => n6, C(25) => n6, C(24) => n6, C(23) 
                           => n6, C(22) => n6, C(21) => n6, C(20) => n6, C(19) 
                           => n6, C(18) => n6, C(17) => n6, C(16) => n6, C(15) 
                           => A_neg_0_15_port, C(14) => A_neg_0_14_port, C(13) 
                           => A_neg_0_13_port, C(12) => A_neg_0_12_port, C(11) 
                           => A_neg_0_11_port, C(10) => A_neg_0_10_port, C(9) 
                           => A_neg_0_9_port, C(8) => A_neg_0_8_port, C(7) => 
                           A_neg_0_7_port, C(6) => A_neg_0_6_port, C(5) => 
                           A_neg_0_5_port, C(4) => A_neg_0_4_port, C(3) => 
                           A_neg_0_3_port, C(2) => A_neg_0_2_port, C(1) => 
                           A_neg_0_1_port, C(0) => n21, D(31) => X_Logic0_port,
                           D(30) => X_Logic0_port, D(29) => X_Logic0_port, 
                           D(28) => X_Logic0_port, D(27) => X_Logic0_port, 
                           D(26) => X_Logic0_port, D(25) => X_Logic0_port, 
                           D(24) => X_Logic0_port, D(23) => X_Logic0_port, 
                           D(22) => X_Logic0_port, D(21) => X_Logic0_port, 
                           D(20) => X_Logic0_port, D(19) => X_Logic0_port, 
                           D(18) => X_Logic0_port, D(17) => X_Logic0_port, 
                           D(16) => A(15), D(15) => A(14), D(14) => A(13), 
                           D(13) => A(12), D(12) => A(11), D(11) => A(10), 
                           D(10) => A(9), D(9) => A(8), D(8) => A(7), D(7) => 
                           A(6), D(6) => A(5), D(5) => A(4), D(4) => A(3), D(3)
                           => A(2), D(2) => A(1), D(1) => A(0), D(0) => 
                           X_Logic0_port, E(31) => n8, E(30) => n8, E(29) => n8
                           , E(28) => n8, E(27) => n8, E(26) => n8, E(25) => n8
                           , E(24) => n8, E(23) => n8, E(22) => n8, E(21) => n8
                           , E(20) => n8, E(19) => n8, E(18) => n8, E(17) => n8
                           , E(16) => A_neg_1_16_port, E(15) => A_neg_1_15_port
                           , E(14) => A_neg_1_14_port, E(13) => A_neg_1_13_port
                           , E(12) => A_neg_1_12_port, E(11) => A_neg_1_11_port
                           , E(10) => A_neg_1_10_port, E(9) => A_neg_1_9_port, 
                           E(8) => A_neg_1_8_port, E(7) => A_neg_1_7_port, E(6)
                           => A_neg_1_6_port, E(5) => A_neg_1_5_port, E(4) => 
                           A_neg_1_4_port, E(3) => A_neg_1_3_port, E(2) => 
                           A_neg_1_2_port, E(1) => A(0), E(0) => n70, SEL(2) =>
                           selector_2_port, SEL(1) => selector_1_port, SEL(0) 
                           => selector_0_port, Y(31) => addends_0_31_port, 
                           Y(30) => addends_0_30_port, Y(29) => 
                           addends_0_29_port, Y(28) => addends_0_28_port, Y(27)
                           => addends_0_27_port, Y(26) => addends_0_26_port, 
                           Y(25) => addends_0_25_port, Y(24) => 
                           addends_0_24_port, Y(23) => addends_0_23_port, Y(22)
                           => addends_0_22_port, Y(21) => addends_0_21_port, 
                           Y(20) => addends_0_20_port, Y(19) => 
                           addends_0_19_port, Y(18) => addends_0_18_port, Y(17)
                           => addends_0_17_port, Y(16) => addends_0_16_port, 
                           Y(15) => addends_0_15_port, Y(14) => 
                           addends_0_14_port, Y(13) => addends_0_13_port, Y(12)
                           => addends_0_12_port, Y(11) => addends_0_11_port, 
                           Y(10) => addends_0_10_port, Y(9) => addends_0_9_port
                           , Y(8) => addends_0_8_port, Y(7) => addends_0_7_port
                           , Y(6) => addends_0_6_port, Y(5) => addends_0_5_port
                           , Y(4) => addends_0_4_port, Y(3) => addends_0_3_port
                           , Y(2) => addends_0_2_port, Y(1) => addends_0_1_port
                           , Y(0) => addends_0_0_port);
   MUX_I_1 : MUX5to1_NBIT32_7 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => A(15), B(16) => A(14), B(15)
                           => A(13), B(14) => A(12), B(13) => A(11), B(12) => 
                           A(10), B(11) => A(9), B(10) => A(8), B(9) => A(7), 
                           B(8) => A(6), B(7) => A(5), B(6) => A(4), B(5) => 
                           A(3), B(4) => A(2), B(3) => A(1), B(2) => A(0), B(1)
                           => X_Logic0_port, B(0) => X_Logic0_port, C(31) => n9
                           , C(30) => n9, C(29) => n9, C(28) => n9, C(27) => n9
                           , C(26) => n9, C(25) => n9, C(24) => n9, C(23) => n9
                           , C(22) => n9, C(21) => n9, C(20) => n9, C(19) => n9
                           , C(18) => n9, C(17) => A_neg_2_17_port, C(16) => 
                           A_neg_2_16_port, C(15) => A_neg_2_15_port, C(14) => 
                           A_neg_2_14_port, C(13) => A_neg_2_13_port, C(12) => 
                           A_neg_2_12_port, C(11) => A_neg_2_11_port, C(10) => 
                           A_neg_2_10_port, C(9) => A_neg_2_9_port, C(8) => 
                           A_neg_2_8_port, C(7) => A_neg_2_7_port, C(6) => 
                           A_neg_2_6_port, C(5) => A_neg_2_5_port, C(4) => 
                           A_neg_2_4_port, C(3) => A_neg_2_3_port, C(2) => n21,
                           C(1) => n70, C(0) => n70, D(31) => X_Logic0_port, 
                           D(30) => X_Logic0_port, D(29) => X_Logic0_port, 
                           D(28) => X_Logic0_port, D(27) => X_Logic0_port, 
                           D(26) => X_Logic0_port, D(25) => X_Logic0_port, 
                           D(24) => X_Logic0_port, D(23) => X_Logic0_port, 
                           D(22) => X_Logic0_port, D(21) => X_Logic0_port, 
                           D(20) => X_Logic0_port, D(19) => X_Logic0_port, 
                           D(18) => A(15), D(17) => A(14), D(16) => A(13), 
                           D(15) => A(12), D(14) => A(11), D(13) => A(10), 
                           D(12) => A(9), D(11) => A(8), D(10) => A(7), D(9) =>
                           A(6), D(8) => A(5), D(7) => A(4), D(6) => A(3), D(5)
                           => A(2), D(4) => A(1), D(3) => A(0), D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n11, E(30) => n11, E(29) => 
                           n11, E(28) => n11, E(27) => n11, E(26) => n11, E(25)
                           => n11, E(24) => n11, E(23) => n11, E(22) => n11, 
                           E(21) => n11, E(20) => n11, E(19) => n11, E(18) => 
                           A_neg_3_18_port, E(17) => A_neg_3_17_port, E(16) => 
                           A_neg_3_16_port, E(15) => A_neg_3_15_port, E(14) => 
                           A_neg_3_14_port, E(13) => A_neg_3_13_port, E(12) => 
                           A_neg_3_12_port, E(11) => A_neg_3_11_port, E(10) => 
                           A_neg_3_10_port, E(9) => A_neg_3_9_port, E(8) => 
                           A_neg_3_8_port, E(7) => A_neg_3_7_port, E(6) => 
                           A_neg_3_6_port, E(5) => A_neg_3_5_port, E(4) => 
                           A_neg_3_4_port, E(3) => A(0), E(2) => n70, E(1) => 
                           n70, E(0) => n70, SEL(2) => selector_5_port, SEL(1) 
                           => selector_4_port, SEL(0) => selector_3_port, Y(31)
                           => addends_1_31_port, Y(30) => addends_1_30_port, 
                           Y(29) => addends_1_29_port, Y(28) => 
                           addends_1_28_port, Y(27) => addends_1_27_port, Y(26)
                           => addends_1_26_port, Y(25) => addends_1_25_port, 
                           Y(24) => addends_1_24_port, Y(23) => 
                           addends_1_23_port, Y(22) => addends_1_22_port, Y(21)
                           => addends_1_21_port, Y(20) => addends_1_20_port, 
                           Y(19) => addends_1_19_port, Y(18) => 
                           addends_1_18_port, Y(17) => addends_1_17_port, Y(16)
                           => addends_1_16_port, Y(15) => addends_1_15_port, 
                           Y(14) => addends_1_14_port, Y(13) => 
                           addends_1_13_port, Y(12) => addends_1_12_port, Y(11)
                           => addends_1_11_port, Y(10) => addends_1_10_port, 
                           Y(9) => addends_1_9_port, Y(8) => addends_1_8_port, 
                           Y(7) => addends_1_7_port, Y(6) => addends_1_6_port, 
                           Y(5) => addends_1_5_port, Y(4) => addends_1_4_port, 
                           Y(3) => addends_1_3_port, Y(2) => addends_1_2_port, 
                           Y(1) => addends_1_1_port, Y(0) => addends_1_0_port);
   MUX_I_2 : MUX5to1_NBIT32_6 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => A(15), B(18) => A(14), B(17)
                           => A(13), B(16) => A(12), B(15) => A(11), B(14) => 
                           A(10), B(13) => A(9), B(12) => A(8), B(11) => A(7), 
                           B(10) => A(6), B(9) => A(5), B(8) => A(4), B(7) => 
                           A(3), B(6) => A(2), B(5) => A(1), B(4) => A(0), B(3)
                           => X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n12, 
                           C(30) => n12, C(29) => n12, C(28) => n12, C(27) => 
                           n12, C(26) => n12, C(25) => n12, C(24) => n12, C(23)
                           => n12, C(22) => n12, C(21) => n12, C(20) => n12, 
                           C(19) => A_neg_4_19_port, C(18) => A_neg_4_18_port, 
                           C(17) => A_neg_4_17_port, C(16) => A_neg_4_16_port, 
                           C(15) => A_neg_4_15_port, C(14) => A_neg_4_14_port, 
                           C(13) => A_neg_4_13_port, C(12) => A_neg_4_12_port, 
                           C(11) => A_neg_4_11_port, C(10) => A_neg_4_10_port, 
                           C(9) => A_neg_4_9_port, C(8) => A_neg_4_8_port, C(7)
                           => A_neg_4_7_port, C(6) => A_neg_4_6_port, C(5) => 
                           A_neg_4_5_port, C(4) => n21, C(3) => n70, C(2) => 
                           n70, C(1) => n70, C(0) => n70, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => A(15), D(19) => A(14), D(18)
                           => A(13), D(17) => A(12), D(16) => A(11), D(15) => 
                           A(10), D(14) => A(9), D(13) => A(8), D(12) => A(7), 
                           D(11) => A(6), D(10) => A(5), D(9) => A(4), D(8) => 
                           A(3), D(7) => A(2), D(6) => A(1), D(5) => A(0), D(4)
                           => X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n3, E(30) => n3, E(29) => n3
                           , E(28) => n3, E(27) => n3, E(26) => n3, E(25) => n3
                           , E(24) => n3, E(23) => n3, E(22) => n3, E(21) => n3
                           , E(20) => A_neg_5_20_port, E(19) => A_neg_5_19_port
                           , E(18) => A_neg_5_18_port, E(17) => A_neg_5_17_port
                           , E(16) => A_neg_5_16_port, E(15) => A_neg_5_15_port
                           , E(14) => A_neg_5_14_port, E(13) => A_neg_5_13_port
                           , E(12) => A_neg_5_12_port, E(11) => A_neg_5_11_port
                           , E(10) => A_neg_5_10_port, E(9) => A_neg_5_9_port, 
                           E(8) => A_neg_5_8_port, E(7) => A_neg_5_7_port, E(6)
                           => A_neg_5_6_port, E(5) => A(0), E(4) => n70, E(3) 
                           => n70, E(2) => n70, E(1) => n70, E(0) => n70, 
                           SEL(2) => selector_8_port, SEL(1) => selector_7_port
                           , SEL(0) => selector_6_port, Y(31) => 
                           mux_out_2_31_port, Y(30) => mux_out_2_30_port, Y(29)
                           => mux_out_2_29_port, Y(28) => mux_out_2_28_port, 
                           Y(27) => mux_out_2_27_port, Y(26) => 
                           mux_out_2_26_port, Y(25) => mux_out_2_25_port, Y(24)
                           => mux_out_2_24_port, Y(23) => mux_out_2_23_port, 
                           Y(22) => mux_out_2_22_port, Y(21) => 
                           mux_out_2_21_port, Y(20) => mux_out_2_20_port, Y(19)
                           => mux_out_2_19_port, Y(18) => mux_out_2_18_port, 
                           Y(17) => mux_out_2_17_port, Y(16) => 
                           mux_out_2_16_port, Y(15) => mux_out_2_15_port, Y(14)
                           => mux_out_2_14_port, Y(13) => mux_out_2_13_port, 
                           Y(12) => mux_out_2_12_port, Y(11) => 
                           mux_out_2_11_port, Y(10) => mux_out_2_10_port, Y(9) 
                           => mux_out_2_9_port, Y(8) => mux_out_2_8_port, Y(7) 
                           => mux_out_2_7_port, Y(6) => mux_out_2_6_port, Y(5) 
                           => mux_out_2_5_port, Y(4) => mux_out_2_4_port, Y(3) 
                           => mux_out_2_3_port, Y(2) => mux_out_2_2_port, Y(1) 
                           => mux_out_2_1_port, Y(0) => mux_out_2_0_port);
   MUX_I_3 : MUX5to1_NBIT32_5 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => A(15), B(20) => A(14), B(19)
                           => A(13), B(18) => A(12), B(17) => A(11), B(16) => 
                           A(10), B(15) => A(9), B(14) => A(8), B(13) => A(7), 
                           B(12) => A(6), B(11) => A(5), B(10) => A(4), B(9) =>
                           A(3), B(8) => A(2), B(7) => A(1), B(6) => n21, B(5) 
                           => X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n4, 
                           C(30) => n4, C(29) => n4, C(28) => n4, C(27) => n4, 
                           C(26) => n4, C(25) => n4, C(24) => n4, C(23) => n4, 
                           C(22) => n4, C(21) => A_neg_6_21_port, C(20) => 
                           A_neg_6_20_port, C(19) => A_neg_6_19_port, C(18) => 
                           A_neg_6_18_port, C(17) => A_neg_6_17_port, C(16) => 
                           A_neg_6_16_port, C(15) => A_neg_6_15_port, C(14) => 
                           A_neg_6_14_port, C(13) => A_neg_6_13_port, C(12) => 
                           A_neg_6_12_port, C(11) => A_neg_6_11_port, C(10) => 
                           A_neg_6_10_port, C(9) => A_neg_6_9_port, C(8) => 
                           A_neg_6_8_port, C(7) => A_neg_6_7_port, C(6) => n21,
                           C(5) => n70, C(4) => n70, C(3) => n70, C(2) => n70, 
                           C(1) => n70, C(0) => n70, D(31) => X_Logic0_port, 
                           D(30) => X_Logic0_port, D(29) => X_Logic0_port, 
                           D(28) => X_Logic0_port, D(27) => X_Logic0_port, 
                           D(26) => X_Logic0_port, D(25) => X_Logic0_port, 
                           D(24) => X_Logic0_port, D(23) => X_Logic0_port, 
                           D(22) => A(15), D(21) => A(14), D(20) => A(13), 
                           D(19) => A(12), D(18) => A(11), D(17) => A(10), 
                           D(16) => A(9), D(15) => A(8), D(14) => A(7), D(13) 
                           => A(6), D(12) => A(5), D(11) => A(4), D(10) => A(3)
                           , D(9) => A(2), D(8) => A(1), D(7) => A(0), D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n5, E(30) => n5, E(29) => n5
                           , E(28) => n5, E(27) => n5, E(26) => n5, E(25) => n5
                           , E(24) => n5, E(23) => n5, E(22) => A_neg_7_22_port
                           , E(21) => A_neg_7_21_port, E(20) => A_neg_7_20_port
                           , E(19) => A_neg_7_19_port, E(18) => A_neg_7_18_port
                           , E(17) => A_neg_7_17_port, E(16) => A_neg_7_16_port
                           , E(15) => A_neg_7_15_port, E(14) => A_neg_7_14_port
                           , E(13) => A_neg_7_13_port, E(12) => A_neg_7_12_port
                           , E(11) => A_neg_7_11_port, E(10) => A_neg_7_10_port
                           , E(9) => A_neg_7_9_port, E(8) => A_neg_7_8_port, 
                           E(7) => A(0), E(6) => n70, E(5) => n70, E(4) => n70,
                           E(3) => n70, E(2) => n70, E(1) => n70, E(0) => n70, 
                           SEL(2) => selector_11_port, SEL(1) => 
                           selector_10_port, SEL(0) => selector_9_port, Y(31) 
                           => mux_out_3_31_port, Y(30) => mux_out_3_30_port, 
                           Y(29) => mux_out_3_29_port, Y(28) => 
                           mux_out_3_28_port, Y(27) => mux_out_3_27_port, Y(26)
                           => mux_out_3_26_port, Y(25) => mux_out_3_25_port, 
                           Y(24) => mux_out_3_24_port, Y(23) => 
                           mux_out_3_23_port, Y(22) => mux_out_3_22_port, Y(21)
                           => mux_out_3_21_port, Y(20) => mux_out_3_20_port, 
                           Y(19) => mux_out_3_19_port, Y(18) => 
                           mux_out_3_18_port, Y(17) => mux_out_3_17_port, Y(16)
                           => mux_out_3_16_port, Y(15) => mux_out_3_15_port, 
                           Y(14) => mux_out_3_14_port, Y(13) => 
                           mux_out_3_13_port, Y(12) => mux_out_3_12_port, Y(11)
                           => mux_out_3_11_port, Y(10) => mux_out_3_10_port, 
                           Y(9) => mux_out_3_9_port, Y(8) => mux_out_3_8_port, 
                           Y(7) => mux_out_3_7_port, Y(6) => mux_out_3_6_port, 
                           Y(5) => mux_out_3_5_port, Y(4) => mux_out_3_4_port, 
                           Y(3) => mux_out_3_3_port, Y(2) => mux_out_3_2_port, 
                           Y(1) => mux_out_3_1_port, Y(0) => mux_out_3_0_port);
   MUX_I_4 : MUX5to1_NBIT32_4 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => A(15), B(22) => A(14), B(21)
                           => A(13), B(20) => A(12), B(19) => A(11), B(18) => 
                           A(10), B(17) => A(9), B(16) => A(8), B(15) => A(7), 
                           B(14) => A(6), B(13) => A(5), B(12) => A(4), B(11) 
                           => A(3), B(10) => A(2), B(9) => A(1), B(8) => n21, 
                           B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) 
                           => X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n7, 
                           C(30) => n7, C(29) => n7, C(28) => n7, C(27) => n7, 
                           C(26) => n7, C(25) => n7, C(24) => n7, C(23) => 
                           A_neg_8_23_port, C(22) => A_neg_8_22_port, C(21) => 
                           A_neg_8_21_port, C(20) => A_neg_8_20_port, C(19) => 
                           A_neg_8_19_port, C(18) => A_neg_8_18_port, C(17) => 
                           A_neg_8_17_port, C(16) => A_neg_8_16_port, C(15) => 
                           A_neg_8_15_port, C(14) => A_neg_8_14_port, C(13) => 
                           A_neg_8_13_port, C(12) => A_neg_8_12_port, C(11) => 
                           A_neg_8_11_port, C(10) => A_neg_8_10_port, C(9) => 
                           A_neg_8_9_port, C(8) => n21, C(7) => n70, C(6) => 
                           n70, C(5) => n70, C(4) => n70, C(3) => n70, C(2) => 
                           n70, C(1) => n70, C(0) => n70, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => A(15), D(23) => A(14), D(22)
                           => A(13), D(21) => A(12), D(20) => A(11), D(19) => 
                           A(10), D(18) => A(9), D(17) => A(8), D(16) => A(7), 
                           D(15) => A(6), D(14) => A(5), D(13) => A(4), D(12) 
                           => A(3), D(11) => A(2), D(10) => A(1), D(9) => A(0),
                           D(8) => X_Logic0_port, D(7) => X_Logic0_port, D(6) 
                           => X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n10, E(30) => n10, E(29) => 
                           n10, E(28) => n10, E(27) => n10, E(26) => n10, E(25)
                           => n10, E(24) => A_neg_9_24_port, E(23) => 
                           A_neg_9_23_port, E(22) => A_neg_9_22_port, E(21) => 
                           A_neg_9_21_port, E(20) => A_neg_9_20_port, E(19) => 
                           A_neg_9_19_port, E(18) => A_neg_9_18_port, E(17) => 
                           A_neg_9_17_port, E(16) => A_neg_9_16_port, E(15) => 
                           A_neg_9_15_port, E(14) => A_neg_9_14_port, E(13) => 
                           A_neg_9_13_port, E(12) => A_neg_9_12_port, E(11) => 
                           A_neg_9_11_port, E(10) => A_neg_9_10_port, E(9) => 
                           A(0), E(8) => n70, E(7) => n70, E(6) => n70, E(5) =>
                           n70, E(4) => n70, E(3) => n70, E(2) => n70, E(1) => 
                           n70, E(0) => n70, SEL(2) => selector_14_port, SEL(1)
                           => selector_13_port, SEL(0) => selector_12_port, 
                           Y(31) => mux_out_4_31_port, Y(30) => 
                           mux_out_4_30_port, Y(29) => mux_out_4_29_port, Y(28)
                           => mux_out_4_28_port, Y(27) => mux_out_4_27_port, 
                           Y(26) => mux_out_4_26_port, Y(25) => 
                           mux_out_4_25_port, Y(24) => mux_out_4_24_port, Y(23)
                           => mux_out_4_23_port, Y(22) => mux_out_4_22_port, 
                           Y(21) => mux_out_4_21_port, Y(20) => 
                           mux_out_4_20_port, Y(19) => mux_out_4_19_port, Y(18)
                           => mux_out_4_18_port, Y(17) => mux_out_4_17_port, 
                           Y(16) => mux_out_4_16_port, Y(15) => 
                           mux_out_4_15_port, Y(14) => mux_out_4_14_port, Y(13)
                           => mux_out_4_13_port, Y(12) => mux_out_4_12_port, 
                           Y(11) => mux_out_4_11_port, Y(10) => 
                           mux_out_4_10_port, Y(9) => mux_out_4_9_port, Y(8) =>
                           mux_out_4_8_port, Y(7) => mux_out_4_7_port, Y(6) => 
                           mux_out_4_6_port, Y(5) => mux_out_4_5_port, Y(4) => 
                           mux_out_4_4_port, Y(3) => mux_out_4_3_port, Y(2) => 
                           mux_out_4_2_port, Y(1) => mux_out_4_1_port, Y(0) => 
                           mux_out_4_0_port);
   MUX_I_5 : MUX5to1_NBIT32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => A(15), B(24) => A(14), B(23)
                           => A(13), B(22) => A(12), B(21) => A(11), B(20) => 
                           A(10), B(19) => A(9), B(18) => A(8), B(17) => A(7), 
                           B(16) => A(6), B(15) => A(5), B(14) => A(4), B(13) 
                           => A(3), B(12) => A(2), B(11) => A(1), B(10) => n21,
                           B(9) => X_Logic0_port, B(8) => X_Logic0_port, B(7) 
                           => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n13, 
                           C(30) => n13, C(29) => n13, C(28) => n13, C(27) => 
                           n13, C(26) => n13, C(25) => A_neg_10_25_port, C(24) 
                           => A_neg_10_24_port, C(23) => A_neg_10_23_port, 
                           C(22) => A_neg_10_22_port, C(21) => A_neg_10_21_port
                           , C(20) => A_neg_10_20_port, C(19) => 
                           A_neg_10_19_port, C(18) => A_neg_10_18_port, C(17) 
                           => A_neg_10_17_port, C(16) => A_neg_10_16_port, 
                           C(15) => A_neg_10_15_port, C(14) => A_neg_10_14_port
                           , C(13) => A_neg_10_13_port, C(12) => 
                           A_neg_10_12_port, C(11) => A_neg_10_11_port, C(10) 
                           => n21, C(9) => n70, C(8) => n70, C(7) => n70, C(6) 
                           => n70, C(5) => n70, C(4) => n70, C(3) => n70, C(2) 
                           => n70, C(1) => n70, C(0) => n70, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => A(15), D(25) => A(14), D(24)
                           => A(13), D(23) => A(12), D(22) => A(11), D(21) => 
                           A(10), D(20) => A(9), D(19) => A(8), D(18) => A(7), 
                           D(17) => A(6), D(16) => A(5), D(15) => A(4), D(14) 
                           => A(3), D(13) => A(2), D(12) => A(1), D(11) => A(0)
                           , D(10) => X_Logic0_port, D(9) => X_Logic0_port, 
                           D(8) => X_Logic0_port, D(7) => X_Logic0_port, D(6) 
                           => X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n14, E(30) => n14, E(29) => 
                           n14, E(28) => n14, E(27) => n14, E(26) => 
                           A_neg_11_26_port, E(25) => A_neg_11_25_port, E(24) 
                           => A_neg_11_24_port, E(23) => A_neg_11_23_port, 
                           E(22) => A_neg_11_22_port, E(21) => A_neg_11_21_port
                           , E(20) => A_neg_11_20_port, E(19) => 
                           A_neg_11_19_port, E(18) => A_neg_11_18_port, E(17) 
                           => A_neg_11_17_port, E(16) => A_neg_11_16_port, 
                           E(15) => A_neg_11_15_port, E(14) => A_neg_11_14_port
                           , E(13) => A_neg_11_13_port, E(12) => 
                           A_neg_11_12_port, E(11) => A(0), E(10) => n70, E(9) 
                           => n70, E(8) => n70, E(7) => n70, E(6) => n70, E(5) 
                           => n70, E(4) => n70, E(3) => n70, E(2) => n70, E(1) 
                           => n70, E(0) => n70, SEL(2) => selector_17_port, 
                           SEL(1) => selector_16_port, SEL(0) => 
                           selector_15_port, Y(31) => mux_out_5_31_port, Y(30) 
                           => mux_out_5_30_port, Y(29) => mux_out_5_29_port, 
                           Y(28) => mux_out_5_28_port, Y(27) => 
                           mux_out_5_27_port, Y(26) => mux_out_5_26_port, Y(25)
                           => mux_out_5_25_port, Y(24) => mux_out_5_24_port, 
                           Y(23) => mux_out_5_23_port, Y(22) => 
                           mux_out_5_22_port, Y(21) => mux_out_5_21_port, Y(20)
                           => mux_out_5_20_port, Y(19) => mux_out_5_19_port, 
                           Y(18) => mux_out_5_18_port, Y(17) => 
                           mux_out_5_17_port, Y(16) => mux_out_5_16_port, Y(15)
                           => mux_out_5_15_port, Y(14) => mux_out_5_14_port, 
                           Y(13) => mux_out_5_13_port, Y(12) => 
                           mux_out_5_12_port, Y(11) => mux_out_5_11_port, Y(10)
                           => mux_out_5_10_port, Y(9) => mux_out_5_9_port, Y(8)
                           => mux_out_5_8_port, Y(7) => mux_out_5_7_port, Y(6) 
                           => mux_out_5_6_port, Y(5) => mux_out_5_5_port, Y(4) 
                           => mux_out_5_4_port, Y(3) => mux_out_5_3_port, Y(2) 
                           => mux_out_5_2_port, Y(1) => mux_out_5_1_port, Y(0) 
                           => mux_out_5_0_port);
   MUX_I_6 : MUX5to1_NBIT32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => A(15), B(26) => A(14), B(25)
                           => A(13), B(24) => A(12), B(23) => A(11), B(22) => 
                           A(10), B(21) => A(9), B(20) => A(8), B(19) => A(7), 
                           B(18) => A(6), B(17) => A(5), B(16) => A(4), B(15) 
                           => A(3), B(14) => A(2), B(13) => A(1), B(12) => n21,
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n15, 
                           C(30) => n15, C(29) => n15, C(28) => n15, C(27) => 
                           A_neg_12_27_port, C(26) => A_neg_12_26_port, C(25) 
                           => A_neg_12_25_port, C(24) => A_neg_12_24_port, 
                           C(23) => A_neg_12_23_port, C(22) => A_neg_12_22_port
                           , C(21) => A_neg_12_21_port, C(20) => 
                           A_neg_12_20_port, C(19) => A_neg_12_19_port, C(18) 
                           => A_neg_12_18_port, C(17) => A_neg_12_17_port, 
                           C(16) => A_neg_12_16_port, C(15) => A_neg_12_15_port
                           , C(14) => A_neg_12_14_port, C(13) => 
                           A_neg_12_13_port, C(12) => n21, C(11) => n70, C(10) 
                           => n70, C(9) => n70, C(8) => n70, C(7) => n70, C(6) 
                           => n70, C(5) => n70, C(4) => n70, C(3) => n70, C(2) 
                           => n70, C(1) => n70, C(0) => n70, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => A(15), D(27) => A(14), D(26)
                           => A(13), D(25) => A(12), D(24) => A(11), D(23) => 
                           A(10), D(22) => A(9), D(21) => A(8), D(20) => A(7), 
                           D(19) => A(6), D(18) => A(5), D(17) => A(4), D(16) 
                           => A(3), D(15) => A(2), D(14) => A(1), D(13) => A(0)
                           , D(12) => X_Logic0_port, D(11) => X_Logic0_port, 
                           D(10) => X_Logic0_port, D(9) => X_Logic0_port, D(8) 
                           => X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n16, E(30) => n16, E(29) => 
                           n16, E(28) => A_neg_13_28_port, E(27) => 
                           A_neg_13_27_port, E(26) => A_neg_13_26_port, E(25) 
                           => A_neg_13_25_port, E(24) => A_neg_13_24_port, 
                           E(23) => A_neg_13_23_port, E(22) => A_neg_13_22_port
                           , E(21) => A_neg_13_21_port, E(20) => 
                           A_neg_13_20_port, E(19) => A_neg_13_19_port, E(18) 
                           => A_neg_13_18_port, E(17) => A_neg_13_17_port, 
                           E(16) => A_neg_13_16_port, E(15) => A_neg_13_15_port
                           , E(14) => A_neg_13_14_port, E(13) => n21, E(12) => 
                           n70, E(11) => n70, E(10) => n70, E(9) => n70, E(8) 
                           => n70, E(7) => n70, E(6) => n70, E(5) => n70, E(4) 
                           => n70, E(3) => n70, E(2) => n70, E(1) => n70, E(0) 
                           => n70, SEL(2) => selector_20_port, SEL(1) => 
                           selector_19_port, SEL(0) => selector_18_port, Y(31) 
                           => mux_out_6_31_port, Y(30) => mux_out_6_30_port, 
                           Y(29) => mux_out_6_29_port, Y(28) => 
                           mux_out_6_28_port, Y(27) => mux_out_6_27_port, Y(26)
                           => mux_out_6_26_port, Y(25) => mux_out_6_25_port, 
                           Y(24) => mux_out_6_24_port, Y(23) => 
                           mux_out_6_23_port, Y(22) => mux_out_6_22_port, Y(21)
                           => mux_out_6_21_port, Y(20) => mux_out_6_20_port, 
                           Y(19) => mux_out_6_19_port, Y(18) => 
                           mux_out_6_18_port, Y(17) => mux_out_6_17_port, Y(16)
                           => mux_out_6_16_port, Y(15) => mux_out_6_15_port, 
                           Y(14) => mux_out_6_14_port, Y(13) => 
                           mux_out_6_13_port, Y(12) => mux_out_6_12_port, Y(11)
                           => mux_out_6_11_port, Y(10) => mux_out_6_10_port, 
                           Y(9) => mux_out_6_9_port, Y(8) => mux_out_6_8_port, 
                           Y(7) => mux_out_6_7_port, Y(6) => mux_out_6_6_port, 
                           Y(5) => mux_out_6_5_port, Y(4) => mux_out_6_4_port, 
                           Y(3) => mux_out_6_3_port, Y(2) => mux_out_6_2_port, 
                           Y(1) => mux_out_6_1_port, Y(0) => mux_out_6_0_port);
   MUX_I_7 : MUX5to1_NBIT32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => A(15), B(28) => A(14), B(27)
                           => A(13), B(26) => A(12), B(25) => A(11), B(24) => 
                           A(10), B(23) => A(9), B(22) => A(8), B(21) => A(7), 
                           B(20) => A(6), B(19) => A(5), B(18) => A(4), B(17) 
                           => A(3), B(16) => A(2), B(15) => A(1), B(14) => n21,
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n17, 
                           C(30) => n17, C(29) => A_neg_14_29_port, C(28) => 
                           A_neg_14_28_port, C(27) => A_neg_14_27_port, C(26) 
                           => A_neg_14_26_port, C(25) => A_neg_14_25_port, 
                           C(24) => A_neg_14_24_port, C(23) => A_neg_14_23_port
                           , C(22) => A_neg_14_22_port, C(21) => 
                           A_neg_14_21_port, C(20) => A_neg_14_20_port, C(19) 
                           => A_neg_14_19_port, C(18) => A_neg_14_18_port, 
                           C(17) => A_neg_14_17_port, C(16) => A_neg_14_16_port
                           , C(15) => A_neg_14_15_port, C(14) => n21, C(13) => 
                           n70, C(12) => n70, C(11) => n70, C(10) => n70, C(9) 
                           => n70, C(8) => n70, C(7) => n70, C(6) => n70, C(5) 
                           => n70, C(4) => n70, C(3) => n70, C(2) => n70, C(1) 
                           => n70, C(0) => n70, D(31) => X_Logic0_port, D(30) 
                           => A(15), D(29) => A(14), D(28) => A(13), D(27) => 
                           A(12), D(26) => A(11), D(25) => A(10), D(24) => A(9)
                           , D(23) => A(8), D(22) => A(7), D(21) => A(6), D(20)
                           => A(5), D(19) => A(4), D(18) => A(3), D(17) => A(2)
                           , D(16) => A(1), D(15) => A(0), D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n1, E(30) => 
                           A_neg_15_30_port, E(29) => A_neg_15_29_port, E(28) 
                           => A_neg_15_28_port, E(27) => A_neg_15_27_port, 
                           E(26) => A_neg_15_26_port, E(25) => A_neg_15_25_port
                           , E(24) => A_neg_15_24_port, E(23) => 
                           A_neg_15_23_port, E(22) => A_neg_15_22_port, E(21) 
                           => A_neg_15_21_port, E(20) => A_neg_15_20_port, 
                           E(19) => A_neg_15_19_port, E(18) => A_neg_15_18_port
                           , E(17) => A_neg_15_17_port, E(16) => 
                           A_neg_15_16_port, E(15) => n21, E(14) => n70, E(13) 
                           => n70, E(12) => n70, E(11) => n70, E(10) => n70, 
                           E(9) => n70, E(8) => n70, E(7) => n70, E(6) => n70, 
                           E(5) => n70, E(4) => n70, E(3) => n70, E(2) => n70, 
                           E(1) => n70, E(0) => n70, SEL(2) => selector_23_port
                           , SEL(1) => selector_22_port, SEL(0) => 
                           selector_21_port, Y(31) => mux_out_7_31_port, Y(30) 
                           => mux_out_7_30_port, Y(29) => mux_out_7_29_port, 
                           Y(28) => mux_out_7_28_port, Y(27) => 
                           mux_out_7_27_port, Y(26) => mux_out_7_26_port, Y(25)
                           => mux_out_7_25_port, Y(24) => mux_out_7_24_port, 
                           Y(23) => mux_out_7_23_port, Y(22) => 
                           mux_out_7_22_port, Y(21) => mux_out_7_21_port, Y(20)
                           => mux_out_7_20_port, Y(19) => mux_out_7_19_port, 
                           Y(18) => mux_out_7_18_port, Y(17) => 
                           mux_out_7_17_port, Y(16) => mux_out_7_16_port, Y(15)
                           => mux_out_7_15_port, Y(14) => mux_out_7_14_port, 
                           Y(13) => mux_out_7_13_port, Y(12) => 
                           mux_out_7_12_port, Y(11) => mux_out_7_11_port, Y(10)
                           => mux_out_7_10_port, Y(9) => mux_out_7_9_port, Y(8)
                           => mux_out_7_8_port, Y(7) => mux_out_7_7_port, Y(6) 
                           => mux_out_7_6_port, Y(5) => mux_out_7_5_port, Y(4) 
                           => mux_out_7_4_port, Y(3) => mux_out_7_3_port, Y(2) 
                           => mux_out_7_2_port, Y(1) => mux_out_7_1_port, Y(0) 
                           => mux_out_7_0_port);
   ADD0 : ADDER_NBIT32_NBIT_PER_BLOCK4_7 port map( A(31) => addends_0_31_port, 
                           A(30) => addends_0_30_port, A(29) => 
                           addends_0_29_port, A(28) => addends_0_28_port, A(27)
                           => addends_0_27_port, A(26) => addends_0_26_port, 
                           A(25) => addends_0_25_port, A(24) => 
                           addends_0_24_port, A(23) => addends_0_23_port, A(22)
                           => addends_0_22_port, A(21) => addends_0_21_port, 
                           A(20) => addends_0_20_port, A(19) => 
                           addends_0_19_port, A(18) => addends_0_18_port, A(17)
                           => addends_0_17_port, A(16) => addends_0_16_port, 
                           A(15) => addends_0_15_port, A(14) => 
                           addends_0_14_port, A(13) => addends_0_13_port, A(12)
                           => addends_0_12_port, A(11) => addends_0_11_port, 
                           A(10) => addends_0_10_port, A(9) => addends_0_9_port
                           , A(8) => addends_0_8_port, A(7) => addends_0_7_port
                           , A(6) => addends_0_6_port, A(5) => addends_0_5_port
                           , A(4) => addends_0_4_port, A(3) => addends_0_3_port
                           , A(2) => addends_0_2_port, A(1) => addends_0_1_port
                           , A(0) => addends_0_0_port, B(31) => 
                           addends_1_31_port, B(30) => addends_1_30_port, B(29)
                           => addends_1_29_port, B(28) => addends_1_28_port, 
                           B(27) => addends_1_27_port, B(26) => 
                           addends_1_26_port, B(25) => addends_1_25_port, B(24)
                           => addends_1_24_port, B(23) => addends_1_23_port, 
                           B(22) => addends_1_22_port, B(21) => 
                           addends_1_21_port, B(20) => addends_1_20_port, B(19)
                           => addends_1_19_port, B(18) => addends_1_18_port, 
                           B(17) => addends_1_17_port, B(16) => 
                           addends_1_16_port, B(15) => addends_1_15_port, B(14)
                           => addends_1_14_port, B(13) => addends_1_13_port, 
                           B(12) => addends_1_12_port, B(11) => 
                           addends_1_11_port, B(10) => addends_1_10_port, B(9) 
                           => addends_1_9_port, B(8) => addends_1_8_port, B(7) 
                           => addends_1_7_port, B(6) => addends_1_6_port, B(5) 
                           => addends_1_5_port, B(4) => addends_1_4_port, B(3) 
                           => addends_1_3_port, B(2) => addends_1_2_port, B(1) 
                           => addends_1_1_port, B(0) => addends_1_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_0_31_port, S(30) => reg_in_0_30_port
                           , S(29) => reg_in_0_29_port, S(28) => 
                           reg_in_0_28_port, S(27) => reg_in_0_27_port, S(26) 
                           => reg_in_0_26_port, S(25) => reg_in_0_25_port, 
                           S(24) => reg_in_0_24_port, S(23) => reg_in_0_23_port
                           , S(22) => reg_in_0_22_port, S(21) => 
                           reg_in_0_21_port, S(20) => reg_in_0_20_port, S(19) 
                           => reg_in_0_19_port, S(18) => reg_in_0_18_port, 
                           S(17) => reg_in_0_17_port, S(16) => reg_in_0_16_port
                           , S(15) => reg_in_0_15_port, S(14) => 
                           reg_in_0_14_port, S(13) => reg_in_0_13_port, S(12) 
                           => reg_in_0_12_port, S(11) => reg_in_0_11_port, 
                           S(10) => reg_in_0_10_port, S(9) => reg_in_0_9_port, 
                           S(8) => reg_in_0_8_port, S(7) => reg_in_0_7_port, 
                           S(6) => reg_in_0_6_port, S(5) => reg_in_0_5_port, 
                           S(4) => reg_in_0_4_port, S(3) => reg_in_0_3_port, 
                           S(2) => reg_in_0_2_port, S(1) => reg_in_0_1_port, 
                           S(0) => reg_in_0_0_port, Cout => n_1687);
   REG0 : REG_NBIT32_3 port map( clk => CLOCK, reset => X_Logic0_port, enable 
                           => X_Logic1_port, data_in(31) => reg_in_0_31_port, 
                           data_in(30) => reg_in_0_30_port, data_in(29) => 
                           reg_in_0_29_port, data_in(28) => reg_in_0_28_port, 
                           data_in(27) => reg_in_0_27_port, data_in(26) => 
                           reg_in_0_26_port, data_in(25) => reg_in_0_25_port, 
                           data_in(24) => reg_in_0_24_port, data_in(23) => 
                           reg_in_0_23_port, data_in(22) => reg_in_0_22_port, 
                           data_in(21) => reg_in_0_21_port, data_in(20) => 
                           reg_in_0_20_port, data_in(19) => reg_in_0_19_port, 
                           data_in(18) => reg_in_0_18_port, data_in(17) => 
                           reg_in_0_17_port, data_in(16) => reg_in_0_16_port, 
                           data_in(15) => reg_in_0_15_port, data_in(14) => 
                           reg_in_0_14_port, data_in(13) => reg_in_0_13_port, 
                           data_in(12) => reg_in_0_12_port, data_in(11) => 
                           reg_in_0_11_port, data_in(10) => reg_in_0_10_port, 
                           data_in(9) => reg_in_0_9_port, data_in(8) => 
                           reg_in_0_8_port, data_in(7) => reg_in_0_7_port, 
                           data_in(6) => reg_in_0_6_port, data_in(5) => 
                           reg_in_0_5_port, data_in(4) => reg_in_0_4_port, 
                           data_in(3) => reg_in_0_3_port, data_in(2) => 
                           reg_in_0_2_port, data_in(1) => reg_in_0_1_port, 
                           data_in(0) => reg_in_0_0_port, data_out(31) => 
                           reg_out_0_31_port, data_out(30) => reg_out_0_30_port
                           , data_out(29) => reg_out_0_29_port, data_out(28) =>
                           reg_out_0_28_port, data_out(27) => reg_out_0_27_port
                           , data_out(26) => reg_out_0_26_port, data_out(25) =>
                           reg_out_0_25_port, data_out(24) => reg_out_0_24_port
                           , data_out(23) => reg_out_0_23_port, data_out(22) =>
                           reg_out_0_22_port, data_out(21) => reg_out_0_21_port
                           , data_out(20) => reg_out_0_20_port, data_out(19) =>
                           reg_out_0_19_port, data_out(18) => reg_out_0_18_port
                           , data_out(17) => reg_out_0_17_port, data_out(16) =>
                           reg_out_0_16_port, data_out(15) => reg_out_0_15_port
                           , data_out(14) => reg_out_0_14_port, data_out(13) =>
                           reg_out_0_13_port, data_out(12) => reg_out_0_12_port
                           , data_out(11) => reg_out_0_11_port, data_out(10) =>
                           reg_out_0_10_port, data_out(9) => reg_out_0_9_port, 
                           data_out(8) => reg_out_0_8_port, data_out(7) => 
                           reg_out_0_7_port, data_out(6) => reg_out_0_6_port, 
                           data_out(5) => reg_out_0_5_port, data_out(4) => 
                           reg_out_0_4_port, data_out(3) => reg_out_0_3_port, 
                           data_out(2) => reg_out_0_2_port, data_out(1) => 
                           reg_out_0_1_port, data_out(0) => reg_out_0_0_port);
   ADD_0i_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_6 port map( A(31) => 
                           reg_out_0_31_port, A(30) => reg_out_0_30_port, A(29)
                           => reg_out_0_29_port, A(28) => reg_out_0_28_port, 
                           A(27) => reg_out_0_27_port, A(26) => 
                           reg_out_0_26_port, A(25) => reg_out_0_25_port, A(24)
                           => reg_out_0_24_port, A(23) => reg_out_0_23_port, 
                           A(22) => reg_out_0_22_port, A(21) => 
                           reg_out_0_21_port, A(20) => reg_out_0_20_port, A(19)
                           => reg_out_0_19_port, A(18) => reg_out_0_18_port, 
                           A(17) => reg_out_0_17_port, A(16) => 
                           reg_out_0_16_port, A(15) => reg_out_0_15_port, A(14)
                           => reg_out_0_14_port, A(13) => reg_out_0_13_port, 
                           A(12) => reg_out_0_12_port, A(11) => 
                           reg_out_0_11_port, A(10) => reg_out_0_10_port, A(9) 
                           => reg_out_0_9_port, A(8) => reg_out_0_8_port, A(7) 
                           => reg_out_0_7_port, A(6) => reg_out_0_6_port, A(5) 
                           => reg_out_0_5_port, A(4) => reg_out_0_4_port, A(3) 
                           => reg_out_0_3_port, A(2) => reg_out_0_2_port, A(1) 
                           => reg_out_0_1_port, A(0) => reg_out_0_0_port, B(31)
                           => addends_2_31_port, B(30) => addends_2_30_port, 
                           B(29) => addends_2_29_port, B(28) => 
                           addends_2_28_port, B(27) => addends_2_27_port, B(26)
                           => addends_2_26_port, B(25) => addends_2_25_port, 
                           B(24) => addends_2_24_port, B(23) => 
                           addends_2_23_port, B(22) => addends_2_22_port, B(21)
                           => addends_2_21_port, B(20) => addends_2_20_port, 
                           B(19) => addends_2_19_port, B(18) => 
                           addends_2_18_port, B(17) => addends_2_17_port, B(16)
                           => addends_2_16_port, B(15) => addends_2_15_port, 
                           B(14) => addends_2_14_port, B(13) => 
                           addends_2_13_port, B(12) => addends_2_12_port, B(11)
                           => addends_2_11_port, B(10) => addends_2_10_port, 
                           B(9) => addends_2_9_port, B(8) => addends_2_8_port, 
                           B(7) => addends_2_7_port, B(6) => addends_2_6_port, 
                           B(5) => addends_2_5_port, B(4) => addends_2_4_port, 
                           B(3) => addends_2_3_port, B(2) => addends_2_2_port, 
                           B(1) => addends_2_1_port, B(0) => addends_2_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_0_31_port, S(30) => 
                           add_out_0_30_port, S(29) => add_out_0_29_port, S(28)
                           => add_out_0_28_port, S(27) => add_out_0_27_port, 
                           S(26) => add_out_0_26_port, S(25) => 
                           add_out_0_25_port, S(24) => add_out_0_24_port, S(23)
                           => add_out_0_23_port, S(22) => add_out_0_22_port, 
                           S(21) => add_out_0_21_port, S(20) => 
                           add_out_0_20_port, S(19) => add_out_0_19_port, S(18)
                           => add_out_0_18_port, S(17) => add_out_0_17_port, 
                           S(16) => add_out_0_16_port, S(15) => 
                           add_out_0_15_port, S(14) => add_out_0_14_port, S(13)
                           => add_out_0_13_port, S(12) => add_out_0_12_port, 
                           S(11) => add_out_0_11_port, S(10) => 
                           add_out_0_10_port, S(9) => add_out_0_9_port, S(8) =>
                           add_out_0_8_port, S(7) => add_out_0_7_port, S(6) => 
                           add_out_0_6_port, S(5) => add_out_0_5_port, S(4) => 
                           add_out_0_4_port, S(3) => add_out_0_3_port, S(2) => 
                           add_out_0_2_port, S(1) => add_out_0_1_port, S(0) => 
                           add_out_0_0_port, Cout => n_1688);
   ADD_1i_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_5 port map( A(31) => 
                           add_out_0_31_port, A(30) => add_out_0_30_port, A(29)
                           => add_out_0_29_port, A(28) => add_out_0_28_port, 
                           A(27) => add_out_0_27_port, A(26) => 
                           add_out_0_26_port, A(25) => add_out_0_25_port, A(24)
                           => add_out_0_24_port, A(23) => add_out_0_23_port, 
                           A(22) => add_out_0_22_port, A(21) => 
                           add_out_0_21_port, A(20) => add_out_0_20_port, A(19)
                           => add_out_0_19_port, A(18) => add_out_0_18_port, 
                           A(17) => add_out_0_17_port, A(16) => 
                           add_out_0_16_port, A(15) => add_out_0_15_port, A(14)
                           => add_out_0_14_port, A(13) => add_out_0_13_port, 
                           A(12) => add_out_0_12_port, A(11) => 
                           add_out_0_11_port, A(10) => add_out_0_10_port, A(9) 
                           => add_out_0_9_port, A(8) => add_out_0_8_port, A(7) 
                           => add_out_0_7_port, A(6) => add_out_0_6_port, A(5) 
                           => add_out_0_5_port, A(4) => add_out_0_4_port, A(3) 
                           => add_out_0_3_port, A(2) => add_out_0_2_port, A(1) 
                           => add_out_0_1_port, A(0) => add_out_0_0_port, B(31)
                           => addends_3_31_port, B(30) => addends_3_30_port, 
                           B(29) => addends_3_29_port, B(28) => 
                           addends_3_28_port, B(27) => addends_3_27_port, B(26)
                           => addends_3_26_port, B(25) => addends_3_25_port, 
                           B(24) => addends_3_24_port, B(23) => 
                           addends_3_23_port, B(22) => addends_3_22_port, B(21)
                           => addends_3_21_port, B(20) => addends_3_20_port, 
                           B(19) => addends_3_19_port, B(18) => 
                           addends_3_18_port, B(17) => addends_3_17_port, B(16)
                           => addends_3_16_port, B(15) => addends_3_15_port, 
                           B(14) => addends_3_14_port, B(13) => 
                           addends_3_13_port, B(12) => addends_3_12_port, B(11)
                           => addends_3_11_port, B(10) => addends_3_10_port, 
                           B(9) => addends_3_9_port, B(8) => addends_3_8_port, 
                           B(7) => addends_3_7_port, B(6) => addends_3_6_port, 
                           B(5) => addends_3_5_port, B(4) => addends_3_4_port, 
                           B(3) => addends_3_3_port, B(2) => addends_3_2_port, 
                           B(1) => addends_3_1_port, B(0) => addends_3_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_1_31_port, S(30) => reg_in_1_30_port
                           , S(29) => reg_in_1_29_port, S(28) => 
                           reg_in_1_28_port, S(27) => reg_in_1_27_port, S(26) 
                           => reg_in_1_26_port, S(25) => reg_in_1_25_port, 
                           S(24) => reg_in_1_24_port, S(23) => reg_in_1_23_port
                           , S(22) => reg_in_1_22_port, S(21) => 
                           reg_in_1_21_port, S(20) => reg_in_1_20_port, S(19) 
                           => reg_in_1_19_port, S(18) => reg_in_1_18_port, 
                           S(17) => reg_in_1_17_port, S(16) => reg_in_1_16_port
                           , S(15) => reg_in_1_15_port, S(14) => 
                           reg_in_1_14_port, S(13) => reg_in_1_13_port, S(12) 
                           => reg_in_1_12_port, S(11) => reg_in_1_11_port, 
                           S(10) => reg_in_1_10_port, S(9) => reg_in_1_9_port, 
                           S(8) => reg_in_1_8_port, S(7) => reg_in_1_7_port, 
                           S(6) => reg_in_1_6_port, S(5) => reg_in_1_5_port, 
                           S(4) => reg_in_1_4_port, S(3) => reg_in_1_3_port, 
                           S(2) => reg_in_1_2_port, S(1) => reg_in_1_1_port, 
                           S(0) => reg_in_1_0_port, Cout => n_1689);
   REG_i_1 : REG_NBIT32_2 port map( clk => CLOCK, reset => X_Logic0_port, 
                           enable => X_Logic1_port, data_in(31) => 
                           reg_in_1_31_port, data_in(30) => reg_in_1_30_port, 
                           data_in(29) => reg_in_1_29_port, data_in(28) => 
                           reg_in_1_28_port, data_in(27) => reg_in_1_27_port, 
                           data_in(26) => reg_in_1_26_port, data_in(25) => 
                           reg_in_1_25_port, data_in(24) => reg_in_1_24_port, 
                           data_in(23) => reg_in_1_23_port, data_in(22) => 
                           reg_in_1_22_port, data_in(21) => reg_in_1_21_port, 
                           data_in(20) => reg_in_1_20_port, data_in(19) => 
                           reg_in_1_19_port, data_in(18) => reg_in_1_18_port, 
                           data_in(17) => reg_in_1_17_port, data_in(16) => 
                           reg_in_1_16_port, data_in(15) => reg_in_1_15_port, 
                           data_in(14) => reg_in_1_14_port, data_in(13) => 
                           reg_in_1_13_port, data_in(12) => reg_in_1_12_port, 
                           data_in(11) => reg_in_1_11_port, data_in(10) => 
                           reg_in_1_10_port, data_in(9) => reg_in_1_9_port, 
                           data_in(8) => reg_in_1_8_port, data_in(7) => 
                           reg_in_1_7_port, data_in(6) => reg_in_1_6_port, 
                           data_in(5) => reg_in_1_5_port, data_in(4) => 
                           reg_in_1_4_port, data_in(3) => reg_in_1_3_port, 
                           data_in(2) => reg_in_1_2_port, data_in(1) => 
                           reg_in_1_1_port, data_in(0) => reg_in_1_0_port, 
                           data_out(31) => reg_out_1_31_port, data_out(30) => 
                           reg_out_1_30_port, data_out(29) => reg_out_1_29_port
                           , data_out(28) => reg_out_1_28_port, data_out(27) =>
                           reg_out_1_27_port, data_out(26) => reg_out_1_26_port
                           , data_out(25) => reg_out_1_25_port, data_out(24) =>
                           reg_out_1_24_port, data_out(23) => reg_out_1_23_port
                           , data_out(22) => reg_out_1_22_port, data_out(21) =>
                           reg_out_1_21_port, data_out(20) => reg_out_1_20_port
                           , data_out(19) => reg_out_1_19_port, data_out(18) =>
                           reg_out_1_18_port, data_out(17) => reg_out_1_17_port
                           , data_out(16) => reg_out_1_16_port, data_out(15) =>
                           reg_out_1_15_port, data_out(14) => reg_out_1_14_port
                           , data_out(13) => reg_out_1_13_port, data_out(12) =>
                           reg_out_1_12_port, data_out(11) => reg_out_1_11_port
                           , data_out(10) => reg_out_1_10_port, data_out(9) => 
                           reg_out_1_9_port, data_out(8) => reg_out_1_8_port, 
                           data_out(7) => reg_out_1_7_port, data_out(6) => 
                           reg_out_1_6_port, data_out(5) => reg_out_1_5_port, 
                           data_out(4) => reg_out_1_4_port, data_out(3) => 
                           reg_out_1_3_port, data_out(2) => reg_out_1_2_port, 
                           data_out(1) => reg_out_1_1_port, data_out(0) => 
                           reg_out_1_0_port);
   ADD_0i_2 : ADDER_NBIT32_NBIT_PER_BLOCK4_4 port map( A(31) => 
                           reg_out_1_31_port, A(30) => reg_out_1_30_port, A(29)
                           => reg_out_1_29_port, A(28) => reg_out_1_28_port, 
                           A(27) => reg_out_1_27_port, A(26) => 
                           reg_out_1_26_port, A(25) => reg_out_1_25_port, A(24)
                           => reg_out_1_24_port, A(23) => reg_out_1_23_port, 
                           A(22) => reg_out_1_22_port, A(21) => 
                           reg_out_1_21_port, A(20) => reg_out_1_20_port, A(19)
                           => reg_out_1_19_port, A(18) => reg_out_1_18_port, 
                           A(17) => reg_out_1_17_port, A(16) => 
                           reg_out_1_16_port, A(15) => reg_out_1_15_port, A(14)
                           => reg_out_1_14_port, A(13) => reg_out_1_13_port, 
                           A(12) => reg_out_1_12_port, A(11) => 
                           reg_out_1_11_port, A(10) => reg_out_1_10_port, A(9) 
                           => reg_out_1_9_port, A(8) => reg_out_1_8_port, A(7) 
                           => reg_out_1_7_port, A(6) => reg_out_1_6_port, A(5) 
                           => reg_out_1_5_port, A(4) => reg_out_1_4_port, A(3) 
                           => reg_out_1_3_port, A(2) => reg_out_1_2_port, A(1) 
                           => reg_out_1_1_port, A(0) => reg_out_1_0_port, B(31)
                           => addends_4_31_port, B(30) => addends_4_30_port, 
                           B(29) => addends_4_29_port, B(28) => 
                           addends_4_28_port, B(27) => addends_4_27_port, B(26)
                           => addends_4_26_port, B(25) => addends_4_25_port, 
                           B(24) => addends_4_24_port, B(23) => 
                           addends_4_23_port, B(22) => addends_4_22_port, B(21)
                           => addends_4_21_port, B(20) => addends_4_20_port, 
                           B(19) => addends_4_19_port, B(18) => 
                           addends_4_18_port, B(17) => addends_4_17_port, B(16)
                           => addends_4_16_port, B(15) => addends_4_15_port, 
                           B(14) => addends_4_14_port, B(13) => 
                           addends_4_13_port, B(12) => addends_4_12_port, B(11)
                           => addends_4_11_port, B(10) => addends_4_10_port, 
                           B(9) => addends_4_9_port, B(8) => addends_4_8_port, 
                           B(7) => addends_4_7_port, B(6) => addends_4_6_port, 
                           B(5) => addends_4_5_port, B(4) => addends_4_4_port, 
                           B(3) => addends_4_3_port, B(2) => addends_4_2_port, 
                           B(1) => addends_4_1_port, B(0) => addends_4_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_1_31_port, S(30) => 
                           add_out_1_30_port, S(29) => add_out_1_29_port, S(28)
                           => add_out_1_28_port, S(27) => add_out_1_27_port, 
                           S(26) => add_out_1_26_port, S(25) => 
                           add_out_1_25_port, S(24) => add_out_1_24_port, S(23)
                           => add_out_1_23_port, S(22) => add_out_1_22_port, 
                           S(21) => add_out_1_21_port, S(20) => 
                           add_out_1_20_port, S(19) => add_out_1_19_port, S(18)
                           => add_out_1_18_port, S(17) => add_out_1_17_port, 
                           S(16) => add_out_1_16_port, S(15) => 
                           add_out_1_15_port, S(14) => add_out_1_14_port, S(13)
                           => add_out_1_13_port, S(12) => add_out_1_12_port, 
                           S(11) => add_out_1_11_port, S(10) => 
                           add_out_1_10_port, S(9) => add_out_1_9_port, S(8) =>
                           add_out_1_8_port, S(7) => add_out_1_7_port, S(6) => 
                           add_out_1_6_port, S(5) => add_out_1_5_port, S(4) => 
                           add_out_1_4_port, S(3) => add_out_1_3_port, S(2) => 
                           add_out_1_2_port, S(1) => add_out_1_1_port, S(0) => 
                           add_out_1_0_port, Cout => n_1690);
   ADD_1i_2 : ADDER_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => 
                           add_out_1_31_port, A(30) => add_out_1_30_port, A(29)
                           => add_out_1_29_port, A(28) => add_out_1_28_port, 
                           A(27) => add_out_1_27_port, A(26) => 
                           add_out_1_26_port, A(25) => add_out_1_25_port, A(24)
                           => add_out_1_24_port, A(23) => add_out_1_23_port, 
                           A(22) => add_out_1_22_port, A(21) => 
                           add_out_1_21_port, A(20) => add_out_1_20_port, A(19)
                           => add_out_1_19_port, A(18) => add_out_1_18_port, 
                           A(17) => add_out_1_17_port, A(16) => 
                           add_out_1_16_port, A(15) => add_out_1_15_port, A(14)
                           => add_out_1_14_port, A(13) => add_out_1_13_port, 
                           A(12) => add_out_1_12_port, A(11) => 
                           add_out_1_11_port, A(10) => add_out_1_10_port, A(9) 
                           => add_out_1_9_port, A(8) => add_out_1_8_port, A(7) 
                           => add_out_1_7_port, A(6) => add_out_1_6_port, A(5) 
                           => add_out_1_5_port, A(4) => add_out_1_4_port, A(3) 
                           => add_out_1_3_port, A(2) => add_out_1_2_port, A(1) 
                           => add_out_1_1_port, A(0) => add_out_1_0_port, B(31)
                           => addends_5_31_port, B(30) => addends_5_30_port, 
                           B(29) => addends_5_29_port, B(28) => 
                           addends_5_28_port, B(27) => addends_5_27_port, B(26)
                           => addends_5_26_port, B(25) => addends_5_25_port, 
                           B(24) => addends_5_24_port, B(23) => 
                           addends_5_23_port, B(22) => addends_5_22_port, B(21)
                           => addends_5_21_port, B(20) => addends_5_20_port, 
                           B(19) => addends_5_19_port, B(18) => 
                           addends_5_18_port, B(17) => addends_5_17_port, B(16)
                           => addends_5_16_port, B(15) => addends_5_15_port, 
                           B(14) => addends_5_14_port, B(13) => 
                           addends_5_13_port, B(12) => addends_5_12_port, B(11)
                           => addends_5_11_port, B(10) => addends_5_10_port, 
                           B(9) => addends_5_9_port, B(8) => addends_5_8_port, 
                           B(7) => addends_5_7_port, B(6) => addends_5_6_port, 
                           B(5) => addends_5_5_port, B(4) => addends_5_4_port, 
                           B(3) => addends_5_3_port, B(2) => addends_5_2_port, 
                           B(1) => addends_5_1_port, B(0) => addends_5_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_2_31_port, S(30) => reg_in_2_30_port
                           , S(29) => reg_in_2_29_port, S(28) => 
                           reg_in_2_28_port, S(27) => reg_in_2_27_port, S(26) 
                           => reg_in_2_26_port, S(25) => reg_in_2_25_port, 
                           S(24) => reg_in_2_24_port, S(23) => reg_in_2_23_port
                           , S(22) => reg_in_2_22_port, S(21) => 
                           reg_in_2_21_port, S(20) => reg_in_2_20_port, S(19) 
                           => reg_in_2_19_port, S(18) => reg_in_2_18_port, 
                           S(17) => reg_in_2_17_port, S(16) => reg_in_2_16_port
                           , S(15) => reg_in_2_15_port, S(14) => 
                           reg_in_2_14_port, S(13) => reg_in_2_13_port, S(12) 
                           => reg_in_2_12_port, S(11) => reg_in_2_11_port, 
                           S(10) => reg_in_2_10_port, S(9) => reg_in_2_9_port, 
                           S(8) => reg_in_2_8_port, S(7) => reg_in_2_7_port, 
                           S(6) => reg_in_2_6_port, S(5) => reg_in_2_5_port, 
                           S(4) => reg_in_2_4_port, S(3) => reg_in_2_3_port, 
                           S(2) => reg_in_2_2_port, S(1) => reg_in_2_1_port, 
                           S(0) => reg_in_2_0_port, Cout => n_1691);
   REG_i_2 : REG_NBIT32_1 port map( clk => CLOCK, reset => X_Logic0_port, 
                           enable => X_Logic1_port, data_in(31) => 
                           reg_in_2_31_port, data_in(30) => reg_in_2_30_port, 
                           data_in(29) => reg_in_2_29_port, data_in(28) => 
                           reg_in_2_28_port, data_in(27) => reg_in_2_27_port, 
                           data_in(26) => reg_in_2_26_port, data_in(25) => 
                           reg_in_2_25_port, data_in(24) => reg_in_2_24_port, 
                           data_in(23) => reg_in_2_23_port, data_in(22) => 
                           reg_in_2_22_port, data_in(21) => reg_in_2_21_port, 
                           data_in(20) => reg_in_2_20_port, data_in(19) => 
                           reg_in_2_19_port, data_in(18) => reg_in_2_18_port, 
                           data_in(17) => reg_in_2_17_port, data_in(16) => 
                           reg_in_2_16_port, data_in(15) => reg_in_2_15_port, 
                           data_in(14) => reg_in_2_14_port, data_in(13) => 
                           reg_in_2_13_port, data_in(12) => reg_in_2_12_port, 
                           data_in(11) => reg_in_2_11_port, data_in(10) => 
                           reg_in_2_10_port, data_in(9) => reg_in_2_9_port, 
                           data_in(8) => reg_in_2_8_port, data_in(7) => 
                           reg_in_2_7_port, data_in(6) => reg_in_2_6_port, 
                           data_in(5) => reg_in_2_5_port, data_in(4) => 
                           reg_in_2_4_port, data_in(3) => reg_in_2_3_port, 
                           data_in(2) => reg_in_2_2_port, data_in(1) => 
                           reg_in_2_1_port, data_in(0) => reg_in_2_0_port, 
                           data_out(31) => reg_out_2_31_port, data_out(30) => 
                           reg_out_2_30_port, data_out(29) => reg_out_2_29_port
                           , data_out(28) => reg_out_2_28_port, data_out(27) =>
                           reg_out_2_27_port, data_out(26) => reg_out_2_26_port
                           , data_out(25) => reg_out_2_25_port, data_out(24) =>
                           reg_out_2_24_port, data_out(23) => reg_out_2_23_port
                           , data_out(22) => reg_out_2_22_port, data_out(21) =>
                           reg_out_2_21_port, data_out(20) => reg_out_2_20_port
                           , data_out(19) => reg_out_2_19_port, data_out(18) =>
                           reg_out_2_18_port, data_out(17) => reg_out_2_17_port
                           , data_out(16) => reg_out_2_16_port, data_out(15) =>
                           reg_out_2_15_port, data_out(14) => reg_out_2_14_port
                           , data_out(13) => reg_out_2_13_port, data_out(12) =>
                           reg_out_2_12_port, data_out(11) => reg_out_2_11_port
                           , data_out(10) => reg_out_2_10_port, data_out(9) => 
                           reg_out_2_9_port, data_out(8) => reg_out_2_8_port, 
                           data_out(7) => reg_out_2_7_port, data_out(6) => 
                           reg_out_2_6_port, data_out(5) => reg_out_2_5_port, 
                           data_out(4) => reg_out_2_4_port, data_out(3) => 
                           reg_out_2_3_port, data_out(2) => reg_out_2_2_port, 
                           data_out(1) => reg_out_2_1_port, data_out(0) => 
                           reg_out_2_0_port);
   ADD_N_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => 
                           reg_out_2_31_port, A(30) => reg_out_2_30_port, A(29)
                           => reg_out_2_29_port, A(28) => reg_out_2_28_port, 
                           A(27) => reg_out_2_27_port, A(26) => 
                           reg_out_2_26_port, A(25) => reg_out_2_25_port, A(24)
                           => reg_out_2_24_port, A(23) => reg_out_2_23_port, 
                           A(22) => reg_out_2_22_port, A(21) => 
                           reg_out_2_21_port, A(20) => reg_out_2_20_port, A(19)
                           => reg_out_2_19_port, A(18) => reg_out_2_18_port, 
                           A(17) => reg_out_2_17_port, A(16) => 
                           reg_out_2_16_port, A(15) => reg_out_2_15_port, A(14)
                           => reg_out_2_14_port, A(13) => reg_out_2_13_port, 
                           A(12) => reg_out_2_12_port, A(11) => 
                           reg_out_2_11_port, A(10) => reg_out_2_10_port, A(9) 
                           => reg_out_2_9_port, A(8) => reg_out_2_8_port, A(7) 
                           => reg_out_2_7_port, A(6) => reg_out_2_6_port, A(5) 
                           => reg_out_2_5_port, A(4) => reg_out_2_4_port, A(3) 
                           => reg_out_2_3_port, A(2) => reg_out_2_2_port, A(1) 
                           => reg_out_2_1_port, A(0) => reg_out_2_0_port, B(31)
                           => addends_6_31_port, B(30) => addends_6_30_port, 
                           B(29) => addends_6_29_port, B(28) => 
                           addends_6_28_port, B(27) => addends_6_27_port, B(26)
                           => addends_6_26_port, B(25) => addends_6_25_port, 
                           B(24) => addends_6_24_port, B(23) => 
                           addends_6_23_port, B(22) => addends_6_22_port, B(21)
                           => addends_6_21_port, B(20) => addends_6_20_port, 
                           B(19) => addends_6_19_port, B(18) => 
                           addends_6_18_port, B(17) => addends_6_17_port, B(16)
                           => addends_6_16_port, B(15) => addends_6_15_port, 
                           B(14) => addends_6_14_port, B(13) => 
                           addends_6_13_port, B(12) => addends_6_12_port, B(11)
                           => addends_6_11_port, B(10) => addends_6_10_port, 
                           B(9) => addends_6_9_port, B(8) => addends_6_8_port, 
                           B(7) => addends_6_7_port, B(6) => addends_6_6_port, 
                           B(5) => addends_6_5_port, B(4) => addends_6_4_port, 
                           B(3) => addends_6_3_port, B(2) => addends_6_2_port, 
                           B(1) => addends_6_1_port, B(0) => addends_6_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_2_31_port, S(30) => 
                           add_out_2_30_port, S(29) => add_out_2_29_port, S(28)
                           => add_out_2_28_port, S(27) => add_out_2_27_port, 
                           S(26) => add_out_2_26_port, S(25) => 
                           add_out_2_25_port, S(24) => add_out_2_24_port, S(23)
                           => add_out_2_23_port, S(22) => add_out_2_22_port, 
                           S(21) => add_out_2_21_port, S(20) => 
                           add_out_2_20_port, S(19) => add_out_2_19_port, S(18)
                           => add_out_2_18_port, S(17) => add_out_2_17_port, 
                           S(16) => add_out_2_16_port, S(15) => 
                           add_out_2_15_port, S(14) => add_out_2_14_port, S(13)
                           => add_out_2_13_port, S(12) => add_out_2_12_port, 
                           S(11) => add_out_2_11_port, S(10) => 
                           add_out_2_10_port, S(9) => add_out_2_9_port, S(8) =>
                           add_out_2_8_port, S(7) => add_out_2_7_port, S(6) => 
                           add_out_2_6_port, S(5) => add_out_2_5_port, S(4) => 
                           add_out_2_4_port, S(3) => add_out_2_3_port, S(2) => 
                           add_out_2_2_port, S(1) => add_out_2_1_port, S(0) => 
                           add_out_2_0_port, Cout => n_1692);
   ADD_N : ADDER_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => add_out_2_31_port,
                           A(30) => add_out_2_30_port, A(29) => 
                           add_out_2_29_port, A(28) => add_out_2_28_port, A(27)
                           => add_out_2_27_port, A(26) => add_out_2_26_port, 
                           A(25) => add_out_2_25_port, A(24) => 
                           add_out_2_24_port, A(23) => add_out_2_23_port, A(22)
                           => add_out_2_22_port, A(21) => add_out_2_21_port, 
                           A(20) => add_out_2_20_port, A(19) => 
                           add_out_2_19_port, A(18) => add_out_2_18_port, A(17)
                           => add_out_2_17_port, A(16) => add_out_2_16_port, 
                           A(15) => add_out_2_15_port, A(14) => 
                           add_out_2_14_port, A(13) => add_out_2_13_port, A(12)
                           => add_out_2_12_port, A(11) => add_out_2_11_port, 
                           A(10) => add_out_2_10_port, A(9) => add_out_2_9_port
                           , A(8) => add_out_2_8_port, A(7) => add_out_2_7_port
                           , A(6) => add_out_2_6_port, A(5) => add_out_2_5_port
                           , A(4) => add_out_2_4_port, A(3) => add_out_2_3_port
                           , A(2) => add_out_2_2_port, A(1) => add_out_2_1_port
                           , A(0) => add_out_2_0_port, B(31) => 
                           addends_7_31_port, B(30) => addends_7_30_port, B(29)
                           => addends_7_29_port, B(28) => addends_7_28_port, 
                           B(27) => addends_7_27_port, B(26) => 
                           addends_7_26_port, B(25) => addends_7_25_port, B(24)
                           => addends_7_24_port, B(23) => addends_7_23_port, 
                           B(22) => addends_7_22_port, B(21) => 
                           addends_7_21_port, B(20) => addends_7_20_port, B(19)
                           => addends_7_19_port, B(18) => addends_7_18_port, 
                           B(17) => addends_7_17_port, B(16) => 
                           addends_7_16_port, B(15) => addends_7_15_port, B(14)
                           => addends_7_14_port, B(13) => addends_7_13_port, 
                           B(12) => addends_7_12_port, B(11) => 
                           addends_7_11_port, B(10) => addends_7_10_port, B(9) 
                           => addends_7_9_port, B(8) => addends_7_8_port, B(7) 
                           => addends_7_7_port, B(6) => addends_7_6_port, B(5) 
                           => addends_7_5_port, B(4) => addends_7_4_port, B(3) 
                           => addends_7_3_port, B(2) => addends_7_2_port, B(1) 
                           => addends_7_1_port, B(0) => addends_7_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => Y(31), S(30) => Y(30), S(29) => Y(29), 
                           S(28) => Y(28), S(27) => Y(27), S(26) => Y(26), 
                           S(25) => Y(25), S(24) => Y(24), S(23) => Y(23), 
                           S(22) => Y(22), S(21) => Y(21), S(20) => Y(20), 
                           S(19) => Y(19), S(18) => Y(18), S(17) => Y(17), 
                           S(16) => Y(16), S(15) => Y(15), S(14) => Y(14), 
                           S(13) => Y(13), S(12) => Y(12), S(11) => Y(11), 
                           S(10) => Y(10), S(9) => Y(9), S(8) => Y(8), S(7) => 
                           Y(7), S(6) => Y(6), S(5) => Y(5), S(4) => Y(4), S(3)
                           => Y(3), S(2) => Y(2), S(1) => Y(1), S(0) => Y(0), 
                           Cout => n_1693);
   addends_reg_6_15_inst : DFF_X1 port map( D => pipe2_0_15_port, CK => CLOCK, 
                           Q => addends_6_15_port, QN => n_1694);
   addends_reg_6_6_inst : DFF_X1 port map( D => pipe2_0_6_port, CK => CLOCK, Q 
                           => addends_6_6_port, QN => n_1695);
   addends_reg_6_4_inst : DFF_X1 port map( D => pipe2_0_4_port, CK => CLOCK, Q 
                           => addends_6_4_port, QN => n_1696);
   addends_reg_6_1_inst : DFF_X1 port map( D => pipe2_0_1_port, CK => CLOCK, Q 
                           => addends_6_1_port, QN => n_1697);
   addends_reg_6_0_inst : DFF_X1 port map( D => pipe2_0_0_port, CK => CLOCK, Q 
                           => addends_6_0_port, QN => n_1698);
   addends_reg_5_31_inst : DFF_X1 port map( D => pipe1_1_31_port, CK => CLOCK, 
                           Q => addends_5_31_port, QN => n_1699);
   addends_reg_5_30_inst : DFF_X1 port map( D => pipe1_1_30_port, CK => CLOCK, 
                           Q => addends_5_30_port, QN => n_1700);
   addends_reg_5_29_inst : DFF_X1 port map( D => pipe1_1_29_port, CK => CLOCK, 
                           Q => addends_5_29_port, QN => n_1701);
   addends_reg_4_30_inst : DFF_X1 port map( D => pipe1_0_30_port, CK => CLOCK, 
                           Q => addends_4_30_port, QN => n_1702);
   addends_reg_5_4_inst : DFF_X1 port map( D => pipe1_1_4_port, CK => CLOCK, Q 
                           => addends_5_4_port, QN => n_1703);
   addends_reg_4_0_inst : SDFF_X1 port map( D => pipe1_0_0_port, SI => n2, SE 
                           => n2, CK => CLOCK, Q => addends_4_0_port, QN => 
                           n_1704);
   U3 : NAND2_X1 port map( A1 => sub_126_G16_carry_30_port, A2 => n67, ZN => n1
                           );
   n2 <= '0';
   U5 : BUF_X1 port map( A => n69, Z => n67);
   U6 : BUF_X1 port map( A => n27, Z => n25);
   U7 : BUF_X1 port map( A => n30, Z => n28);
   U8 : BUF_X1 port map( A => n33, Z => n31);
   U9 : BUF_X1 port map( A => n36, Z => n34);
   U10 : BUF_X1 port map( A => n39, Z => n37);
   U11 : BUF_X1 port map( A => n42, Z => n40);
   U12 : BUF_X1 port map( A => n45, Z => n43);
   U13 : BUF_X1 port map( A => n48, Z => n46);
   U14 : BUF_X1 port map( A => n51, Z => n49);
   U15 : BUF_X1 port map( A => n54, Z => n52);
   U16 : BUF_X1 port map( A => n57, Z => n55);
   U17 : BUF_X1 port map( A => n60, Z => n58);
   U18 : BUF_X1 port map( A => n63, Z => n61);
   U19 : BUF_X1 port map( A => n66, Z => n64);
   U20 : BUF_X1 port map( A => n24, Z => n22);
   U21 : BUF_X1 port map( A => n24, Z => n23);
   U22 : NAND2_X1 port map( A1 => sub_126_G6_carry_20_port, A2 => n68, ZN => n3
                           );
   U23 : NAND2_X1 port map( A1 => sub_126_G7_carry_21_port, A2 => n68, ZN => n4
                           );
   U24 : NAND2_X1 port map( A1 => sub_126_G8_carry_22_port, A2 => n68, ZN => n5
                           );
   U25 : NAND2_X1 port map( A1 => sub_126_carry_15_port, A2 => n67, ZN => n6);
   U26 : NAND2_X1 port map( A1 => sub_126_G9_carry_23_port, A2 => n68, ZN => n7
                           );
   U27 : NAND2_X1 port map( A1 => sub_126_G2_carry_16_port, A2 => n68, ZN => n8
                           );
   U28 : NAND2_X1 port map( A1 => sub_126_G3_carry_17_port, A2 => n68, ZN => n9
                           );
   U29 : NAND2_X1 port map( A1 => sub_126_G10_carry_24_port, A2 => n68, ZN => 
                           n10);
   U30 : NAND2_X1 port map( A1 => sub_126_G4_carry_18_port, A2 => n68, ZN => 
                           n11);
   U31 : NAND2_X1 port map( A1 => sub_126_G5_carry_19_port, A2 => n68, ZN => 
                           n12);
   U32 : NAND2_X1 port map( A1 => sub_126_G11_carry_25_port, A2 => n68, ZN => 
                           n13);
   U33 : NAND2_X1 port map( A1 => sub_126_G12_carry_26_port, A2 => n68, ZN => 
                           n14);
   U34 : NAND2_X1 port map( A1 => sub_126_G13_carry_27_port, A2 => n68, ZN => 
                           n15);
   U35 : NAND2_X1 port map( A1 => sub_126_G14_carry_28_port, A2 => n68, ZN => 
                           n16);
   U36 : NAND2_X1 port map( A1 => sub_126_G15_carry_29_port, A2 => n68, ZN => 
                           n17);
   U37 : INV_X1 port map( A => n22, ZN => n21);
   U38 : BUF_X1 port map( A => n23, Z => n18);
   U39 : BUF_X1 port map( A => n23, Z => n19);
   U40 : BUF_X1 port map( A => n23, Z => n20);
   U41 : BUF_X1 port map( A => n27, Z => n26);
   U42 : BUF_X1 port map( A => n30, Z => n29);
   U43 : BUF_X1 port map( A => n33, Z => n32);
   U44 : BUF_X1 port map( A => n36, Z => n35);
   U45 : BUF_X1 port map( A => n39, Z => n38);
   U46 : BUF_X1 port map( A => n42, Z => n41);
   U47 : BUF_X1 port map( A => n45, Z => n44);
   U48 : BUF_X1 port map( A => n48, Z => n47);
   U49 : BUF_X1 port map( A => n51, Z => n50);
   U50 : BUF_X1 port map( A => n54, Z => n53);
   U51 : BUF_X1 port map( A => n57, Z => n56);
   U52 : BUF_X1 port map( A => n60, Z => n59);
   U53 : BUF_X1 port map( A => n63, Z => n62);
   U54 : BUF_X1 port map( A => n66, Z => n65);
   U55 : BUF_X1 port map( A => n69, Z => n68);
   U56 : INV_X1 port map( A => A(0), ZN => n24);
   U57 : INV_X1 port map( A => A(1), ZN => n27);
   U58 : INV_X1 port map( A => A(2), ZN => n30);
   U59 : INV_X1 port map( A => A(3), ZN => n33);
   U60 : INV_X1 port map( A => A(4), ZN => n36);
   U61 : INV_X1 port map( A => A(5), ZN => n39);
   U62 : INV_X1 port map( A => A(6), ZN => n42);
   U63 : INV_X1 port map( A => A(7), ZN => n45);
   U64 : INV_X1 port map( A => A(8), ZN => n48);
   U65 : INV_X1 port map( A => A(9), ZN => n51);
   U66 : INV_X1 port map( A => A(10), ZN => n54);
   U67 : INV_X1 port map( A => A(11), ZN => n57);
   U68 : INV_X1 port map( A => A(12), ZN => n60);
   U69 : INV_X1 port map( A => A(13), ZN => n63);
   U70 : INV_X1 port map( A => A(14), ZN => n66);
   U71 : INV_X1 port map( A => A(15), ZN => n69);
   U72 : XOR2_X1 port map( A => n67, B => sub_126_G2_carry_16_port, Z => 
                           A_neg_1_16_port);
   U73 : AND2_X1 port map( A1 => sub_126_G2_carry_15_port, A2 => n65, ZN => 
                           sub_126_G2_carry_16_port);
   U74 : XOR2_X1 port map( A => n64, B => sub_126_G2_carry_15_port, Z => 
                           A_neg_1_15_port);
   U75 : AND2_X1 port map( A1 => sub_126_G2_carry_14_port, A2 => n62, ZN => 
                           sub_126_G2_carry_15_port);
   U76 : XOR2_X1 port map( A => n61, B => sub_126_G2_carry_14_port, Z => 
                           A_neg_1_14_port);
   U77 : AND2_X1 port map( A1 => sub_126_G2_carry_13_port, A2 => n59, ZN => 
                           sub_126_G2_carry_14_port);
   U78 : XOR2_X1 port map( A => n58, B => sub_126_G2_carry_13_port, Z => 
                           A_neg_1_13_port);
   U79 : AND2_X1 port map( A1 => sub_126_G2_carry_12_port, A2 => n56, ZN => 
                           sub_126_G2_carry_13_port);
   U80 : XOR2_X1 port map( A => n55, B => sub_126_G2_carry_12_port, Z => 
                           A_neg_1_12_port);
   U81 : AND2_X1 port map( A1 => sub_126_G2_carry_11_port, A2 => n53, ZN => 
                           sub_126_G2_carry_12_port);
   U82 : XOR2_X1 port map( A => n52, B => sub_126_G2_carry_11_port, Z => 
                           A_neg_1_11_port);
   U83 : AND2_X1 port map( A1 => sub_126_G2_carry_10_port, A2 => n50, ZN => 
                           sub_126_G2_carry_11_port);
   U84 : XOR2_X1 port map( A => n49, B => sub_126_G2_carry_10_port, Z => 
                           A_neg_1_10_port);
   U85 : AND2_X1 port map( A1 => sub_126_G2_carry_9_port, A2 => n47, ZN => 
                           sub_126_G2_carry_10_port);
   U86 : XOR2_X1 port map( A => n46, B => sub_126_G2_carry_9_port, Z => 
                           A_neg_1_9_port);
   U87 : AND2_X1 port map( A1 => sub_126_G2_carry_8_port, A2 => n44, ZN => 
                           sub_126_G2_carry_9_port);
   U88 : XOR2_X1 port map( A => n43, B => sub_126_G2_carry_8_port, Z => 
                           A_neg_1_8_port);
   U89 : AND2_X1 port map( A1 => sub_126_G2_carry_7_port, A2 => n41, ZN => 
                           sub_126_G2_carry_8_port);
   U90 : XOR2_X1 port map( A => n40, B => sub_126_G2_carry_7_port, Z => 
                           A_neg_1_7_port);
   U91 : AND2_X1 port map( A1 => sub_126_G2_carry_6_port, A2 => n38, ZN => 
                           sub_126_G2_carry_7_port);
   U92 : XOR2_X1 port map( A => n37, B => sub_126_G2_carry_6_port, Z => 
                           A_neg_1_6_port);
   U93 : AND2_X1 port map( A1 => sub_126_G2_carry_5_port, A2 => n35, ZN => 
                           sub_126_G2_carry_6_port);
   U94 : XOR2_X1 port map( A => n34, B => sub_126_G2_carry_5_port, Z => 
                           A_neg_1_5_port);
   U95 : AND2_X1 port map( A1 => sub_126_G2_carry_4_port, A2 => n32, ZN => 
                           sub_126_G2_carry_5_port);
   U96 : XOR2_X1 port map( A => n31, B => sub_126_G2_carry_4_port, Z => 
                           A_neg_1_4_port);
   U97 : AND2_X1 port map( A1 => sub_126_G2_carry_3_port, A2 => n29, ZN => 
                           sub_126_G2_carry_4_port);
   U98 : XOR2_X1 port map( A => n28, B => sub_126_G2_carry_3_port, Z => 
                           A_neg_1_3_port);
   U99 : AND2_X1 port map( A1 => n20, A2 => n26, ZN => sub_126_G2_carry_3_port)
                           ;
   U100 : XOR2_X1 port map( A => n25, B => n19, Z => A_neg_1_2_port);
   U101 : XOR2_X1 port map( A => n67, B => sub_126_carry_15_port, Z => 
                           A_neg_0_15_port);
   U102 : AND2_X1 port map( A1 => sub_126_carry_14_port, A2 => n64, ZN => 
                           sub_126_carry_15_port);
   U103 : XOR2_X1 port map( A => n64, B => sub_126_carry_14_port, Z => 
                           A_neg_0_14_port);
   U104 : AND2_X1 port map( A1 => sub_126_carry_13_port, A2 => n61, ZN => 
                           sub_126_carry_14_port);
   U105 : XOR2_X1 port map( A => n61, B => sub_126_carry_13_port, Z => 
                           A_neg_0_13_port);
   U106 : AND2_X1 port map( A1 => sub_126_carry_12_port, A2 => n58, ZN => 
                           sub_126_carry_13_port);
   U107 : XOR2_X1 port map( A => n58, B => sub_126_carry_12_port, Z => 
                           A_neg_0_12_port);
   U108 : AND2_X1 port map( A1 => sub_126_carry_11_port, A2 => n55, ZN => 
                           sub_126_carry_12_port);
   U109 : XOR2_X1 port map( A => n55, B => sub_126_carry_11_port, Z => 
                           A_neg_0_11_port);
   U110 : AND2_X1 port map( A1 => sub_126_carry_10_port, A2 => n52, ZN => 
                           sub_126_carry_11_port);
   U111 : XOR2_X1 port map( A => n52, B => sub_126_carry_10_port, Z => 
                           A_neg_0_10_port);
   U112 : AND2_X1 port map( A1 => sub_126_carry_9_port, A2 => n49, ZN => 
                           sub_126_carry_10_port);
   U113 : XOR2_X1 port map( A => n49, B => sub_126_carry_9_port, Z => 
                           A_neg_0_9_port);
   U114 : AND2_X1 port map( A1 => sub_126_carry_8_port, A2 => n46, ZN => 
                           sub_126_carry_9_port);
   U115 : XOR2_X1 port map( A => n46, B => sub_126_carry_8_port, Z => 
                           A_neg_0_8_port);
   U116 : AND2_X1 port map( A1 => sub_126_carry_7_port, A2 => n43, ZN => 
                           sub_126_carry_8_port);
   U117 : XOR2_X1 port map( A => n43, B => sub_126_carry_7_port, Z => 
                           A_neg_0_7_port);
   U118 : AND2_X1 port map( A1 => sub_126_carry_6_port, A2 => n40, ZN => 
                           sub_126_carry_7_port);
   U119 : XOR2_X1 port map( A => n40, B => sub_126_carry_6_port, Z => 
                           A_neg_0_6_port);
   U120 : AND2_X1 port map( A1 => sub_126_carry_5_port, A2 => n37, ZN => 
                           sub_126_carry_6_port);
   U121 : XOR2_X1 port map( A => n37, B => sub_126_carry_5_port, Z => 
                           A_neg_0_5_port);
   U122 : AND2_X1 port map( A1 => sub_126_carry_4_port, A2 => n34, ZN => 
                           sub_126_carry_5_port);
   U123 : XOR2_X1 port map( A => n34, B => sub_126_carry_4_port, Z => 
                           A_neg_0_4_port);
   U124 : AND2_X1 port map( A1 => sub_126_carry_3_port, A2 => n31, ZN => 
                           sub_126_carry_4_port);
   U125 : XOR2_X1 port map( A => n31, B => sub_126_carry_3_port, Z => 
                           A_neg_0_3_port);
   U126 : AND2_X1 port map( A1 => sub_126_carry_2_port, A2 => n28, ZN => 
                           sub_126_carry_3_port);
   U127 : XOR2_X1 port map( A => n28, B => sub_126_carry_2_port, Z => 
                           A_neg_0_2_port);
   U128 : AND2_X1 port map( A1 => n20, A2 => n25, ZN => sub_126_carry_2_port);
   U129 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_0_1_port);
   U130 : XOR2_X1 port map( A => n67, B => sub_126_G4_carry_18_port, Z => 
                           A_neg_3_18_port);
   U131 : AND2_X1 port map( A1 => sub_126_G4_carry_17_port, A2 => n65, ZN => 
                           sub_126_G4_carry_18_port);
   U132 : XOR2_X1 port map( A => n64, B => sub_126_G4_carry_17_port, Z => 
                           A_neg_3_17_port);
   U133 : AND2_X1 port map( A1 => sub_126_G4_carry_16_port, A2 => n62, ZN => 
                           sub_126_G4_carry_17_port);
   U134 : XOR2_X1 port map( A => n61, B => sub_126_G4_carry_16_port, Z => 
                           A_neg_3_16_port);
   U135 : AND2_X1 port map( A1 => sub_126_G4_carry_15_port, A2 => n59, ZN => 
                           sub_126_G4_carry_16_port);
   U136 : XOR2_X1 port map( A => n58, B => sub_126_G4_carry_15_port, Z => 
                           A_neg_3_15_port);
   U137 : AND2_X1 port map( A1 => sub_126_G4_carry_14_port, A2 => n56, ZN => 
                           sub_126_G4_carry_15_port);
   U138 : XOR2_X1 port map( A => n55, B => sub_126_G4_carry_14_port, Z => 
                           A_neg_3_14_port);
   U139 : AND2_X1 port map( A1 => sub_126_G4_carry_13_port, A2 => n53, ZN => 
                           sub_126_G4_carry_14_port);
   U140 : XOR2_X1 port map( A => n52, B => sub_126_G4_carry_13_port, Z => 
                           A_neg_3_13_port);
   U141 : AND2_X1 port map( A1 => sub_126_G4_carry_12_port, A2 => n50, ZN => 
                           sub_126_G4_carry_13_port);
   U142 : XOR2_X1 port map( A => n49, B => sub_126_G4_carry_12_port, Z => 
                           A_neg_3_12_port);
   U143 : AND2_X1 port map( A1 => sub_126_G4_carry_11_port, A2 => n47, ZN => 
                           sub_126_G4_carry_12_port);
   U144 : XOR2_X1 port map( A => n46, B => sub_126_G4_carry_11_port, Z => 
                           A_neg_3_11_port);
   U145 : AND2_X1 port map( A1 => sub_126_G4_carry_10_port, A2 => n44, ZN => 
                           sub_126_G4_carry_11_port);
   U146 : XOR2_X1 port map( A => n43, B => sub_126_G4_carry_10_port, Z => 
                           A_neg_3_10_port);
   U147 : AND2_X1 port map( A1 => sub_126_G4_carry_9_port, A2 => n41, ZN => 
                           sub_126_G4_carry_10_port);
   U148 : XOR2_X1 port map( A => n40, B => sub_126_G4_carry_9_port, Z => 
                           A_neg_3_9_port);
   U149 : AND2_X1 port map( A1 => sub_126_G4_carry_8_port, A2 => n38, ZN => 
                           sub_126_G4_carry_9_port);
   U150 : XOR2_X1 port map( A => n37, B => sub_126_G4_carry_8_port, Z => 
                           A_neg_3_8_port);
   U151 : AND2_X1 port map( A1 => sub_126_G4_carry_7_port, A2 => n35, ZN => 
                           sub_126_G4_carry_8_port);
   U152 : XOR2_X1 port map( A => n34, B => sub_126_G4_carry_7_port, Z => 
                           A_neg_3_7_port);
   U153 : AND2_X1 port map( A1 => sub_126_G4_carry_6_port, A2 => n32, ZN => 
                           sub_126_G4_carry_7_port);
   U154 : XOR2_X1 port map( A => n31, B => sub_126_G4_carry_6_port, Z => 
                           A_neg_3_6_port);
   U155 : AND2_X1 port map( A1 => sub_126_G4_carry_5_port, A2 => n29, ZN => 
                           sub_126_G4_carry_6_port);
   U156 : XOR2_X1 port map( A => n28, B => sub_126_G4_carry_5_port, Z => 
                           A_neg_3_5_port);
   U157 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => sub_126_G4_carry_5_port
                           );
   U158 : XOR2_X1 port map( A => n25, B => n19, Z => A_neg_3_4_port);
   U159 : XOR2_X1 port map( A => n67, B => sub_126_G3_carry_17_port, Z => 
                           A_neg_2_17_port);
   U160 : AND2_X1 port map( A1 => sub_126_G3_carry_16_port, A2 => n65, ZN => 
                           sub_126_G3_carry_17_port);
   U161 : XOR2_X1 port map( A => n64, B => sub_126_G3_carry_16_port, Z => 
                           A_neg_2_16_port);
   U162 : AND2_X1 port map( A1 => sub_126_G3_carry_15_port, A2 => n62, ZN => 
                           sub_126_G3_carry_16_port);
   U163 : XOR2_X1 port map( A => n61, B => sub_126_G3_carry_15_port, Z => 
                           A_neg_2_15_port);
   U164 : AND2_X1 port map( A1 => sub_126_G3_carry_14_port, A2 => n59, ZN => 
                           sub_126_G3_carry_15_port);
   U165 : XOR2_X1 port map( A => n58, B => sub_126_G3_carry_14_port, Z => 
                           A_neg_2_14_port);
   U166 : AND2_X1 port map( A1 => sub_126_G3_carry_13_port, A2 => n56, ZN => 
                           sub_126_G3_carry_14_port);
   U167 : XOR2_X1 port map( A => n55, B => sub_126_G3_carry_13_port, Z => 
                           A_neg_2_13_port);
   U168 : AND2_X1 port map( A1 => sub_126_G3_carry_12_port, A2 => n53, ZN => 
                           sub_126_G3_carry_13_port);
   U169 : XOR2_X1 port map( A => n52, B => sub_126_G3_carry_12_port, Z => 
                           A_neg_2_12_port);
   U170 : AND2_X1 port map( A1 => sub_126_G3_carry_11_port, A2 => n50, ZN => 
                           sub_126_G3_carry_12_port);
   U171 : XOR2_X1 port map( A => n49, B => sub_126_G3_carry_11_port, Z => 
                           A_neg_2_11_port);
   U172 : AND2_X1 port map( A1 => sub_126_G3_carry_10_port, A2 => n47, ZN => 
                           sub_126_G3_carry_11_port);
   U173 : XOR2_X1 port map( A => n46, B => sub_126_G3_carry_10_port, Z => 
                           A_neg_2_10_port);
   U174 : AND2_X1 port map( A1 => sub_126_G3_carry_9_port, A2 => n44, ZN => 
                           sub_126_G3_carry_10_port);
   U175 : XOR2_X1 port map( A => n43, B => sub_126_G3_carry_9_port, Z => 
                           A_neg_2_9_port);
   U176 : AND2_X1 port map( A1 => sub_126_G3_carry_8_port, A2 => n41, ZN => 
                           sub_126_G3_carry_9_port);
   U177 : XOR2_X1 port map( A => n40, B => sub_126_G3_carry_8_port, Z => 
                           A_neg_2_8_port);
   U178 : AND2_X1 port map( A1 => sub_126_G3_carry_7_port, A2 => n38, ZN => 
                           sub_126_G3_carry_8_port);
   U179 : XOR2_X1 port map( A => n37, B => sub_126_G3_carry_7_port, Z => 
                           A_neg_2_7_port);
   U180 : AND2_X1 port map( A1 => sub_126_G3_carry_6_port, A2 => n35, ZN => 
                           sub_126_G3_carry_7_port);
   U181 : XOR2_X1 port map( A => n34, B => sub_126_G3_carry_6_port, Z => 
                           A_neg_2_6_port);
   U182 : AND2_X1 port map( A1 => sub_126_G3_carry_5_port, A2 => n32, ZN => 
                           sub_126_G3_carry_6_port);
   U183 : XOR2_X1 port map( A => n31, B => sub_126_G3_carry_5_port, Z => 
                           A_neg_2_5_port);
   U184 : AND2_X1 port map( A1 => sub_126_G3_carry_4_port, A2 => n29, ZN => 
                           sub_126_G3_carry_5_port);
   U185 : XOR2_X1 port map( A => n28, B => sub_126_G3_carry_4_port, Z => 
                           A_neg_2_4_port);
   U186 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => sub_126_G3_carry_4_port
                           );
   U187 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_2_3_port);
   U188 : XOR2_X1 port map( A => n67, B => sub_126_G6_carry_20_port, Z => 
                           A_neg_5_20_port);
   U189 : AND2_X1 port map( A1 => sub_126_G6_carry_19_port, A2 => n65, ZN => 
                           sub_126_G6_carry_20_port);
   U190 : XOR2_X1 port map( A => n64, B => sub_126_G6_carry_19_port, Z => 
                           A_neg_5_19_port);
   U191 : AND2_X1 port map( A1 => sub_126_G6_carry_18_port, A2 => n62, ZN => 
                           sub_126_G6_carry_19_port);
   U192 : XOR2_X1 port map( A => n61, B => sub_126_G6_carry_18_port, Z => 
                           A_neg_5_18_port);
   U193 : AND2_X1 port map( A1 => sub_126_G6_carry_17_port, A2 => n59, ZN => 
                           sub_126_G6_carry_18_port);
   U194 : XOR2_X1 port map( A => n58, B => sub_126_G6_carry_17_port, Z => 
                           A_neg_5_17_port);
   U195 : AND2_X1 port map( A1 => sub_126_G6_carry_16_port, A2 => n56, ZN => 
                           sub_126_G6_carry_17_port);
   U196 : XOR2_X1 port map( A => n55, B => sub_126_G6_carry_16_port, Z => 
                           A_neg_5_16_port);
   U197 : AND2_X1 port map( A1 => sub_126_G6_carry_15_port, A2 => n53, ZN => 
                           sub_126_G6_carry_16_port);
   U198 : XOR2_X1 port map( A => n52, B => sub_126_G6_carry_15_port, Z => 
                           A_neg_5_15_port);
   U199 : AND2_X1 port map( A1 => sub_126_G6_carry_14_port, A2 => n50, ZN => 
                           sub_126_G6_carry_15_port);
   U200 : XOR2_X1 port map( A => n49, B => sub_126_G6_carry_14_port, Z => 
                           A_neg_5_14_port);
   U201 : AND2_X1 port map( A1 => sub_126_G6_carry_13_port, A2 => n47, ZN => 
                           sub_126_G6_carry_14_port);
   U202 : XOR2_X1 port map( A => n46, B => sub_126_G6_carry_13_port, Z => 
                           A_neg_5_13_port);
   U203 : AND2_X1 port map( A1 => sub_126_G6_carry_12_port, A2 => n44, ZN => 
                           sub_126_G6_carry_13_port);
   U204 : XOR2_X1 port map( A => n43, B => sub_126_G6_carry_12_port, Z => 
                           A_neg_5_12_port);
   U205 : AND2_X1 port map( A1 => sub_126_G6_carry_11_port, A2 => n41, ZN => 
                           sub_126_G6_carry_12_port);
   U206 : XOR2_X1 port map( A => n40, B => sub_126_G6_carry_11_port, Z => 
                           A_neg_5_11_port);
   U207 : AND2_X1 port map( A1 => sub_126_G6_carry_10_port, A2 => n38, ZN => 
                           sub_126_G6_carry_11_port);
   U208 : XOR2_X1 port map( A => n37, B => sub_126_G6_carry_10_port, Z => 
                           A_neg_5_10_port);
   U209 : AND2_X1 port map( A1 => sub_126_G6_carry_9_port, A2 => n35, ZN => 
                           sub_126_G6_carry_10_port);
   U210 : XOR2_X1 port map( A => n34, B => sub_126_G6_carry_9_port, Z => 
                           A_neg_5_9_port);
   U211 : AND2_X1 port map( A1 => sub_126_G6_carry_8_port, A2 => n32, ZN => 
                           sub_126_G6_carry_9_port);
   U212 : XOR2_X1 port map( A => n31, B => sub_126_G6_carry_8_port, Z => 
                           A_neg_5_8_port);
   U213 : AND2_X1 port map( A1 => sub_126_G6_carry_7_port, A2 => n29, ZN => 
                           sub_126_G6_carry_8_port);
   U214 : XOR2_X1 port map( A => n28, B => sub_126_G6_carry_7_port, Z => 
                           A_neg_5_7_port);
   U215 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => sub_126_G6_carry_7_port
                           );
   U216 : XOR2_X1 port map( A => n25, B => n19, Z => A_neg_5_6_port);
   U217 : XOR2_X1 port map( A => n67, B => sub_126_G5_carry_19_port, Z => 
                           A_neg_4_19_port);
   U218 : AND2_X1 port map( A1 => sub_126_G5_carry_18_port, A2 => n65, ZN => 
                           sub_126_G5_carry_19_port);
   U219 : XOR2_X1 port map( A => n64, B => sub_126_G5_carry_18_port, Z => 
                           A_neg_4_18_port);
   U220 : AND2_X1 port map( A1 => sub_126_G5_carry_17_port, A2 => n62, ZN => 
                           sub_126_G5_carry_18_port);
   U221 : XOR2_X1 port map( A => n61, B => sub_126_G5_carry_17_port, Z => 
                           A_neg_4_17_port);
   U222 : AND2_X1 port map( A1 => sub_126_G5_carry_16_port, A2 => n59, ZN => 
                           sub_126_G5_carry_17_port);
   U223 : XOR2_X1 port map( A => n58, B => sub_126_G5_carry_16_port, Z => 
                           A_neg_4_16_port);
   U224 : AND2_X1 port map( A1 => sub_126_G5_carry_15_port, A2 => n56, ZN => 
                           sub_126_G5_carry_16_port);
   U225 : XOR2_X1 port map( A => n55, B => sub_126_G5_carry_15_port, Z => 
                           A_neg_4_15_port);
   U226 : AND2_X1 port map( A1 => sub_126_G5_carry_14_port, A2 => n53, ZN => 
                           sub_126_G5_carry_15_port);
   U227 : XOR2_X1 port map( A => n52, B => sub_126_G5_carry_14_port, Z => 
                           A_neg_4_14_port);
   U228 : AND2_X1 port map( A1 => sub_126_G5_carry_13_port, A2 => n50, ZN => 
                           sub_126_G5_carry_14_port);
   U229 : XOR2_X1 port map( A => n49, B => sub_126_G5_carry_13_port, Z => 
                           A_neg_4_13_port);
   U230 : AND2_X1 port map( A1 => sub_126_G5_carry_12_port, A2 => n47, ZN => 
                           sub_126_G5_carry_13_port);
   U231 : XOR2_X1 port map( A => n46, B => sub_126_G5_carry_12_port, Z => 
                           A_neg_4_12_port);
   U232 : AND2_X1 port map( A1 => sub_126_G5_carry_11_port, A2 => n44, ZN => 
                           sub_126_G5_carry_12_port);
   U233 : XOR2_X1 port map( A => n43, B => sub_126_G5_carry_11_port, Z => 
                           A_neg_4_11_port);
   U234 : AND2_X1 port map( A1 => sub_126_G5_carry_10_port, A2 => n41, ZN => 
                           sub_126_G5_carry_11_port);
   U235 : XOR2_X1 port map( A => n40, B => sub_126_G5_carry_10_port, Z => 
                           A_neg_4_10_port);
   U236 : AND2_X1 port map( A1 => sub_126_G5_carry_9_port, A2 => n38, ZN => 
                           sub_126_G5_carry_10_port);
   U237 : XOR2_X1 port map( A => n37, B => sub_126_G5_carry_9_port, Z => 
                           A_neg_4_9_port);
   U238 : AND2_X1 port map( A1 => sub_126_G5_carry_8_port, A2 => n35, ZN => 
                           sub_126_G5_carry_9_port);
   U239 : XOR2_X1 port map( A => n34, B => sub_126_G5_carry_8_port, Z => 
                           A_neg_4_8_port);
   U240 : AND2_X1 port map( A1 => sub_126_G5_carry_7_port, A2 => n32, ZN => 
                           sub_126_G5_carry_8_port);
   U241 : XOR2_X1 port map( A => n31, B => sub_126_G5_carry_7_port, Z => 
                           A_neg_4_7_port);
   U242 : AND2_X1 port map( A1 => sub_126_G5_carry_6_port, A2 => n29, ZN => 
                           sub_126_G5_carry_7_port);
   U243 : XOR2_X1 port map( A => n28, B => sub_126_G5_carry_6_port, Z => 
                           A_neg_4_6_port);
   U244 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => sub_126_G5_carry_6_port
                           );
   U245 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_4_5_port);
   U246 : XOR2_X1 port map( A => n67, B => sub_126_G8_carry_22_port, Z => 
                           A_neg_7_22_port);
   U247 : AND2_X1 port map( A1 => sub_126_G8_carry_21_port, A2 => n65, ZN => 
                           sub_126_G8_carry_22_port);
   U248 : XOR2_X1 port map( A => n64, B => sub_126_G8_carry_21_port, Z => 
                           A_neg_7_21_port);
   U249 : AND2_X1 port map( A1 => sub_126_G8_carry_20_port, A2 => n62, ZN => 
                           sub_126_G8_carry_21_port);
   U250 : XOR2_X1 port map( A => n61, B => sub_126_G8_carry_20_port, Z => 
                           A_neg_7_20_port);
   U251 : AND2_X1 port map( A1 => sub_126_G8_carry_19_port, A2 => n59, ZN => 
                           sub_126_G8_carry_20_port);
   U252 : XOR2_X1 port map( A => n58, B => sub_126_G8_carry_19_port, Z => 
                           A_neg_7_19_port);
   U253 : AND2_X1 port map( A1 => sub_126_G8_carry_18_port, A2 => n56, ZN => 
                           sub_126_G8_carry_19_port);
   U254 : XOR2_X1 port map( A => n55, B => sub_126_G8_carry_18_port, Z => 
                           A_neg_7_18_port);
   U255 : AND2_X1 port map( A1 => sub_126_G8_carry_17_port, A2 => n53, ZN => 
                           sub_126_G8_carry_18_port);
   U256 : XOR2_X1 port map( A => n52, B => sub_126_G8_carry_17_port, Z => 
                           A_neg_7_17_port);
   U257 : AND2_X1 port map( A1 => sub_126_G8_carry_16_port, A2 => n50, ZN => 
                           sub_126_G8_carry_17_port);
   U258 : XOR2_X1 port map( A => n49, B => sub_126_G8_carry_16_port, Z => 
                           A_neg_7_16_port);
   U259 : AND2_X1 port map( A1 => sub_126_G8_carry_15_port, A2 => n47, ZN => 
                           sub_126_G8_carry_16_port);
   U260 : XOR2_X1 port map( A => n46, B => sub_126_G8_carry_15_port, Z => 
                           A_neg_7_15_port);
   U261 : AND2_X1 port map( A1 => sub_126_G8_carry_14_port, A2 => n44, ZN => 
                           sub_126_G8_carry_15_port);
   U262 : XOR2_X1 port map( A => n43, B => sub_126_G8_carry_14_port, Z => 
                           A_neg_7_14_port);
   U263 : AND2_X1 port map( A1 => sub_126_G8_carry_13_port, A2 => n41, ZN => 
                           sub_126_G8_carry_14_port);
   U264 : XOR2_X1 port map( A => n40, B => sub_126_G8_carry_13_port, Z => 
                           A_neg_7_13_port);
   U265 : AND2_X1 port map( A1 => sub_126_G8_carry_12_port, A2 => n38, ZN => 
                           sub_126_G8_carry_13_port);
   U266 : XOR2_X1 port map( A => n37, B => sub_126_G8_carry_12_port, Z => 
                           A_neg_7_12_port);
   U267 : AND2_X1 port map( A1 => sub_126_G8_carry_11_port, A2 => n35, ZN => 
                           sub_126_G8_carry_12_port);
   U268 : XOR2_X1 port map( A => n34, B => sub_126_G8_carry_11_port, Z => 
                           A_neg_7_11_port);
   U269 : AND2_X1 port map( A1 => sub_126_G8_carry_10_port, A2 => n32, ZN => 
                           sub_126_G8_carry_11_port);
   U270 : XOR2_X1 port map( A => n31, B => sub_126_G8_carry_10_port, Z => 
                           A_neg_7_10_port);
   U271 : AND2_X1 port map( A1 => sub_126_G8_carry_9_port, A2 => n29, ZN => 
                           sub_126_G8_carry_10_port);
   U272 : XOR2_X1 port map( A => n28, B => sub_126_G8_carry_9_port, Z => 
                           A_neg_7_9_port);
   U273 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => sub_126_G8_carry_9_port
                           );
   U274 : XOR2_X1 port map( A => n25, B => n19, Z => A_neg_7_8_port);
   U275 : XOR2_X1 port map( A => n67, B => sub_126_G7_carry_21_port, Z => 
                           A_neg_6_21_port);
   U276 : AND2_X1 port map( A1 => sub_126_G7_carry_20_port, A2 => n65, ZN => 
                           sub_126_G7_carry_21_port);
   U277 : XOR2_X1 port map( A => n64, B => sub_126_G7_carry_20_port, Z => 
                           A_neg_6_20_port);
   U278 : AND2_X1 port map( A1 => sub_126_G7_carry_19_port, A2 => n62, ZN => 
                           sub_126_G7_carry_20_port);
   U279 : XOR2_X1 port map( A => n61, B => sub_126_G7_carry_19_port, Z => 
                           A_neg_6_19_port);
   U280 : AND2_X1 port map( A1 => sub_126_G7_carry_18_port, A2 => n59, ZN => 
                           sub_126_G7_carry_19_port);
   U281 : XOR2_X1 port map( A => n58, B => sub_126_G7_carry_18_port, Z => 
                           A_neg_6_18_port);
   U282 : AND2_X1 port map( A1 => sub_126_G7_carry_17_port, A2 => n56, ZN => 
                           sub_126_G7_carry_18_port);
   U283 : XOR2_X1 port map( A => n55, B => sub_126_G7_carry_17_port, Z => 
                           A_neg_6_17_port);
   U284 : AND2_X1 port map( A1 => sub_126_G7_carry_16_port, A2 => n53, ZN => 
                           sub_126_G7_carry_17_port);
   U285 : XOR2_X1 port map( A => n52, B => sub_126_G7_carry_16_port, Z => 
                           A_neg_6_16_port);
   U286 : AND2_X1 port map( A1 => sub_126_G7_carry_15_port, A2 => n50, ZN => 
                           sub_126_G7_carry_16_port);
   U287 : XOR2_X1 port map( A => n49, B => sub_126_G7_carry_15_port, Z => 
                           A_neg_6_15_port);
   U288 : AND2_X1 port map( A1 => sub_126_G7_carry_14_port, A2 => n47, ZN => 
                           sub_126_G7_carry_15_port);
   U289 : XOR2_X1 port map( A => n46, B => sub_126_G7_carry_14_port, Z => 
                           A_neg_6_14_port);
   U290 : AND2_X1 port map( A1 => sub_126_G7_carry_13_port, A2 => n44, ZN => 
                           sub_126_G7_carry_14_port);
   U291 : XOR2_X1 port map( A => n43, B => sub_126_G7_carry_13_port, Z => 
                           A_neg_6_13_port);
   U292 : AND2_X1 port map( A1 => sub_126_G7_carry_12_port, A2 => n41, ZN => 
                           sub_126_G7_carry_13_port);
   U293 : XOR2_X1 port map( A => n40, B => sub_126_G7_carry_12_port, Z => 
                           A_neg_6_12_port);
   U294 : AND2_X1 port map( A1 => sub_126_G7_carry_11_port, A2 => n38, ZN => 
                           sub_126_G7_carry_12_port);
   U295 : XOR2_X1 port map( A => n37, B => sub_126_G7_carry_11_port, Z => 
                           A_neg_6_11_port);
   U296 : AND2_X1 port map( A1 => sub_126_G7_carry_10_port, A2 => n35, ZN => 
                           sub_126_G7_carry_11_port);
   U297 : XOR2_X1 port map( A => n34, B => sub_126_G7_carry_10_port, Z => 
                           A_neg_6_10_port);
   U298 : AND2_X1 port map( A1 => sub_126_G7_carry_9_port, A2 => n32, ZN => 
                           sub_126_G7_carry_10_port);
   U299 : XOR2_X1 port map( A => n31, B => sub_126_G7_carry_9_port, Z => 
                           A_neg_6_9_port);
   U300 : AND2_X1 port map( A1 => sub_126_G7_carry_8_port, A2 => n29, ZN => 
                           sub_126_G7_carry_9_port);
   U301 : XOR2_X1 port map( A => n28, B => sub_126_G7_carry_8_port, Z => 
                           A_neg_6_8_port);
   U302 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => sub_126_G7_carry_8_port
                           );
   U303 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_6_7_port);
   U304 : XOR2_X1 port map( A => n67, B => sub_126_G10_carry_24_port, Z => 
                           A_neg_9_24_port);
   U305 : AND2_X1 port map( A1 => sub_126_G10_carry_23_port, A2 => n65, ZN => 
                           sub_126_G10_carry_24_port);
   U306 : XOR2_X1 port map( A => n64, B => sub_126_G10_carry_23_port, Z => 
                           A_neg_9_23_port);
   U307 : AND2_X1 port map( A1 => sub_126_G10_carry_22_port, A2 => n62, ZN => 
                           sub_126_G10_carry_23_port);
   U308 : XOR2_X1 port map( A => n61, B => sub_126_G10_carry_22_port, Z => 
                           A_neg_9_22_port);
   U309 : AND2_X1 port map( A1 => sub_126_G10_carry_21_port, A2 => n59, ZN => 
                           sub_126_G10_carry_22_port);
   U310 : XOR2_X1 port map( A => n58, B => sub_126_G10_carry_21_port, Z => 
                           A_neg_9_21_port);
   U311 : AND2_X1 port map( A1 => sub_126_G10_carry_20_port, A2 => n56, ZN => 
                           sub_126_G10_carry_21_port);
   U312 : XOR2_X1 port map( A => n55, B => sub_126_G10_carry_20_port, Z => 
                           A_neg_9_20_port);
   U313 : AND2_X1 port map( A1 => sub_126_G10_carry_19_port, A2 => n53, ZN => 
                           sub_126_G10_carry_20_port);
   U314 : XOR2_X1 port map( A => n52, B => sub_126_G10_carry_19_port, Z => 
                           A_neg_9_19_port);
   U315 : AND2_X1 port map( A1 => sub_126_G10_carry_18_port, A2 => n50, ZN => 
                           sub_126_G10_carry_19_port);
   U316 : XOR2_X1 port map( A => n49, B => sub_126_G10_carry_18_port, Z => 
                           A_neg_9_18_port);
   U317 : AND2_X1 port map( A1 => sub_126_G10_carry_17_port, A2 => n47, ZN => 
                           sub_126_G10_carry_18_port);
   U318 : XOR2_X1 port map( A => n46, B => sub_126_G10_carry_17_port, Z => 
                           A_neg_9_17_port);
   U319 : AND2_X1 port map( A1 => sub_126_G10_carry_16_port, A2 => n44, ZN => 
                           sub_126_G10_carry_17_port);
   U320 : XOR2_X1 port map( A => n43, B => sub_126_G10_carry_16_port, Z => 
                           A_neg_9_16_port);
   U321 : AND2_X1 port map( A1 => sub_126_G10_carry_15_port, A2 => n41, ZN => 
                           sub_126_G10_carry_16_port);
   U322 : XOR2_X1 port map( A => n40, B => sub_126_G10_carry_15_port, Z => 
                           A_neg_9_15_port);
   U323 : AND2_X1 port map( A1 => sub_126_G10_carry_14_port, A2 => n38, ZN => 
                           sub_126_G10_carry_15_port);
   U324 : XOR2_X1 port map( A => n37, B => sub_126_G10_carry_14_port, Z => 
                           A_neg_9_14_port);
   U325 : AND2_X1 port map( A1 => sub_126_G10_carry_13_port, A2 => n35, ZN => 
                           sub_126_G10_carry_14_port);
   U326 : XOR2_X1 port map( A => n34, B => sub_126_G10_carry_13_port, Z => 
                           A_neg_9_13_port);
   U327 : AND2_X1 port map( A1 => sub_126_G10_carry_12_port, A2 => n32, ZN => 
                           sub_126_G10_carry_13_port);
   U328 : XOR2_X1 port map( A => n31, B => sub_126_G10_carry_12_port, Z => 
                           A_neg_9_12_port);
   U329 : AND2_X1 port map( A1 => sub_126_G10_carry_11_port, A2 => n29, ZN => 
                           sub_126_G10_carry_12_port);
   U330 : XOR2_X1 port map( A => n28, B => sub_126_G10_carry_11_port, Z => 
                           A_neg_9_11_port);
   U331 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G10_carry_11_port);
   U332 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_9_10_port);
   U333 : XOR2_X1 port map( A => n67, B => sub_126_G9_carry_23_port, Z => 
                           A_neg_8_23_port);
   U334 : AND2_X1 port map( A1 => sub_126_G9_carry_22_port, A2 => n65, ZN => 
                           sub_126_G9_carry_23_port);
   U335 : XOR2_X1 port map( A => n64, B => sub_126_G9_carry_22_port, Z => 
                           A_neg_8_22_port);
   U336 : AND2_X1 port map( A1 => sub_126_G9_carry_21_port, A2 => n62, ZN => 
                           sub_126_G9_carry_22_port);
   U337 : XOR2_X1 port map( A => n61, B => sub_126_G9_carry_21_port, Z => 
                           A_neg_8_21_port);
   U338 : AND2_X1 port map( A1 => sub_126_G9_carry_20_port, A2 => n59, ZN => 
                           sub_126_G9_carry_21_port);
   U339 : XOR2_X1 port map( A => n58, B => sub_126_G9_carry_20_port, Z => 
                           A_neg_8_20_port);
   U340 : AND2_X1 port map( A1 => sub_126_G9_carry_19_port, A2 => n56, ZN => 
                           sub_126_G9_carry_20_port);
   U341 : XOR2_X1 port map( A => n55, B => sub_126_G9_carry_19_port, Z => 
                           A_neg_8_19_port);
   U342 : AND2_X1 port map( A1 => sub_126_G9_carry_18_port, A2 => n53, ZN => 
                           sub_126_G9_carry_19_port);
   U343 : XOR2_X1 port map( A => n52, B => sub_126_G9_carry_18_port, Z => 
                           A_neg_8_18_port);
   U344 : AND2_X1 port map( A1 => sub_126_G9_carry_17_port, A2 => n50, ZN => 
                           sub_126_G9_carry_18_port);
   U345 : XOR2_X1 port map( A => n49, B => sub_126_G9_carry_17_port, Z => 
                           A_neg_8_17_port);
   U346 : AND2_X1 port map( A1 => sub_126_G9_carry_16_port, A2 => n47, ZN => 
                           sub_126_G9_carry_17_port);
   U347 : XOR2_X1 port map( A => n46, B => sub_126_G9_carry_16_port, Z => 
                           A_neg_8_16_port);
   U348 : AND2_X1 port map( A1 => sub_126_G9_carry_15_port, A2 => n44, ZN => 
                           sub_126_G9_carry_16_port);
   U349 : XOR2_X1 port map( A => n43, B => sub_126_G9_carry_15_port, Z => 
                           A_neg_8_15_port);
   U350 : AND2_X1 port map( A1 => sub_126_G9_carry_14_port, A2 => n41, ZN => 
                           sub_126_G9_carry_15_port);
   U351 : XOR2_X1 port map( A => n40, B => sub_126_G9_carry_14_port, Z => 
                           A_neg_8_14_port);
   U352 : AND2_X1 port map( A1 => sub_126_G9_carry_13_port, A2 => n38, ZN => 
                           sub_126_G9_carry_14_port);
   U353 : XOR2_X1 port map( A => n37, B => sub_126_G9_carry_13_port, Z => 
                           A_neg_8_13_port);
   U354 : AND2_X1 port map( A1 => sub_126_G9_carry_12_port, A2 => n35, ZN => 
                           sub_126_G9_carry_13_port);
   U355 : XOR2_X1 port map( A => n34, B => sub_126_G9_carry_12_port, Z => 
                           A_neg_8_12_port);
   U356 : AND2_X1 port map( A1 => sub_126_G9_carry_11_port, A2 => n32, ZN => 
                           sub_126_G9_carry_12_port);
   U357 : XOR2_X1 port map( A => n31, B => sub_126_G9_carry_11_port, Z => 
                           A_neg_8_11_port);
   U358 : AND2_X1 port map( A1 => sub_126_G9_carry_10_port, A2 => n29, ZN => 
                           sub_126_G9_carry_11_port);
   U359 : XOR2_X1 port map( A => n28, B => sub_126_G9_carry_10_port, Z => 
                           A_neg_8_10_port);
   U360 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G9_carry_10_port);
   U361 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_8_9_port);
   U362 : XOR2_X1 port map( A => n67, B => sub_126_G12_carry_26_port, Z => 
                           A_neg_11_26_port);
   U363 : AND2_X1 port map( A1 => sub_126_G12_carry_25_port, A2 => n65, ZN => 
                           sub_126_G12_carry_26_port);
   U364 : XOR2_X1 port map( A => n64, B => sub_126_G12_carry_25_port, Z => 
                           A_neg_11_25_port);
   U365 : AND2_X1 port map( A1 => sub_126_G12_carry_24_port, A2 => n62, ZN => 
                           sub_126_G12_carry_25_port);
   U366 : XOR2_X1 port map( A => n61, B => sub_126_G12_carry_24_port, Z => 
                           A_neg_11_24_port);
   U367 : AND2_X1 port map( A1 => sub_126_G12_carry_23_port, A2 => n59, ZN => 
                           sub_126_G12_carry_24_port);
   U368 : XOR2_X1 port map( A => n58, B => sub_126_G12_carry_23_port, Z => 
                           A_neg_11_23_port);
   U369 : AND2_X1 port map( A1 => sub_126_G12_carry_22_port, A2 => n56, ZN => 
                           sub_126_G12_carry_23_port);
   U370 : XOR2_X1 port map( A => n55, B => sub_126_G12_carry_22_port, Z => 
                           A_neg_11_22_port);
   U371 : AND2_X1 port map( A1 => sub_126_G12_carry_21_port, A2 => n53, ZN => 
                           sub_126_G12_carry_22_port);
   U372 : XOR2_X1 port map( A => n52, B => sub_126_G12_carry_21_port, Z => 
                           A_neg_11_21_port);
   U373 : AND2_X1 port map( A1 => sub_126_G12_carry_20_port, A2 => n50, ZN => 
                           sub_126_G12_carry_21_port);
   U374 : XOR2_X1 port map( A => n49, B => sub_126_G12_carry_20_port, Z => 
                           A_neg_11_20_port);
   U375 : AND2_X1 port map( A1 => sub_126_G12_carry_19_port, A2 => n47, ZN => 
                           sub_126_G12_carry_20_port);
   U376 : XOR2_X1 port map( A => n46, B => sub_126_G12_carry_19_port, Z => 
                           A_neg_11_19_port);
   U377 : AND2_X1 port map( A1 => sub_126_G12_carry_18_port, A2 => n44, ZN => 
                           sub_126_G12_carry_19_port);
   U378 : XOR2_X1 port map( A => n43, B => sub_126_G12_carry_18_port, Z => 
                           A_neg_11_18_port);
   U379 : AND2_X1 port map( A1 => sub_126_G12_carry_17_port, A2 => n41, ZN => 
                           sub_126_G12_carry_18_port);
   U380 : XOR2_X1 port map( A => n40, B => sub_126_G12_carry_17_port, Z => 
                           A_neg_11_17_port);
   U381 : AND2_X1 port map( A1 => sub_126_G12_carry_16_port, A2 => n38, ZN => 
                           sub_126_G12_carry_17_port);
   U382 : XOR2_X1 port map( A => n37, B => sub_126_G12_carry_16_port, Z => 
                           A_neg_11_16_port);
   U383 : AND2_X1 port map( A1 => sub_126_G12_carry_15_port, A2 => n35, ZN => 
                           sub_126_G12_carry_16_port);
   U384 : XOR2_X1 port map( A => n34, B => sub_126_G12_carry_15_port, Z => 
                           A_neg_11_15_port);
   U385 : AND2_X1 port map( A1 => sub_126_G12_carry_14_port, A2 => n32, ZN => 
                           sub_126_G12_carry_15_port);
   U386 : XOR2_X1 port map( A => n31, B => sub_126_G12_carry_14_port, Z => 
                           A_neg_11_14_port);
   U387 : AND2_X1 port map( A1 => sub_126_G12_carry_13_port, A2 => n29, ZN => 
                           sub_126_G12_carry_14_port);
   U388 : XOR2_X1 port map( A => n28, B => sub_126_G12_carry_13_port, Z => 
                           A_neg_11_13_port);
   U389 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G12_carry_13_port);
   U390 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_11_12_port);
   U391 : XOR2_X1 port map( A => n67, B => sub_126_G11_carry_25_port, Z => 
                           A_neg_10_25_port);
   U392 : AND2_X1 port map( A1 => sub_126_G11_carry_24_port, A2 => n65, ZN => 
                           sub_126_G11_carry_25_port);
   U393 : XOR2_X1 port map( A => n64, B => sub_126_G11_carry_24_port, Z => 
                           A_neg_10_24_port);
   U394 : AND2_X1 port map( A1 => sub_126_G11_carry_23_port, A2 => n62, ZN => 
                           sub_126_G11_carry_24_port);
   U395 : XOR2_X1 port map( A => n61, B => sub_126_G11_carry_23_port, Z => 
                           A_neg_10_23_port);
   U396 : AND2_X1 port map( A1 => sub_126_G11_carry_22_port, A2 => n59, ZN => 
                           sub_126_G11_carry_23_port);
   U397 : XOR2_X1 port map( A => n58, B => sub_126_G11_carry_22_port, Z => 
                           A_neg_10_22_port);
   U398 : AND2_X1 port map( A1 => sub_126_G11_carry_21_port, A2 => n56, ZN => 
                           sub_126_G11_carry_22_port);
   U399 : XOR2_X1 port map( A => n55, B => sub_126_G11_carry_21_port, Z => 
                           A_neg_10_21_port);
   U400 : AND2_X1 port map( A1 => sub_126_G11_carry_20_port, A2 => n53, ZN => 
                           sub_126_G11_carry_21_port);
   U401 : XOR2_X1 port map( A => n52, B => sub_126_G11_carry_20_port, Z => 
                           A_neg_10_20_port);
   U402 : AND2_X1 port map( A1 => sub_126_G11_carry_19_port, A2 => n50, ZN => 
                           sub_126_G11_carry_20_port);
   U403 : XOR2_X1 port map( A => n49, B => sub_126_G11_carry_19_port, Z => 
                           A_neg_10_19_port);
   U404 : AND2_X1 port map( A1 => sub_126_G11_carry_18_port, A2 => n47, ZN => 
                           sub_126_G11_carry_19_port);
   U405 : XOR2_X1 port map( A => n46, B => sub_126_G11_carry_18_port, Z => 
                           A_neg_10_18_port);
   U406 : AND2_X1 port map( A1 => sub_126_G11_carry_17_port, A2 => n44, ZN => 
                           sub_126_G11_carry_18_port);
   U407 : XOR2_X1 port map( A => n43, B => sub_126_G11_carry_17_port, Z => 
                           A_neg_10_17_port);
   U408 : AND2_X1 port map( A1 => sub_126_G11_carry_16_port, A2 => n41, ZN => 
                           sub_126_G11_carry_17_port);
   U409 : XOR2_X1 port map( A => n40, B => sub_126_G11_carry_16_port, Z => 
                           A_neg_10_16_port);
   U410 : AND2_X1 port map( A1 => sub_126_G11_carry_15_port, A2 => n38, ZN => 
                           sub_126_G11_carry_16_port);
   U411 : XOR2_X1 port map( A => n37, B => sub_126_G11_carry_15_port, Z => 
                           A_neg_10_15_port);
   U412 : AND2_X1 port map( A1 => sub_126_G11_carry_14_port, A2 => n35, ZN => 
                           sub_126_G11_carry_15_port);
   U413 : XOR2_X1 port map( A => n34, B => sub_126_G11_carry_14_port, Z => 
                           A_neg_10_14_port);
   U414 : AND2_X1 port map( A1 => sub_126_G11_carry_13_port, A2 => n32, ZN => 
                           sub_126_G11_carry_14_port);
   U415 : XOR2_X1 port map( A => n31, B => sub_126_G11_carry_13_port, Z => 
                           A_neg_10_13_port);
   U416 : AND2_X1 port map( A1 => sub_126_G11_carry_12_port, A2 => n29, ZN => 
                           sub_126_G11_carry_13_port);
   U417 : XOR2_X1 port map( A => n28, B => sub_126_G11_carry_12_port, Z => 
                           A_neg_10_12_port);
   U418 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G11_carry_12_port);
   U419 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_10_11_port);
   U420 : XOR2_X1 port map( A => n67, B => sub_126_G14_carry_28_port, Z => 
                           A_neg_13_28_port);
   U421 : AND2_X1 port map( A1 => sub_126_G14_carry_27_port, A2 => n65, ZN => 
                           sub_126_G14_carry_28_port);
   U422 : XOR2_X1 port map( A => n64, B => sub_126_G14_carry_27_port, Z => 
                           A_neg_13_27_port);
   U423 : AND2_X1 port map( A1 => sub_126_G14_carry_26_port, A2 => n62, ZN => 
                           sub_126_G14_carry_27_port);
   U424 : XOR2_X1 port map( A => n61, B => sub_126_G14_carry_26_port, Z => 
                           A_neg_13_26_port);
   U425 : AND2_X1 port map( A1 => sub_126_G14_carry_25_port, A2 => n59, ZN => 
                           sub_126_G14_carry_26_port);
   U426 : XOR2_X1 port map( A => n58, B => sub_126_G14_carry_25_port, Z => 
                           A_neg_13_25_port);
   U427 : AND2_X1 port map( A1 => sub_126_G14_carry_24_port, A2 => n56, ZN => 
                           sub_126_G14_carry_25_port);
   U428 : XOR2_X1 port map( A => n55, B => sub_126_G14_carry_24_port, Z => 
                           A_neg_13_24_port);
   U429 : AND2_X1 port map( A1 => sub_126_G14_carry_23_port, A2 => n53, ZN => 
                           sub_126_G14_carry_24_port);
   U430 : XOR2_X1 port map( A => n52, B => sub_126_G14_carry_23_port, Z => 
                           A_neg_13_23_port);
   U431 : AND2_X1 port map( A1 => sub_126_G14_carry_22_port, A2 => n50, ZN => 
                           sub_126_G14_carry_23_port);
   U432 : XOR2_X1 port map( A => n49, B => sub_126_G14_carry_22_port, Z => 
                           A_neg_13_22_port);
   U433 : AND2_X1 port map( A1 => sub_126_G14_carry_21_port, A2 => n47, ZN => 
                           sub_126_G14_carry_22_port);
   U434 : XOR2_X1 port map( A => n46, B => sub_126_G14_carry_21_port, Z => 
                           A_neg_13_21_port);
   U435 : AND2_X1 port map( A1 => sub_126_G14_carry_20_port, A2 => n44, ZN => 
                           sub_126_G14_carry_21_port);
   U436 : XOR2_X1 port map( A => n43, B => sub_126_G14_carry_20_port, Z => 
                           A_neg_13_20_port);
   U437 : AND2_X1 port map( A1 => sub_126_G14_carry_19_port, A2 => n41, ZN => 
                           sub_126_G14_carry_20_port);
   U438 : XOR2_X1 port map( A => n40, B => sub_126_G14_carry_19_port, Z => 
                           A_neg_13_19_port);
   U439 : AND2_X1 port map( A1 => sub_126_G14_carry_18_port, A2 => n38, ZN => 
                           sub_126_G14_carry_19_port);
   U440 : XOR2_X1 port map( A => n37, B => sub_126_G14_carry_18_port, Z => 
                           A_neg_13_18_port);
   U441 : AND2_X1 port map( A1 => sub_126_G14_carry_17_port, A2 => n35, ZN => 
                           sub_126_G14_carry_18_port);
   U442 : XOR2_X1 port map( A => n34, B => sub_126_G14_carry_17_port, Z => 
                           A_neg_13_17_port);
   U443 : AND2_X1 port map( A1 => sub_126_G14_carry_16_port, A2 => n32, ZN => 
                           sub_126_G14_carry_17_port);
   U444 : XOR2_X1 port map( A => n31, B => sub_126_G14_carry_16_port, Z => 
                           A_neg_13_16_port);
   U445 : AND2_X1 port map( A1 => sub_126_G14_carry_15_port, A2 => n29, ZN => 
                           sub_126_G14_carry_16_port);
   U446 : XOR2_X1 port map( A => n28, B => sub_126_G14_carry_15_port, Z => 
                           A_neg_13_15_port);
   U447 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G14_carry_15_port);
   U448 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_13_14_port);
   U449 : XOR2_X1 port map( A => n67, B => sub_126_G13_carry_27_port, Z => 
                           A_neg_12_27_port);
   U450 : AND2_X1 port map( A1 => sub_126_G13_carry_26_port, A2 => n65, ZN => 
                           sub_126_G13_carry_27_port);
   U451 : XOR2_X1 port map( A => n64, B => sub_126_G13_carry_26_port, Z => 
                           A_neg_12_26_port);
   U452 : AND2_X1 port map( A1 => sub_126_G13_carry_25_port, A2 => n62, ZN => 
                           sub_126_G13_carry_26_port);
   U453 : XOR2_X1 port map( A => n61, B => sub_126_G13_carry_25_port, Z => 
                           A_neg_12_25_port);
   U454 : AND2_X1 port map( A1 => sub_126_G13_carry_24_port, A2 => n59, ZN => 
                           sub_126_G13_carry_25_port);
   U455 : XOR2_X1 port map( A => n58, B => sub_126_G13_carry_24_port, Z => 
                           A_neg_12_24_port);
   U456 : AND2_X1 port map( A1 => sub_126_G13_carry_23_port, A2 => n56, ZN => 
                           sub_126_G13_carry_24_port);
   U457 : XOR2_X1 port map( A => n55, B => sub_126_G13_carry_23_port, Z => 
                           A_neg_12_23_port);
   U458 : AND2_X1 port map( A1 => sub_126_G13_carry_22_port, A2 => n53, ZN => 
                           sub_126_G13_carry_23_port);
   U459 : XOR2_X1 port map( A => n52, B => sub_126_G13_carry_22_port, Z => 
                           A_neg_12_22_port);
   U460 : AND2_X1 port map( A1 => sub_126_G13_carry_21_port, A2 => n50, ZN => 
                           sub_126_G13_carry_22_port);
   U461 : XOR2_X1 port map( A => n49, B => sub_126_G13_carry_21_port, Z => 
                           A_neg_12_21_port);
   U462 : AND2_X1 port map( A1 => sub_126_G13_carry_20_port, A2 => n47, ZN => 
                           sub_126_G13_carry_21_port);
   U463 : XOR2_X1 port map( A => n46, B => sub_126_G13_carry_20_port, Z => 
                           A_neg_12_20_port);
   U464 : AND2_X1 port map( A1 => sub_126_G13_carry_19_port, A2 => n44, ZN => 
                           sub_126_G13_carry_20_port);
   U465 : XOR2_X1 port map( A => n43, B => sub_126_G13_carry_19_port, Z => 
                           A_neg_12_19_port);
   U466 : AND2_X1 port map( A1 => sub_126_G13_carry_18_port, A2 => n41, ZN => 
                           sub_126_G13_carry_19_port);
   U467 : XOR2_X1 port map( A => n40, B => sub_126_G13_carry_18_port, Z => 
                           A_neg_12_18_port);
   U468 : AND2_X1 port map( A1 => sub_126_G13_carry_17_port, A2 => n38, ZN => 
                           sub_126_G13_carry_18_port);
   U469 : XOR2_X1 port map( A => n37, B => sub_126_G13_carry_17_port, Z => 
                           A_neg_12_17_port);
   U470 : AND2_X1 port map( A1 => sub_126_G13_carry_16_port, A2 => n35, ZN => 
                           sub_126_G13_carry_17_port);
   U471 : XOR2_X1 port map( A => n34, B => sub_126_G13_carry_16_port, Z => 
                           A_neg_12_16_port);
   U472 : AND2_X1 port map( A1 => sub_126_G13_carry_15_port, A2 => n32, ZN => 
                           sub_126_G13_carry_16_port);
   U473 : XOR2_X1 port map( A => n31, B => sub_126_G13_carry_15_port, Z => 
                           A_neg_12_15_port);
   U474 : AND2_X1 port map( A1 => sub_126_G13_carry_14_port, A2 => n29, ZN => 
                           sub_126_G13_carry_15_port);
   U475 : XOR2_X1 port map( A => n28, B => sub_126_G13_carry_14_port, Z => 
                           A_neg_12_14_port);
   U476 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G13_carry_14_port);
   U477 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_12_13_port);
   U478 : XOR2_X1 port map( A => n67, B => sub_126_G16_carry_30_port, Z => 
                           A_neg_15_30_port);
   U479 : AND2_X1 port map( A1 => sub_126_G16_carry_29_port, A2 => n64, ZN => 
                           sub_126_G16_carry_30_port);
   U480 : XOR2_X1 port map( A => n64, B => sub_126_G16_carry_29_port, Z => 
                           A_neg_15_29_port);
   U481 : AND2_X1 port map( A1 => sub_126_G16_carry_28_port, A2 => n61, ZN => 
                           sub_126_G16_carry_29_port);
   U482 : XOR2_X1 port map( A => n61, B => sub_126_G16_carry_28_port, Z => 
                           A_neg_15_28_port);
   U483 : AND2_X1 port map( A1 => sub_126_G16_carry_27_port, A2 => n58, ZN => 
                           sub_126_G16_carry_28_port);
   U484 : XOR2_X1 port map( A => n58, B => sub_126_G16_carry_27_port, Z => 
                           A_neg_15_27_port);
   U485 : AND2_X1 port map( A1 => sub_126_G16_carry_26_port, A2 => n55, ZN => 
                           sub_126_G16_carry_27_port);
   U486 : XOR2_X1 port map( A => n55, B => sub_126_G16_carry_26_port, Z => 
                           A_neg_15_26_port);
   U487 : AND2_X1 port map( A1 => sub_126_G16_carry_25_port, A2 => n52, ZN => 
                           sub_126_G16_carry_26_port);
   U488 : XOR2_X1 port map( A => n52, B => sub_126_G16_carry_25_port, Z => 
                           A_neg_15_25_port);
   U489 : AND2_X1 port map( A1 => sub_126_G16_carry_24_port, A2 => n49, ZN => 
                           sub_126_G16_carry_25_port);
   U490 : XOR2_X1 port map( A => n49, B => sub_126_G16_carry_24_port, Z => 
                           A_neg_15_24_port);
   U491 : AND2_X1 port map( A1 => sub_126_G16_carry_23_port, A2 => n46, ZN => 
                           sub_126_G16_carry_24_port);
   U492 : XOR2_X1 port map( A => n46, B => sub_126_G16_carry_23_port, Z => 
                           A_neg_15_23_port);
   U493 : AND2_X1 port map( A1 => sub_126_G16_carry_22_port, A2 => n43, ZN => 
                           sub_126_G16_carry_23_port);
   U494 : XOR2_X1 port map( A => n43, B => sub_126_G16_carry_22_port, Z => 
                           A_neg_15_22_port);
   U495 : AND2_X1 port map( A1 => sub_126_G16_carry_21_port, A2 => n40, ZN => 
                           sub_126_G16_carry_22_port);
   U496 : XOR2_X1 port map( A => n40, B => sub_126_G16_carry_21_port, Z => 
                           A_neg_15_21_port);
   U497 : AND2_X1 port map( A1 => sub_126_G16_carry_20_port, A2 => n37, ZN => 
                           sub_126_G16_carry_21_port);
   U498 : XOR2_X1 port map( A => n37, B => sub_126_G16_carry_20_port, Z => 
                           A_neg_15_20_port);
   U499 : AND2_X1 port map( A1 => sub_126_G16_carry_19_port, A2 => n34, ZN => 
                           sub_126_G16_carry_20_port);
   U500 : XOR2_X1 port map( A => n34, B => sub_126_G16_carry_19_port, Z => 
                           A_neg_15_19_port);
   U501 : AND2_X1 port map( A1 => sub_126_G16_carry_18_port, A2 => n31, ZN => 
                           sub_126_G16_carry_19_port);
   U502 : XOR2_X1 port map( A => n31, B => sub_126_G16_carry_18_port, Z => 
                           A_neg_15_18_port);
   U503 : AND2_X1 port map( A1 => sub_126_G16_carry_17_port, A2 => n28, ZN => 
                           sub_126_G16_carry_18_port);
   U504 : XOR2_X1 port map( A => n28, B => sub_126_G16_carry_17_port, Z => 
                           A_neg_15_17_port);
   U505 : AND2_X1 port map( A1 => n19, A2 => n25, ZN => 
                           sub_126_G16_carry_17_port);
   U506 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_15_16_port);
   U507 : XOR2_X1 port map( A => n67, B => sub_126_G15_carry_29_port, Z => 
                           A_neg_14_29_port);
   U508 : AND2_X1 port map( A1 => sub_126_G15_carry_28_port, A2 => n65, ZN => 
                           sub_126_G15_carry_29_port);
   U509 : XOR2_X1 port map( A => n64, B => sub_126_G15_carry_28_port, Z => 
                           A_neg_14_28_port);
   U510 : AND2_X1 port map( A1 => sub_126_G15_carry_27_port, A2 => n62, ZN => 
                           sub_126_G15_carry_28_port);
   U511 : XOR2_X1 port map( A => n61, B => sub_126_G15_carry_27_port, Z => 
                           A_neg_14_27_port);
   U512 : AND2_X1 port map( A1 => sub_126_G15_carry_26_port, A2 => n59, ZN => 
                           sub_126_G15_carry_27_port);
   U513 : XOR2_X1 port map( A => n58, B => sub_126_G15_carry_26_port, Z => 
                           A_neg_14_26_port);
   U514 : AND2_X1 port map( A1 => sub_126_G15_carry_25_port, A2 => n56, ZN => 
                           sub_126_G15_carry_26_port);
   U515 : XOR2_X1 port map( A => n55, B => sub_126_G15_carry_25_port, Z => 
                           A_neg_14_25_port);
   U516 : AND2_X1 port map( A1 => sub_126_G15_carry_24_port, A2 => n53, ZN => 
                           sub_126_G15_carry_25_port);
   U517 : XOR2_X1 port map( A => n52, B => sub_126_G15_carry_24_port, Z => 
                           A_neg_14_24_port);
   U518 : AND2_X1 port map( A1 => sub_126_G15_carry_23_port, A2 => n50, ZN => 
                           sub_126_G15_carry_24_port);
   U519 : XOR2_X1 port map( A => n49, B => sub_126_G15_carry_23_port, Z => 
                           A_neg_14_23_port);
   U520 : AND2_X1 port map( A1 => sub_126_G15_carry_22_port, A2 => n47, ZN => 
                           sub_126_G15_carry_23_port);
   U521 : XOR2_X1 port map( A => n46, B => sub_126_G15_carry_22_port, Z => 
                           A_neg_14_22_port);
   U522 : AND2_X1 port map( A1 => sub_126_G15_carry_21_port, A2 => n44, ZN => 
                           sub_126_G15_carry_22_port);
   U523 : XOR2_X1 port map( A => n43, B => sub_126_G15_carry_21_port, Z => 
                           A_neg_14_21_port);
   U524 : AND2_X1 port map( A1 => sub_126_G15_carry_20_port, A2 => n41, ZN => 
                           sub_126_G15_carry_21_port);
   U525 : XOR2_X1 port map( A => n40, B => sub_126_G15_carry_20_port, Z => 
                           A_neg_14_20_port);
   U526 : AND2_X1 port map( A1 => sub_126_G15_carry_19_port, A2 => n38, ZN => 
                           sub_126_G15_carry_20_port);
   U527 : XOR2_X1 port map( A => n37, B => sub_126_G15_carry_19_port, Z => 
                           A_neg_14_19_port);
   U528 : AND2_X1 port map( A1 => sub_126_G15_carry_18_port, A2 => n35, ZN => 
                           sub_126_G15_carry_19_port);
   U529 : XOR2_X1 port map( A => n34, B => sub_126_G15_carry_18_port, Z => 
                           A_neg_14_18_port);
   U530 : AND2_X1 port map( A1 => sub_126_G15_carry_17_port, A2 => n32, ZN => 
                           sub_126_G15_carry_18_port);
   U531 : XOR2_X1 port map( A => n31, B => sub_126_G15_carry_17_port, Z => 
                           A_neg_14_17_port);
   U532 : AND2_X1 port map( A1 => sub_126_G15_carry_16_port, A2 => n29, ZN => 
                           sub_126_G15_carry_17_port);
   U533 : XOR2_X1 port map( A => n28, B => sub_126_G15_carry_16_port, Z => 
                           A_neg_14_16_port);
   U534 : AND2_X1 port map( A1 => n19, A2 => n26, ZN => 
                           sub_126_G15_carry_16_port);
   U535 : XOR2_X1 port map( A => n25, B => n18, Z => A_neg_14_15_port);
   n70 <= '0';

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CMP_NBIT32 is

   port( SUM : in std_logic_vector (31 downto 0);  Cout : in std_logic;  A_L_B,
         A_LE_B, A_G_B, A_GE_B, A_E_B, A_NE_B : out std_logic);

end CMP_NBIT32;

architecture SYN_structural of CMP_NBIT32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N29, A_E_B_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13 :
      std_logic;

begin
   A_E_B <= A_E_B_port;
   A_NE_B <= N29;
   
   U1 : NOR3_X1 port map( A1 => n8, A2 => SUM(29), A3 => SUM(27), ZN => n10);
   U2 : OR4_X1 port map( A1 => SUM(17), A2 => SUM(15), A3 => n7, A4 => SUM(21),
                           ZN => n8);
   U3 : OR3_X1 port map( A1 => SUM(13), A2 => n6, A3 => SUM(19), ZN => n7);
   U4 : AND4_X1 port map( A1 => n12, A2 => n11, A3 => n10, A4 => n9, ZN => 
                           A_E_B_port);
   U5 : OR3_X1 port map( A1 => SUM(5), A2 => SUM(6), A3 => n2, ZN => n3);
   U6 : OR4_X1 port map( A1 => SUM(4), A2 => SUM(0), A3 => SUM(1), A4 => SUM(2)
                           , ZN => n2);
   U7 : NOR4_X1 port map( A1 => SUM(24), A2 => SUM(22), A3 => SUM(20), A4 => n5
                           , ZN => n12);
   U8 : OR4_X1 port map( A1 => SUM(16), A2 => SUM(14), A3 => SUM(18), A4 => n4,
                           ZN => n5);
   U9 : OR4_X1 port map( A1 => SUM(10), A2 => SUM(8), A3 => n3, A4 => SUM(12), 
                           ZN => n4);
   U10 : NOR3_X1 port map( A1 => SUM(26), A2 => SUM(28), A3 => SUM(30), ZN => 
                           n11);
   U11 : OR4_X1 port map( A1 => SUM(11), A2 => SUM(7), A3 => SUM(3), A4 => 
                           SUM(9), ZN => n6);
   U12 : NOR2_X1 port map( A1 => SUM(25), A2 => SUM(23), ZN => n9);
   U13 : NAND4_X1 port map( A1 => n12, A2 => n11, A3 => n10, A4 => n9, ZN => 
                           N29);
   U14 : INV_X1 port map( A => Cout, ZN => n13);
   U15 : NAND2_X1 port map( A1 => n13, A2 => N29, ZN => A_GE_B);
   U16 : NOR2_X1 port map( A1 => A_E_B_port, A2 => n13, ZN => A_G_B);
   U17 : NAND2_X1 port map( A1 => Cout, A2 => N29, ZN => A_LE_B);
   U18 : NOR2_X1 port map( A1 => Cout, A2 => A_E_B_port, ZN => A_L_B);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LOGIC_NBIT32_N_SELECTOR4 is

   port( S : in std_logic_vector (3 downto 0);  A, B : in std_logic_vector (31 
         downto 0);  O : out std_logic_vector (31 downto 0));

end LOGIC_NBIT32_N_SELECTOR4;

architecture SYN_structural of LOGIC_NBIT32_N_SELECTOR4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4_1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_2
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_3
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_4
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_2
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_5
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_6
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_7
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_8
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_3
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_9
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_10
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_11
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_12
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_4
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_13
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_14
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_15
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_16
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_5
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_17
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_18
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_19
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_20
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_6
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_21
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_22
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_23
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_24
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_7
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_25
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_26
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_27
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_28
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_8
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_29
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_30
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_31
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_32
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_9
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_33
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_34
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_35
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_36
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_10
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_37
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_38
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_39
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_40
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_11
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_41
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_42
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_43
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_44
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_12
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_45
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_46
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_47
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_48
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_13
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_49
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_50
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_51
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_52
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_14
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_53
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_54
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_55
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_56
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_15
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_57
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_58
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_59
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_60
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_16
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_61
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_62
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_63
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_64
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_17
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_65
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_66
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_67
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_68
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_18
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_69
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_70
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_71
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_72
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_19
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_73
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_74
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_75
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_76
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_20
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_77
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_78
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_79
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_80
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_21
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_81
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_82
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_83
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_84
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_22
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_85
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_86
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_87
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_88
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_23
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_89
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_90
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_91
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_92
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_24
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_93
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_94
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_95
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_96
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_25
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_97
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_98
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_99
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_100
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_26
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_101
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_102
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_103
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_104
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_27
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_105
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_106
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_107
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_108
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_28
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_109
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_110
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_111
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_112
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_29
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_113
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_114
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_115
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_116
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_30
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_117
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_118
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_119
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_120
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_31
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_121
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_122
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_123
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_124
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_0
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_125
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_126
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_127
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_0
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal An_31_port, An_30_port, An_29_port, An_28_port, An_27_port, 
      An_26_port, An_25_port, An_24_port, An_23_port, An_22_port, An_21_port, 
      An_20_port, An_19_port, An_18_port, An_17_port, An_16_port, An_15_port, 
      An_14_port, An_13_port, An_12_port, An_11_port, An_10_port, An_9_port, 
      An_8_port, An_7_port, An_6_port, An_5_port, An_4_port, An_3_port, 
      An_2_port, An_1_port, An_0_port, Bn_31_port, Bn_30_port, Bn_29_port, 
      Bn_28_port, Bn_27_port, Bn_26_port, Bn_25_port, Bn_24_port, Bn_23_port, 
      Bn_22_port, Bn_21_port, Bn_20_port, Bn_19_port, Bn_18_port, Bn_17_port, 
      Bn_16_port, Bn_15_port, Bn_14_port, Bn_13_port, Bn_12_port, Bn_11_port, 
      Bn_10_port, Bn_9_port, Bn_8_port, Bn_7_port, Bn_6_port, Bn_5_port, 
      Bn_4_port, Bn_3_port, Bn_2_port, Bn_1_port, Bn_0_port, l0_31_port, 
      l0_30_port, l0_29_port, l0_28_port, l0_27_port, l0_26_port, l0_25_port, 
      l0_24_port, l0_23_port, l0_22_port, l0_21_port, l0_20_port, l0_19_port, 
      l0_18_port, l0_17_port, l0_16_port, l0_15_port, l0_14_port, l0_13_port, 
      l0_12_port, l0_11_port, l0_10_port, l0_9_port, l0_8_port, l0_7_port, 
      l0_6_port, l0_5_port, l0_4_port, l0_3_port, l0_2_port, l0_1_port, 
      l0_0_port, l1_31_port, l1_30_port, l1_29_port, l1_28_port, l1_27_port, 
      l1_26_port, l1_25_port, l1_24_port, l1_23_port, l1_22_port, l1_21_port, 
      l1_20_port, l1_19_port, l1_18_port, l1_17_port, l1_16_port, l1_15_port, 
      l1_14_port, l1_13_port, l1_12_port, l1_11_port, l1_10_port, l1_9_port, 
      l1_8_port, l1_7_port, l1_6_port, l1_5_port, l1_4_port, l1_3_port, 
      l1_2_port, l1_1_port, l1_0_port, l2_31_port, l2_30_port, l2_29_port, 
      l2_28_port, l2_27_port, l2_26_port, l2_25_port, l2_24_port, l2_23_port, 
      l2_22_port, l2_21_port, l2_20_port, l2_19_port, l2_18_port, l2_17_port, 
      l2_16_port, l2_15_port, l2_14_port, l2_13_port, l2_12_port, l2_11_port, 
      l2_10_port, l2_9_port, l2_8_port, l2_7_port, l2_6_port, l2_5_port, 
      l2_4_port, l2_3_port, l2_2_port, l2_1_port, l2_0_port, l3_31_port, 
      l3_30_port, l3_29_port, l3_28_port, l3_27_port, l3_26_port, l3_25_port, 
      l3_24_port, l3_23_port, l3_22_port, l3_21_port, l3_20_port, l3_19_port, 
      l3_18_port, l3_17_port, l3_16_port, l3_15_port, l3_14_port, l3_13_port, 
      l3_12_port, l3_11_port, l3_10_port, l3_9_port, l3_8_port, l3_7_port, 
      l3_6_port, l3_5_port, l3_4_port, l3_3_port, l3_2_port, l3_1_port, 
      l3_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16 : std_logic;

begin
   
   A_i_0 : IV_0 port map( A => A(0), Y => An_0_port);
   A_i_1 : IV_63 port map( A => A(1), Y => An_1_port);
   A_i_2 : IV_62 port map( A => A(2), Y => An_2_port);
   A_i_3 : IV_61 port map( A => A(3), Y => An_3_port);
   A_i_4 : IV_60 port map( A => A(4), Y => An_4_port);
   A_i_5 : IV_59 port map( A => A(5), Y => An_5_port);
   A_i_6 : IV_58 port map( A => A(6), Y => An_6_port);
   A_i_7 : IV_57 port map( A => A(7), Y => An_7_port);
   A_i_8 : IV_56 port map( A => A(8), Y => An_8_port);
   A_i_9 : IV_55 port map( A => A(9), Y => An_9_port);
   A_i_10 : IV_54 port map( A => A(10), Y => An_10_port);
   A_i_11 : IV_53 port map( A => A(11), Y => An_11_port);
   A_i_12 : IV_52 port map( A => A(12), Y => An_12_port);
   A_i_13 : IV_51 port map( A => A(13), Y => An_13_port);
   A_i_14 : IV_50 port map( A => A(14), Y => An_14_port);
   A_i_15 : IV_49 port map( A => A(15), Y => An_15_port);
   A_i_16 : IV_48 port map( A => A(16), Y => An_16_port);
   A_i_17 : IV_47 port map( A => A(17), Y => An_17_port);
   A_i_18 : IV_46 port map( A => A(18), Y => An_18_port);
   A_i_19 : IV_45 port map( A => A(19), Y => An_19_port);
   A_i_20 : IV_44 port map( A => A(20), Y => An_20_port);
   A_i_21 : IV_43 port map( A => A(21), Y => An_21_port);
   A_i_22 : IV_42 port map( A => A(22), Y => An_22_port);
   A_i_23 : IV_41 port map( A => A(23), Y => An_23_port);
   A_i_24 : IV_40 port map( A => A(24), Y => An_24_port);
   A_i_25 : IV_39 port map( A => A(25), Y => An_25_port);
   A_i_26 : IV_38 port map( A => A(26), Y => An_26_port);
   A_i_27 : IV_37 port map( A => A(27), Y => An_27_port);
   A_i_28 : IV_36 port map( A => A(28), Y => An_28_port);
   A_i_29 : IV_35 port map( A => A(29), Y => An_29_port);
   A_i_30 : IV_34 port map( A => A(30), Y => An_30_port);
   A_i_31 : IV_33 port map( A => A(31), Y => An_31_port);
   B_i_0 : IV_32 port map( A => B(0), Y => Bn_0_port);
   B_i_1 : IV_31 port map( A => B(1), Y => Bn_1_port);
   B_i_2 : IV_30 port map( A => B(2), Y => Bn_2_port);
   B_i_3 : IV_29 port map( A => B(3), Y => Bn_3_port);
   B_i_4 : IV_28 port map( A => B(4), Y => Bn_4_port);
   B_i_5 : IV_27 port map( A => B(5), Y => Bn_5_port);
   B_i_6 : IV_26 port map( A => B(6), Y => Bn_6_port);
   B_i_7 : IV_25 port map( A => B(7), Y => Bn_7_port);
   B_i_8 : IV_24 port map( A => B(8), Y => Bn_8_port);
   B_i_9 : IV_23 port map( A => B(9), Y => Bn_9_port);
   B_i_10 : IV_22 port map( A => B(10), Y => Bn_10_port);
   B_i_11 : IV_21 port map( A => B(11), Y => Bn_11_port);
   B_i_12 : IV_20 port map( A => B(12), Y => Bn_12_port);
   B_i_13 : IV_19 port map( A => B(13), Y => Bn_13_port);
   B_i_14 : IV_18 port map( A => B(14), Y => Bn_14_port);
   B_i_15 : IV_17 port map( A => B(15), Y => Bn_15_port);
   B_i_16 : IV_16 port map( A => B(16), Y => Bn_16_port);
   B_i_17 : IV_15 port map( A => B(17), Y => Bn_17_port);
   B_i_18 : IV_14 port map( A => B(18), Y => Bn_18_port);
   B_i_19 : IV_13 port map( A => B(19), Y => Bn_19_port);
   B_i_20 : IV_12 port map( A => B(20), Y => Bn_20_port);
   B_i_21 : IV_11 port map( A => B(21), Y => Bn_21_port);
   B_i_22 : IV_10 port map( A => B(22), Y => Bn_22_port);
   B_i_23 : IV_9 port map( A => B(23), Y => Bn_23_port);
   B_i_24 : IV_8 port map( A => B(24), Y => Bn_24_port);
   B_i_25 : IV_7 port map( A => B(25), Y => Bn_25_port);
   B_i_26 : IV_6 port map( A => B(26), Y => Bn_26_port);
   B_i_27 : IV_5 port map( A => B(27), Y => Bn_27_port);
   B_i_28 : IV_4 port map( A => B(28), Y => Bn_28_port);
   B_i_29 : IV_3 port map( A => B(29), Y => Bn_29_port);
   B_i_30 : IV_2 port map( A => B(30), Y => Bn_30_port);
   B_i_31 : IV_1 port map( A => B(31), Y => Bn_31_port);
   U0_0 : ND3_0 port map( A => n3, B => An_0_port, C => Bn_0_port, Y => 
                           l0_0_port);
   U1_0 : ND3_127 port map( A => n5, B => An_0_port, C => B(0), Y => l1_0_port)
                           ;
   U2_0 : ND3_126 port map( A => n9, B => A(0), C => Bn_0_port, Y => l2_0_port)
                           ;
   U3_0 : ND3_125 port map( A => n13, B => A(0), C => B(0), Y => l3_0_port);
   U4_0 : ND4_0 port map( A => l0_0_port, B => l1_0_port, C => l2_0_port, D => 
                           l3_0_port, Y => O(0));
   U0_1 : ND3_124 port map( A => n1, B => An_1_port, C => Bn_1_port, Y => 
                           l0_1_port);
   U1_1 : ND3_123 port map( A => n5, B => An_1_port, C => B(1), Y => l1_1_port)
                           ;
   U2_1 : ND3_122 port map( A => n9, B => A(1), C => Bn_1_port, Y => l2_1_port)
                           ;
   U3_1 : ND3_121 port map( A => n13, B => A(1), C => B(1), Y => l3_1_port);
   U4_1 : ND4_31 port map( A => l0_1_port, B => l1_1_port, C => l2_1_port, D =>
                           l3_1_port, Y => O(1));
   U0_2 : ND3_120 port map( A => n1, B => An_2_port, C => Bn_2_port, Y => 
                           l0_2_port);
   U1_2 : ND3_119 port map( A => n5, B => An_2_port, C => B(2), Y => l1_2_port)
                           ;
   U2_2 : ND3_118 port map( A => n9, B => A(2), C => Bn_2_port, Y => l2_2_port)
                           ;
   U3_2 : ND3_117 port map( A => n13, B => A(2), C => B(2), Y => l3_2_port);
   U4_2 : ND4_30 port map( A => l0_2_port, B => l1_2_port, C => l2_2_port, D =>
                           l3_2_port, Y => O(2));
   U0_3 : ND3_116 port map( A => n1, B => An_3_port, C => Bn_3_port, Y => 
                           l0_3_port);
   U1_3 : ND3_115 port map( A => n5, B => An_3_port, C => B(3), Y => l1_3_port)
                           ;
   U2_3 : ND3_114 port map( A => n9, B => A(3), C => Bn_3_port, Y => l2_3_port)
                           ;
   U3_3 : ND3_113 port map( A => n13, B => A(3), C => B(3), Y => l3_3_port);
   U4_3 : ND4_29 port map( A => l0_3_port, B => l1_3_port, C => l2_3_port, D =>
                           l3_3_port, Y => O(3));
   U0_4 : ND3_112 port map( A => n1, B => An_4_port, C => Bn_4_port, Y => 
                           l0_4_port);
   U1_4 : ND3_111 port map( A => n5, B => An_4_port, C => B(4), Y => l1_4_port)
                           ;
   U2_4 : ND3_110 port map( A => n9, B => A(4), C => Bn_4_port, Y => l2_4_port)
                           ;
   U3_4 : ND3_109 port map( A => n13, B => A(4), C => B(4), Y => l3_4_port);
   U4_4 : ND4_28 port map( A => l0_4_port, B => l1_4_port, C => l2_4_port, D =>
                           l3_4_port, Y => O(4));
   U0_5 : ND3_108 port map( A => n1, B => An_5_port, C => Bn_5_port, Y => 
                           l0_5_port);
   U1_5 : ND3_107 port map( A => n5, B => An_5_port, C => B(5), Y => l1_5_port)
                           ;
   U2_5 : ND3_106 port map( A => n9, B => A(5), C => Bn_5_port, Y => l2_5_port)
                           ;
   U3_5 : ND3_105 port map( A => n13, B => A(5), C => B(5), Y => l3_5_port);
   U4_5 : ND4_27 port map( A => l0_5_port, B => l1_5_port, C => l2_5_port, D =>
                           l3_5_port, Y => O(5));
   U0_6 : ND3_104 port map( A => n1, B => An_6_port, C => Bn_6_port, Y => 
                           l0_6_port);
   U1_6 : ND3_103 port map( A => n5, B => An_6_port, C => B(6), Y => l1_6_port)
                           ;
   U2_6 : ND3_102 port map( A => n9, B => A(6), C => Bn_6_port, Y => l2_6_port)
                           ;
   U3_6 : ND3_101 port map( A => n13, B => A(6), C => B(6), Y => l3_6_port);
   U4_6 : ND4_26 port map( A => l0_6_port, B => l1_6_port, C => l2_6_port, D =>
                           l3_6_port, Y => O(6));
   U0_7 : ND3_100 port map( A => n1, B => An_7_port, C => Bn_7_port, Y => 
                           l0_7_port);
   U1_7 : ND3_99 port map( A => n5, B => An_7_port, C => B(7), Y => l1_7_port);
   U2_7 : ND3_98 port map( A => n9, B => A(7), C => Bn_7_port, Y => l2_7_port);
   U3_7 : ND3_97 port map( A => n13, B => A(7), C => B(7), Y => l3_7_port);
   U4_7 : ND4_25 port map( A => l0_7_port, B => l1_7_port, C => l2_7_port, D =>
                           l3_7_port, Y => O(7));
   U0_8 : ND3_96 port map( A => n1, B => An_8_port, C => Bn_8_port, Y => 
                           l0_8_port);
   U1_8 : ND3_95 port map( A => n5, B => An_8_port, C => B(8), Y => l1_8_port);
   U2_8 : ND3_94 port map( A => n9, B => A(8), C => Bn_8_port, Y => l2_8_port);
   U3_8 : ND3_93 port map( A => n13, B => A(8), C => B(8), Y => l3_8_port);
   U4_8 : ND4_24 port map( A => l0_8_port, B => l1_8_port, C => l2_8_port, D =>
                           l3_8_port, Y => O(8));
   U0_9 : ND3_92 port map( A => n1, B => An_9_port, C => Bn_9_port, Y => 
                           l0_9_port);
   U1_9 : ND3_91 port map( A => n5, B => An_9_port, C => B(9), Y => l1_9_port);
   U2_9 : ND3_90 port map( A => n9, B => A(9), C => Bn_9_port, Y => l2_9_port);
   U3_9 : ND3_89 port map( A => n13, B => A(9), C => B(9), Y => l3_9_port);
   U4_9 : ND4_23 port map( A => l0_9_port, B => l1_9_port, C => l2_9_port, D =>
                           l3_9_port, Y => O(9));
   U0_10 : ND3_88 port map( A => n1, B => An_10_port, C => Bn_10_port, Y => 
                           l0_10_port);
   U1_10 : ND3_87 port map( A => n5, B => An_10_port, C => B(10), Y => 
                           l1_10_port);
   U2_10 : ND3_86 port map( A => n9, B => A(10), C => Bn_10_port, Y => 
                           l2_10_port);
   U3_10 : ND3_85 port map( A => n13, B => A(10), C => B(10), Y => l3_10_port);
   U4_10 : ND4_22 port map( A => l0_10_port, B => l1_10_port, C => l2_10_port, 
                           D => l3_10_port, Y => O(10));
   U0_11 : ND3_84 port map( A => n1, B => An_11_port, C => Bn_11_port, Y => 
                           l0_11_port);
   U1_11 : ND3_83 port map( A => n5, B => An_11_port, C => B(11), Y => 
                           l1_11_port);
   U2_11 : ND3_82 port map( A => n9, B => A(11), C => Bn_11_port, Y => 
                           l2_11_port);
   U3_11 : ND3_81 port map( A => n13, B => A(11), C => B(11), Y => l3_11_port);
   U4_11 : ND4_21 port map( A => l0_11_port, B => l1_11_port, C => l2_11_port, 
                           D => l3_11_port, Y => O(11));
   U0_12 : ND3_80 port map( A => n1, B => An_12_port, C => Bn_12_port, Y => 
                           l0_12_port);
   U1_12 : ND3_79 port map( A => n6, B => An_12_port, C => B(12), Y => 
                           l1_12_port);
   U2_12 : ND3_78 port map( A => n10, B => A(12), C => Bn_12_port, Y => 
                           l2_12_port);
   U3_12 : ND3_77 port map( A => n14, B => A(12), C => B(12), Y => l3_12_port);
   U4_12 : ND4_20 port map( A => l0_12_port, B => l1_12_port, C => l2_12_port, 
                           D => l3_12_port, Y => O(12));
   U0_13 : ND3_76 port map( A => n2, B => An_13_port, C => Bn_13_port, Y => 
                           l0_13_port);
   U1_13 : ND3_75 port map( A => n6, B => An_13_port, C => B(13), Y => 
                           l1_13_port);
   U2_13 : ND3_74 port map( A => n10, B => A(13), C => Bn_13_port, Y => 
                           l2_13_port);
   U3_13 : ND3_73 port map( A => n14, B => A(13), C => B(13), Y => l3_13_port);
   U4_13 : ND4_19 port map( A => l0_13_port, B => l1_13_port, C => l2_13_port, 
                           D => l3_13_port, Y => O(13));
   U0_14 : ND3_72 port map( A => n2, B => An_14_port, C => Bn_14_port, Y => 
                           l0_14_port);
   U1_14 : ND3_71 port map( A => n6, B => An_14_port, C => B(14), Y => 
                           l1_14_port);
   U2_14 : ND3_70 port map( A => n10, B => A(14), C => Bn_14_port, Y => 
                           l2_14_port);
   U3_14 : ND3_69 port map( A => n14, B => A(14), C => B(14), Y => l3_14_port);
   U4_14 : ND4_18 port map( A => l0_14_port, B => l1_14_port, C => l2_14_port, 
                           D => l3_14_port, Y => O(14));
   U0_15 : ND3_68 port map( A => n2, B => An_15_port, C => Bn_15_port, Y => 
                           l0_15_port);
   U1_15 : ND3_67 port map( A => n6, B => An_15_port, C => B(15), Y => 
                           l1_15_port);
   U2_15 : ND3_66 port map( A => n10, B => A(15), C => Bn_15_port, Y => 
                           l2_15_port);
   U3_15 : ND3_65 port map( A => n14, B => A(15), C => B(15), Y => l3_15_port);
   U4_15 : ND4_17 port map( A => l0_15_port, B => l1_15_port, C => l2_15_port, 
                           D => l3_15_port, Y => O(15));
   U0_16 : ND3_64 port map( A => n2, B => An_16_port, C => Bn_16_port, Y => 
                           l0_16_port);
   U1_16 : ND3_63 port map( A => n6, B => An_16_port, C => B(16), Y => 
                           l1_16_port);
   U2_16 : ND3_62 port map( A => n10, B => A(16), C => Bn_16_port, Y => 
                           l2_16_port);
   U3_16 : ND3_61 port map( A => n14, B => A(16), C => B(16), Y => l3_16_port);
   U4_16 : ND4_16 port map( A => l0_16_port, B => l1_16_port, C => l2_16_port, 
                           D => l3_16_port, Y => O(16));
   U0_17 : ND3_60 port map( A => n2, B => An_17_port, C => Bn_17_port, Y => 
                           l0_17_port);
   U1_17 : ND3_59 port map( A => n6, B => An_17_port, C => B(17), Y => 
                           l1_17_port);
   U2_17 : ND3_58 port map( A => n10, B => A(17), C => Bn_17_port, Y => 
                           l2_17_port);
   U3_17 : ND3_57 port map( A => n14, B => A(17), C => B(17), Y => l3_17_port);
   U4_17 : ND4_15 port map( A => l0_17_port, B => l1_17_port, C => l2_17_port, 
                           D => l3_17_port, Y => O(17));
   U0_18 : ND3_56 port map( A => n2, B => An_18_port, C => Bn_18_port, Y => 
                           l0_18_port);
   U1_18 : ND3_55 port map( A => n6, B => An_18_port, C => B(18), Y => 
                           l1_18_port);
   U2_18 : ND3_54 port map( A => n10, B => A(18), C => Bn_18_port, Y => 
                           l2_18_port);
   U3_18 : ND3_53 port map( A => n14, B => A(18), C => B(18), Y => l3_18_port);
   U4_18 : ND4_14 port map( A => l0_18_port, B => l1_18_port, C => l2_18_port, 
                           D => l3_18_port, Y => O(18));
   U0_19 : ND3_52 port map( A => n2, B => An_19_port, C => Bn_19_port, Y => 
                           l0_19_port);
   U1_19 : ND3_51 port map( A => n6, B => An_19_port, C => B(19), Y => 
                           l1_19_port);
   U2_19 : ND3_50 port map( A => n10, B => A(19), C => Bn_19_port, Y => 
                           l2_19_port);
   U3_19 : ND3_49 port map( A => n14, B => A(19), C => B(19), Y => l3_19_port);
   U4_19 : ND4_13 port map( A => l0_19_port, B => l1_19_port, C => l2_19_port, 
                           D => l3_19_port, Y => O(19));
   U0_20 : ND3_48 port map( A => n2, B => An_20_port, C => Bn_20_port, Y => 
                           l0_20_port);
   U1_20 : ND3_47 port map( A => n6, B => An_20_port, C => B(20), Y => 
                           l1_20_port);
   U2_20 : ND3_46 port map( A => n10, B => A(20), C => Bn_20_port, Y => 
                           l2_20_port);
   U3_20 : ND3_45 port map( A => n14, B => A(20), C => B(20), Y => l3_20_port);
   U4_20 : ND4_12 port map( A => l0_20_port, B => l1_20_port, C => l2_20_port, 
                           D => l3_20_port, Y => O(20));
   U0_21 : ND3_44 port map( A => n2, B => An_21_port, C => Bn_21_port, Y => 
                           l0_21_port);
   U1_21 : ND3_43 port map( A => n6, B => An_21_port, C => B(21), Y => 
                           l1_21_port);
   U2_21 : ND3_42 port map( A => n10, B => A(21), C => Bn_21_port, Y => 
                           l2_21_port);
   U3_21 : ND3_41 port map( A => n14, B => A(21), C => B(21), Y => l3_21_port);
   U4_21 : ND4_11 port map( A => l0_21_port, B => l1_21_port, C => l2_21_port, 
                           D => l3_21_port, Y => O(21));
   U0_22 : ND3_40 port map( A => n2, B => An_22_port, C => Bn_22_port, Y => 
                           l0_22_port);
   U1_22 : ND3_39 port map( A => n6, B => An_22_port, C => B(22), Y => 
                           l1_22_port);
   U2_22 : ND3_38 port map( A => n10, B => A(22), C => Bn_22_port, Y => 
                           l2_22_port);
   U3_22 : ND3_37 port map( A => n14, B => A(22), C => B(22), Y => l3_22_port);
   U4_22 : ND4_10 port map( A => l0_22_port, B => l1_22_port, C => l2_22_port, 
                           D => l3_22_port, Y => O(22));
   U0_23 : ND3_36 port map( A => n2, B => An_23_port, C => Bn_23_port, Y => 
                           l0_23_port);
   U1_23 : ND3_35 port map( A => n6, B => An_23_port, C => B(23), Y => 
                           l1_23_port);
   U2_23 : ND3_34 port map( A => n10, B => A(23), C => Bn_23_port, Y => 
                           l2_23_port);
   U3_23 : ND3_33 port map( A => n14, B => A(23), C => B(23), Y => l3_23_port);
   U4_23 : ND4_9 port map( A => l0_23_port, B => l1_23_port, C => l2_23_port, D
                           => l3_23_port, Y => O(23));
   U0_24 : ND3_32 port map( A => n2, B => An_24_port, C => Bn_24_port, Y => 
                           l0_24_port);
   U1_24 : ND3_31 port map( A => n7, B => An_24_port, C => B(24), Y => 
                           l1_24_port);
   U2_24 : ND3_30 port map( A => n11, B => A(24), C => Bn_24_port, Y => 
                           l2_24_port);
   U3_24 : ND3_29 port map( A => n15, B => A(24), C => B(24), Y => l3_24_port);
   U4_24 : ND4_8 port map( A => l0_24_port, B => l1_24_port, C => l2_24_port, D
                           => l3_24_port, Y => O(24));
   U0_25 : ND3_28 port map( A => n3, B => An_25_port, C => Bn_25_port, Y => 
                           l0_25_port);
   U1_25 : ND3_27 port map( A => n7, B => An_25_port, C => B(25), Y => 
                           l1_25_port);
   U2_25 : ND3_26 port map( A => n11, B => A(25), C => Bn_25_port, Y => 
                           l2_25_port);
   U3_25 : ND3_25 port map( A => n15, B => A(25), C => B(25), Y => l3_25_port);
   U4_25 : ND4_7 port map( A => l0_25_port, B => l1_25_port, C => l2_25_port, D
                           => l3_25_port, Y => O(25));
   U0_26 : ND3_24 port map( A => n3, B => An_26_port, C => Bn_26_port, Y => 
                           l0_26_port);
   U1_26 : ND3_23 port map( A => n7, B => An_26_port, C => B(26), Y => 
                           l1_26_port);
   U2_26 : ND3_22 port map( A => n11, B => A(26), C => Bn_26_port, Y => 
                           l2_26_port);
   U3_26 : ND3_21 port map( A => n15, B => A(26), C => B(26), Y => l3_26_port);
   U4_26 : ND4_6 port map( A => l0_26_port, B => l1_26_port, C => l2_26_port, D
                           => l3_26_port, Y => O(26));
   U0_27 : ND3_20 port map( A => n3, B => An_27_port, C => Bn_27_port, Y => 
                           l0_27_port);
   U1_27 : ND3_19 port map( A => n7, B => An_27_port, C => B(27), Y => 
                           l1_27_port);
   U2_27 : ND3_18 port map( A => n11, B => A(27), C => Bn_27_port, Y => 
                           l2_27_port);
   U3_27 : ND3_17 port map( A => n15, B => A(27), C => B(27), Y => l3_27_port);
   U4_27 : ND4_5 port map( A => l0_27_port, B => l1_27_port, C => l2_27_port, D
                           => l3_27_port, Y => O(27));
   U0_28 : ND3_16 port map( A => n3, B => An_28_port, C => Bn_28_port, Y => 
                           l0_28_port);
   U1_28 : ND3_15 port map( A => n7, B => An_28_port, C => B(28), Y => 
                           l1_28_port);
   U2_28 : ND3_14 port map( A => n11, B => A(28), C => Bn_28_port, Y => 
                           l2_28_port);
   U3_28 : ND3_13 port map( A => n15, B => A(28), C => B(28), Y => l3_28_port);
   U4_28 : ND4_4 port map( A => l0_28_port, B => l1_28_port, C => l2_28_port, D
                           => l3_28_port, Y => O(28));
   U0_29 : ND3_12 port map( A => n3, B => An_29_port, C => Bn_29_port, Y => 
                           l0_29_port);
   U1_29 : ND3_11 port map( A => n7, B => An_29_port, C => B(29), Y => 
                           l1_29_port);
   U2_29 : ND3_10 port map( A => n11, B => A(29), C => Bn_29_port, Y => 
                           l2_29_port);
   U3_29 : ND3_9 port map( A => n15, B => A(29), C => B(29), Y => l3_29_port);
   U4_29 : ND4_3 port map( A => l0_29_port, B => l1_29_port, C => l2_29_port, D
                           => l3_29_port, Y => O(29));
   U0_30 : ND3_8 port map( A => n3, B => An_30_port, C => Bn_30_port, Y => 
                           l0_30_port);
   U1_30 : ND3_7 port map( A => n7, B => An_30_port, C => B(30), Y => 
                           l1_30_port);
   U2_30 : ND3_6 port map( A => n11, B => A(30), C => Bn_30_port, Y => 
                           l2_30_port);
   U3_30 : ND3_5 port map( A => n15, B => A(30), C => B(30), Y => l3_30_port);
   U4_30 : ND4_2 port map( A => l0_30_port, B => l1_30_port, C => l2_30_port, D
                           => l3_30_port, Y => O(30));
   U0_31 : ND3_4 port map( A => n3, B => An_31_port, C => Bn_31_port, Y => 
                           l0_31_port);
   U1_31 : ND3_3 port map( A => n7, B => An_31_port, C => B(31), Y => 
                           l1_31_port);
   U2_31 : ND3_2 port map( A => n11, B => A(31), C => Bn_31_port, Y => 
                           l2_31_port);
   U3_31 : ND3_1 port map( A => n15, B => A(31), C => B(31), Y => l3_31_port);
   U4_31 : ND4_1 port map( A => l0_31_port, B => l1_31_port, C => l2_31_port, D
                           => l3_31_port, Y => O(31));
   U1 : BUF_X1 port map( A => S(3), Z => n16);
   U2 : BUF_X1 port map( A => S(2), Z => n12);
   U3 : BUF_X1 port map( A => S(0), Z => n4);
   U4 : BUF_X1 port map( A => S(1), Z => n8);
   U5 : BUF_X1 port map( A => n16, Z => n14);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n12, Z => n9);
   U8 : BUF_X1 port map( A => n8, Z => n5);
   U9 : BUF_X1 port map( A => n4, Z => n1);
   U10 : BUF_X1 port map( A => n12, Z => n10);
   U11 : BUF_X1 port map( A => n4, Z => n2);
   U12 : BUF_X1 port map( A => n8, Z => n6);
   U13 : BUF_X1 port map( A => n16, Z => n15);
   U14 : BUF_X1 port map( A => n12, Z => n11);
   U15 : BUF_X1 port map( A => n8, Z => n7);
   U16 : BUF_X1 port map( A => n4, Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SHIFTER is

   port( data_in : in std_logic_vector (31 downto 0);  R : in std_logic_vector 
         (4 downto 0);  conf : in std_logic_vector (1 downto 0);  data_out : 
         out std_logic_vector (31 downto 0));

end SHIFTER;

architecture SYN_Behavioral of SHIFTER is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal mask_0_39_port, mask_0_38_port, mask_0_37_port, mask_0_36_port, 
      mask_0_35_port, mask_0_34_port, mask_0_33_port, mask_0_32_port, 
      mask_0_31_port, mask_0_30_port, mask_0_29_port, mask_0_28_port, 
      mask_0_27_port, mask_0_26_port, mask_0_25_port, mask_0_24_port, 
      mask_0_23_port, mask_0_22_port, mask_0_21_port, mask_0_20_port, 
      mask_0_19_port, mask_0_18_port, mask_0_17_port, mask_0_16_port, 
      mask_0_15_port, mask_0_14_port, mask_0_13_port, mask_0_12_port, 
      mask_0_11_port, mask_0_10_port, mask_0_9_port, mask_0_8_port, 
      mask_0_7_port, mask_0_6_port, mask_0_5_port, mask_0_4_port, mask_0_3_port
      , mask_0_2_port, mask_0_1_port, mask_0_0_port, mask_1_39_port, 
      mask_1_38_port, mask_1_37_port, mask_1_36_port, mask_1_35_port, 
      mask_1_34_port, mask_1_33_port, mask_1_32_port, mask_1_31_port, 
      mask_1_30_port, mask_1_29_port, mask_1_28_port, mask_1_27_port, 
      mask_1_26_port, mask_1_25_port, mask_1_24_port, mask_1_23_port, 
      mask_1_22_port, mask_1_21_port, mask_1_20_port, mask_1_19_port, 
      mask_1_18_port, mask_1_17_port, mask_1_16_port, mask_1_15_port, 
      mask_1_14_port, mask_1_13_port, mask_1_12_port, mask_1_11_port, 
      mask_1_10_port, mask_1_9_port, mask_1_8_port, mask_1_7_port, 
      mask_1_6_port, mask_1_5_port, mask_1_4_port, mask_1_3_port, mask_1_2_port
      , mask_1_1_port, mask_1_0_port, mask_2_39_port, mask_2_38_port, 
      mask_2_37_port, mask_2_36_port, mask_2_35_port, mask_2_34_port, 
      mask_2_33_port, mask_2_32_port, mask_2_31_port, mask_2_30_port, 
      mask_2_29_port, mask_2_28_port, mask_2_27_port, mask_2_26_port, 
      mask_2_25_port, mask_2_24_port, mask_2_23_port, mask_2_22_port, 
      mask_2_21_port, mask_2_20_port, mask_2_19_port, mask_2_18_port, 
      mask_2_17_port, mask_2_16_port, mask_2_15_port, mask_2_14_port, 
      mask_2_13_port, mask_2_12_port, mask_2_11_port, mask_2_10_port, 
      mask_2_9_port, mask_2_8_port, mask_2_7_port, mask_2_6_port, mask_2_5_port
      , mask_2_4_port, mask_2_3_port, mask_2_2_port, mask_2_1_port, 
      mask_2_0_port, mask_3_39_port, mask_3_38_port, mask_3_37_port, 
      mask_3_36_port, mask_3_35_port, mask_3_34_port, mask_3_33_port, 
      mask_3_32_port, mask_3_31_port, mask_3_30_port, mask_3_29_port, 
      mask_3_28_port, mask_3_27_port, mask_3_26_port, mask_3_25_port, 
      mask_3_24_port, mask_3_23_port, mask_3_22_port, mask_3_21_port, 
      mask_3_20_port, mask_3_19_port, mask_3_18_port, mask_3_17_port, 
      mask_3_16_port, mask_3_15_port, mask_3_14_port, mask_3_13_port, 
      mask_3_12_port, mask_3_11_port, mask_3_10_port, mask_3_9_port, 
      mask_3_8_port, mask_3_7_port, mask_3_6_port, mask_3_5_port, mask_3_4_port
      , mask_3_3_port, mask_3_2_port, mask_3_1_port, mask_3_0_port, N28, N35, 
      N37, N38, N39, N40, N41, N42, N43, N53, N54, N55, N56, N57, N58, N59, N60
      , N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, 
      N82, N83, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97
      , N98, N99, N108, N109, N110, N111, N112, N113, N114, N115, N116, 
      out_mask_39_port, out_mask_38_port, out_mask_37_port, out_mask_36_port, 
      out_mask_35_port, out_mask_34_port, out_mask_33_port, out_mask_32_port, 
      out_mask_5_port, out_mask_4_port, out_mask_3_port, out_mask_2_port, 
      out_mask_1_port, out_mask_0_port, N158, N159, N160, N161, N162, N163, 
      N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, 
      N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, 
      N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, 
      N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, 
      N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, n219_port, 
      n229, n238, n239, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, 
      n28_port, n29, n30, n31, n32, n33, n34, n35_port, n36, n37_port, n38_port
      , n39_port, n40_port, n41_port, n42_port, n43_port, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53_port, n54_port, n55_port, n56_port, n57_port
      , n58_port, n59_port, n60_port, n61, n62, n63, n64, n65, n66, n67, 
      n68_port, n69_port, n70_port, n71_port, n72_port, n73_port, n74_port, 
      n75_port, n76_port, n77_port, n78_port, n79_port, n80_port, n81_port, 
      n82_port, n83_port, n84, n85_port, n86_port, n87_port, n88_port, n89_port
      , n90_port, n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, 
      n97_port, n98_port, n99_port, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108_port, n109_port, n110_port, n111_port, n112_port, n113_port, 
      n114_port, n115_port, n116_port, n117, n118, n119, n120, n121, n122, n123
      , n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158_port, 
      n159_port, n160_port, n161_port, n162_port, n163_port, n164_port, 
      n165_port, n166_port, n167_port, n168_port, n169_port, n170_port, 
      n171_port, n172_port, n173_port, n174_port, n175_port, n176_port, 
      n177_port, n178_port, n179_port, n180_port, n181_port, n182_port, 
      n183_port, n184_port, n185_port, n186_port, n187_port, n188_port, 
      n189_port, n190_port, n191_port, n192_port, n193_port, n194_port, 
      n195_port, n196_port, n197_port, n198_port, n199_port, n200_port, 
      n201_port, n202_port, n203_port, n204_port, n205_port, n206_port, 
      n207_port, n208_port, n209_port, n210_port, n211_port, n212_port, 
      n213_port, n214_port, n215_port, n216_port, n217_port, n218_port, 
      n220_port, n221_port, n222, n223, n224, n225, n226, n227, n228, n230, 
      n231, n232, n233, n234, n235, n236, n237, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n598 : std_logic;

begin
   
   mask_reg_0_39_inst : DLH_X1 port map( G => n368, D => n542, Q => 
                           mask_0_39_port);
   mask_reg_0_38_inst : DLH_X1 port map( G => n368, D => n543, Q => 
                           mask_0_38_port);
   mask_reg_0_37_inst : DLH_X1 port map( G => n368, D => n544, Q => 
                           mask_0_37_port);
   mask_reg_0_36_inst : DLH_X1 port map( G => n368, D => n545, Q => 
                           mask_0_36_port);
   mask_reg_0_35_inst : DLH_X1 port map( G => n368, D => n546, Q => 
                           mask_0_35_port);
   mask_reg_0_34_inst : DLH_X1 port map( G => n368, D => n547, Q => 
                           mask_0_34_port);
   mask_reg_0_33_inst : DLH_X1 port map( G => n367, D => n548, Q => 
                           mask_0_33_port);
   mask_reg_0_32_inst : DLH_X1 port map( G => n367, D => n549, Q => 
                           mask_0_32_port);
   mask_reg_0_31_inst : DLH_X1 port map( G => n367, D => N116, Q => 
                           mask_0_31_port);
   mask_reg_0_30_inst : DLH_X1 port map( G => n367, D => N115, Q => 
                           mask_0_30_port);
   mask_reg_0_29_inst : DLH_X1 port map( G => n367, D => N114, Q => 
                           mask_0_29_port);
   mask_reg_0_28_inst : DLH_X1 port map( G => n367, D => N113, Q => 
                           mask_0_28_port);
   mask_reg_0_27_inst : DLH_X1 port map( G => n367, D => N112, Q => 
                           mask_0_27_port);
   mask_reg_0_26_inst : DLH_X1 port map( G => n367, D => N111, Q => 
                           mask_0_26_port);
   mask_reg_0_25_inst : DLH_X1 port map( G => n367, D => N110, Q => 
                           mask_0_25_port);
   mask_reg_0_24_inst : DLH_X1 port map( G => n367, D => N109, Q => 
                           mask_0_24_port);
   mask_reg_0_23_inst : DLH_X1 port map( G => n367, D => N108, Q => 
                           mask_0_23_port);
   mask_reg_0_22_inst : DLH_X1 port map( G => n366, D => n551, Q => 
                           mask_0_22_port);
   mask_reg_0_21_inst : DLH_X1 port map( G => n366, D => n552, Q => 
                           mask_0_21_port);
   mask_reg_0_20_inst : DLH_X1 port map( G => n366, D => n553, Q => 
                           mask_0_20_port);
   mask_reg_0_19_inst : DLH_X1 port map( G => n366, D => n554, Q => 
                           mask_0_19_port);
   mask_reg_0_18_inst : DLH_X1 port map( G => n366, D => n555, Q => 
                           mask_0_18_port);
   mask_reg_0_17_inst : DLH_X1 port map( G => n366, D => n556, Q => 
                           mask_0_17_port);
   mask_reg_0_16_inst : DLH_X1 port map( G => n366, D => n557, Q => 
                           mask_0_16_port);
   mask_reg_0_15_inst : DLH_X1 port map( G => n366, D => n558, Q => 
                           mask_0_15_port);
   mask_reg_0_14_inst : DLH_X1 port map( G => n366, D => N99, Q => 
                           mask_0_14_port);
   mask_reg_0_13_inst : DLH_X1 port map( G => n366, D => N98, Q => 
                           mask_0_13_port);
   mask_reg_0_12_inst : DLH_X1 port map( G => n366, D => N97, Q => 
                           mask_0_12_port);
   mask_reg_0_11_inst : DLH_X1 port map( G => n365, D => N96, Q => 
                           mask_0_11_port);
   mask_reg_0_10_inst : DLH_X1 port map( G => n365, D => N95, Q => 
                           mask_0_10_port);
   mask_reg_0_9_inst : DLH_X1 port map( G => n365, D => N94, Q => mask_0_9_port
                           );
   mask_reg_0_8_inst : DLH_X1 port map( G => n365, D => N93, Q => mask_0_8_port
                           );
   mask_reg_0_7_inst : DLH_X1 port map( G => n365, D => N92, Q => mask_0_7_port
                           );
   mask_reg_0_6_inst : DLH_X1 port map( G => n365, D => N91, Q => mask_0_6_port
                           );
   mask_reg_0_5_inst : DLH_X1 port map( G => n365, D => N90, Q => mask_0_5_port
                           );
   mask_reg_0_4_inst : DLH_X1 port map( G => n365, D => N89, Q => mask_0_4_port
                           );
   mask_reg_0_3_inst : DLH_X1 port map( G => n365, D => N88, Q => mask_0_3_port
                           );
   mask_reg_0_2_inst : DLH_X1 port map( G => n365, D => N87, Q => mask_0_2_port
                           );
   mask_reg_0_1_inst : DLH_X1 port map( G => n365, D => N86, Q => mask_0_1_port
                           );
   mask_reg_0_0_inst : DLH_X1 port map( G => n364, D => N85, Q => mask_0_0_port
                           );
   mask_reg_1_39_inst : DLH_X1 port map( G => n364, D => n550, Q => 
                           mask_1_39_port);
   mask_reg_1_38_inst : DLH_X1 port map( G => n364, D => N83, Q => 
                           mask_1_38_port);
   mask_reg_1_37_inst : DLH_X1 port map( G => n364, D => N82, Q => 
                           mask_1_37_port);
   mask_reg_1_36_inst : DLH_X1 port map( G => n364, D => N81, Q => 
                           mask_1_36_port);
   mask_reg_1_35_inst : DLH_X1 port map( G => n364, D => N80, Q => 
                           mask_1_35_port);
   mask_reg_1_34_inst : DLH_X1 port map( G => n364, D => N79, Q => 
                           mask_1_34_port);
   mask_reg_1_33_inst : DLH_X1 port map( G => n364, D => N78, Q => 
                           mask_1_33_port);
   mask_reg_1_32_inst : DLH_X1 port map( G => n364, D => N77, Q => 
                           mask_1_32_port);
   mask_reg_1_31_inst : DLH_X1 port map( G => n364, D => N60, Q => 
                           mask_1_31_port);
   mask_reg_1_30_inst : DLH_X1 port map( G => n364, D => N59, Q => 
                           mask_1_30_port);
   mask_reg_1_29_inst : DLH_X1 port map( G => n363, D => N58, Q => 
                           mask_1_29_port);
   mask_reg_1_28_inst : DLH_X1 port map( G => n363, D => N57, Q => 
                           mask_1_28_port);
   mask_reg_1_27_inst : DLH_X1 port map( G => n363, D => N56, Q => 
                           mask_1_27_port);
   mask_reg_1_26_inst : DLH_X1 port map( G => n363, D => N55, Q => 
                           mask_1_26_port);
   mask_reg_1_25_inst : DLH_X1 port map( G => n363, D => N54, Q => 
                           mask_1_25_port);
   mask_reg_1_24_inst : DLH_X1 port map( G => n363, D => N53, Q => 
                           mask_1_24_port);
   mask_reg_1_23_inst : DLH_X1 port map( G => n363, D => N76, Q => 
                           mask_1_23_port);
   mask_reg_1_22_inst : DLH_X1 port map( G => n363, D => N75, Q => 
                           mask_1_22_port);
   mask_reg_1_21_inst : DLH_X1 port map( G => n363, D => N74, Q => 
                           mask_1_21_port);
   mask_reg_1_20_inst : DLH_X1 port map( G => n363, D => N73, Q => 
                           mask_1_20_port);
   mask_reg_1_19_inst : DLH_X1 port map( G => n363, D => N72, Q => 
                           mask_1_19_port);
   mask_reg_1_18_inst : DLH_X1 port map( G => n362, D => N71, Q => 
                           mask_1_18_port);
   mask_reg_1_17_inst : DLH_X1 port map( G => n362, D => N70, Q => 
                           mask_1_17_port);
   mask_reg_1_16_inst : DLH_X1 port map( G => n362, D => N69, Q => 
                           mask_1_16_port);
   mask_reg_1_15_inst : DLH_X1 port map( G => n362, D => n533, Q => 
                           mask_1_15_port);
   mask_reg_1_14_inst : DLH_X1 port map( G => n362, D => n532, Q => 
                           mask_1_14_port);
   mask_reg_1_13_inst : DLH_X1 port map( G => n362, D => n531, Q => 
                           mask_1_13_port);
   mask_reg_1_12_inst : DLH_X1 port map( G => n362, D => n530, Q => 
                           mask_1_12_port);
   mask_reg_1_11_inst : DLH_X1 port map( G => n362, D => n529, Q => 
                           mask_1_11_port);
   mask_reg_1_10_inst : DLH_X1 port map( G => n362, D => n528, Q => 
                           mask_1_10_port);
   mask_reg_1_9_inst : DLH_X1 port map( G => n362, D => n527, Q => 
                           mask_1_9_port);
   mask_reg_1_8_inst : DLH_X1 port map( G => n362, D => n526, Q => 
                           mask_1_8_port);
   mask_reg_1_7_inst : DLH_X1 port map( G => n361, D => N68, Q => mask_1_7_port
                           );
   mask_reg_1_6_inst : DLH_X1 port map( G => n361, D => n559, Q => 
                           mask_1_6_port);
   mask_reg_1_5_inst : DLH_X1 port map( G => n361, D => n560, Q => 
                           mask_1_5_port);
   mask_reg_1_4_inst : DLH_X1 port map( G => n361, D => n561, Q => 
                           mask_1_4_port);
   mask_reg_1_3_inst : DLH_X1 port map( G => n361, D => n562, Q => 
                           mask_1_3_port);
   mask_reg_1_2_inst : DLH_X1 port map( G => n361, D => n563, Q => 
                           mask_1_2_port);
   mask_reg_1_1_inst : DLH_X1 port map( G => n361, D => n564, Q => 
                           mask_1_1_port);
   mask_reg_1_0_inst : DLH_X1 port map( G => n361, D => n565, Q => 
                           mask_1_0_port);
   mask_reg_2_39_inst : DLH_X1 port map( G => n361, D => N60, Q => 
                           mask_2_39_port);
   mask_reg_2_38_inst : DLH_X1 port map( G => n361, D => N59, Q => 
                           mask_2_38_port);
   mask_reg_2_37_inst : DLH_X1 port map( G => n361, D => N58, Q => 
                           mask_2_37_port);
   mask_reg_2_36_inst : DLH_X1 port map( G => n360, D => N57, Q => 
                           mask_2_36_port);
   mask_reg_2_35_inst : DLH_X1 port map( G => n360, D => N56, Q => 
                           mask_2_35_port);
   mask_reg_2_34_inst : DLH_X1 port map( G => n360, D => N55, Q => 
                           mask_2_34_port);
   mask_reg_2_33_inst : DLH_X1 port map( G => n360, D => N54, Q => 
                           mask_2_33_port);
   mask_reg_2_32_inst : DLH_X1 port map( G => n360, D => N53, Q => 
                           mask_2_32_port);
   mask_reg_2_31_inst : DLH_X1 port map( G => n360, D => n541, Q => 
                           mask_2_31_port);
   mask_reg_2_30_inst : DLH_X1 port map( G => n360, D => N43, Q => 
                           mask_2_30_port);
   mask_reg_2_29_inst : DLH_X1 port map( G => n360, D => N42, Q => 
                           mask_2_29_port);
   mask_reg_2_28_inst : DLH_X1 port map( G => n360, D => N41, Q => 
                           mask_2_28_port);
   mask_reg_2_27_inst : DLH_X1 port map( G => n360, D => N40, Q => 
                           mask_2_27_port);
   mask_reg_2_26_inst : DLH_X1 port map( G => n360, D => N39, Q => 
                           mask_2_26_port);
   mask_reg_2_25_inst : DLH_X1 port map( G => n359, D => N38, Q => 
                           mask_2_25_port);
   mask_reg_2_24_inst : DLH_X1 port map( G => n359, D => N37, Q => 
                           mask_2_24_port);
   mask_reg_2_23_inst : DLH_X1 port map( G => n359, D => n326, Q => 
                           mask_2_23_port);
   mask_reg_2_22_inst : DLH_X1 port map( G => n359, D => n326, Q => 
                           mask_2_22_port);
   mask_reg_2_21_inst : DLH_X1 port map( G => n359, D => n327, Q => 
                           mask_2_21_port);
   mask_reg_2_20_inst : DLH_X1 port map( G => n359, D => n327, Q => 
                           mask_2_20_port);
   mask_reg_2_19_inst : DLH_X1 port map( G => n359, D => n327, Q => 
                           mask_2_19_port);
   mask_reg_2_18_inst : DLH_X1 port map( G => n359, D => n327, Q => 
                           mask_2_18_port);
   mask_reg_2_17_inst : DLH_X1 port map( G => n359, D => n327, Q => 
                           mask_2_17_port);
   mask_reg_2_16_inst : DLH_X1 port map( G => n359, D => n328, Q => 
                           mask_2_16_port);
   mask_reg_2_15_inst : DLH_X1 port map( G => n359, D => N35, Q => 
                           mask_2_15_port);
   mask_reg_2_14_inst : DLH_X1 port map( G => n358, D => n540, Q => 
                           mask_2_14_port);
   mask_reg_2_13_inst : DLH_X1 port map( G => n358, D => n539, Q => 
                           mask_2_13_port);
   mask_reg_2_12_inst : DLH_X1 port map( G => n358, D => n538, Q => 
                           mask_2_12_port);
   mask_reg_2_11_inst : DLH_X1 port map( G => n358, D => n537, Q => 
                           mask_2_11_port);
   mask_reg_2_10_inst : DLH_X1 port map( G => n358, D => n536, Q => 
                           mask_2_10_port);
   mask_reg_2_9_inst : DLH_X1 port map( G => n358, D => n535, Q => 
                           mask_2_9_port);
   mask_reg_2_8_inst : DLH_X1 port map( G => n358, D => n534, Q => 
                           mask_2_8_port);
   mask_reg_2_7_inst : DLH_X1 port map( G => n358, D => n533, Q => 
                           mask_2_7_port);
   mask_reg_2_6_inst : DLH_X1 port map( G => n358, D => n532, Q => 
                           mask_2_6_port);
   mask_reg_2_5_inst : DLH_X1 port map( G => n358, D => n531, Q => 
                           mask_2_5_port);
   mask_reg_2_4_inst : DLH_X1 port map( G => n358, D => n530, Q => 
                           mask_2_4_port);
   mask_reg_2_3_inst : DLH_X1 port map( G => n357, D => n529, Q => 
                           mask_2_3_port);
   mask_reg_2_2_inst : DLH_X1 port map( G => n357, D => n528, Q => 
                           mask_2_2_port);
   mask_reg_2_1_inst : DLH_X1 port map( G => n357, D => n527, Q => 
                           mask_2_1_port);
   mask_reg_2_0_inst : DLH_X1 port map( G => n357, D => n526, Q => 
                           mask_2_0_port);
   mask_reg_3_39_inst : DLH_X1 port map( G => n357, D => n541, Q => 
                           mask_3_39_port);
   mask_reg_3_38_inst : DLH_X1 port map( G => n357, D => N43, Q => 
                           mask_3_38_port);
   mask_reg_3_37_inst : DLH_X1 port map( G => n357, D => N42, Q => 
                           mask_3_37_port);
   mask_reg_3_36_inst : DLH_X1 port map( G => n357, D => N41, Q => 
                           mask_3_36_port);
   mask_reg_3_35_inst : DLH_X1 port map( G => n357, D => N40, Q => 
                           mask_3_35_port);
   mask_reg_3_34_inst : DLH_X1 port map( G => n357, D => N39, Q => 
                           mask_3_34_port);
   mask_reg_3_33_inst : DLH_X1 port map( G => n357, D => N38, Q => 
                           mask_3_33_port);
   mask_reg_3_32_inst : DLH_X1 port map( G => n356, D => N37, Q => 
                           mask_3_32_port);
   mask_reg_3_31_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_31_port);
   mask_reg_3_30_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_30_port);
   mask_reg_3_29_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_29_port);
   mask_reg_3_28_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_28_port);
   mask_reg_3_27_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_27_port);
   mask_reg_3_26_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_26_port);
   mask_reg_3_25_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_25_port);
   mask_reg_3_24_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_24_port);
   mask_reg_3_23_inst : DLH_X1 port map( G => n356, D => n326, Q => 
                           mask_3_23_port);
   mask_reg_3_22_inst : DLH_X1 port map( G => n356, D => n327, Q => 
                           mask_3_22_port);
   mask_reg_3_21_inst : DLH_X1 port map( G => n355, D => n327, Q => 
                           mask_3_21_port);
   mask_reg_3_20_inst : DLH_X1 port map( G => n355, D => n327, Q => 
                           mask_3_20_port);
   mask_reg_3_19_inst : DLH_X1 port map( G => n355, D => n327, Q => 
                           mask_3_19_port);
   mask_reg_3_18_inst : DLH_X1 port map( G => n355, D => n327, Q => 
                           mask_3_18_port);
   mask_reg_3_17_inst : DLH_X1 port map( G => n355, D => n327, Q => 
                           mask_3_17_port);
   mask_reg_3_16_inst : DLH_X1 port map( G => n355, D => n328, Q => 
                           mask_3_16_port);
   mask_reg_3_15_inst : DLH_X1 port map( G => n355, D => n328, Q => 
                           mask_3_15_port);
   mask_reg_3_14_inst : DLH_X1 port map( G => n355, D => n328, Q => 
                           mask_3_14_port);
   mask_reg_3_13_inst : DLH_X1 port map( G => n355, D => n328, Q => 
                           mask_3_13_port);
   mask_reg_3_12_inst : DLH_X1 port map( G => n355, D => n328, Q => 
                           mask_3_12_port);
   mask_reg_3_11_inst : DLH_X1 port map( G => n355, D => n328, Q => 
                           mask_3_11_port);
   mask_reg_3_10_inst : DLH_X1 port map( G => n354, D => n328, Q => 
                           mask_3_10_port);
   mask_reg_3_9_inst : DLH_X1 port map( G => n354, D => n328, Q => 
                           mask_3_9_port);
   mask_reg_3_8_inst : DLH_X1 port map( G => n354, D => n328, Q => 
                           mask_3_8_port);
   mask_reg_3_7_inst : DLH_X1 port map( G => n354, D => N35, Q => mask_3_7_port
                           );
   mask_reg_3_6_inst : DLH_X1 port map( G => n354, D => n540, Q => 
                           mask_3_6_port);
   mask_reg_3_5_inst : DLH_X1 port map( G => n354, D => n539, Q => 
                           mask_3_5_port);
   mask_reg_3_4_inst : DLH_X1 port map( G => n354, D => n538, Q => 
                           mask_3_4_port);
   mask_reg_3_3_inst : DLH_X1 port map( G => n354, D => n537, Q => 
                           mask_3_3_port);
   mask_reg_3_2_inst : DLH_X1 port map( G => n354, D => n536, Q => 
                           mask_3_2_port);
   mask_reg_3_1_inst : DLH_X1 port map( G => n354, D => n535, Q => 
                           mask_3_1_port);
   mask_reg_3_0_inst : DLH_X1 port map( G => n354, D => n534, Q => 
                           mask_3_0_port);
   U3 : BUF_X1 port map( A => n20, Z => n333);
   U4 : AND2_X1 port map( A1 => R(4), A2 => n378, ZN => n1);
   U5 : AND2_X1 port map( A1 => n378, A2 => n379, ZN => n2);
   U6 : AND2_X1 port map( A1 => n301, A2 => n62, ZN => n3);
   U7 : AND2_X1 port map( A1 => n301, A2 => n63, ZN => n4);
   U8 : AND4_X1 port map( A1 => n140, A2 => n141, A3 => n142, A4 => n143, ZN =>
                           n5);
   U9 : AND4_X1 port map( A1 => n148, A2 => n149, A3 => n150, A4 => n151, ZN =>
                           n6);
   U10 : AND4_X1 port map( A1 => n156, A2 => n157, A3 => n158_port, A4 => 
                           n159_port, ZN => n7);
   U11 : AND4_X1 port map( A1 => n160_port, A2 => n130, A3 => n146, A4 => 
                           n109_port, ZN => n8);
   U12 : AND4_X1 port map( A1 => n168_port, A2 => n137, A3 => n154, A4 => n117,
                           ZN => n9);
   U13 : AND4_X1 port map( A1 => n176_port, A2 => n145, A3 => n162_port, A4 => 
                           n127, ZN => n10);
   U14 : AND4_X1 port map( A1 => n136, A2 => n137, A3 => n138, A4 => n139, ZN 
                           => n11);
   U15 : AND4_X1 port map( A1 => n144, A2 => n145, A3 => n146, A4 => n147, ZN 
                           => n12);
   U16 : AND4_X1 port map( A1 => n152, A2 => n153, A3 => n154, A4 => n155, ZN 
                           => n13);
   U17 : AND4_X1 port map( A1 => n160_port, A2 => n161_port, A3 => n162_port, 
                           A4 => n163_port, ZN => n14);
   U18 : AND4_X1 port map( A1 => n156, A2 => n125, A3 => n142, A4 => n102, ZN 
                           => n15);
   U19 : AND4_X1 port map( A1 => n164_port, A2 => n135, A3 => n150, A4 => 
                           n115_port, ZN => n16);
   U20 : AND4_X1 port map( A1 => n172_port, A2 => n141, A3 => n158_port, A4 => 
                           n122, ZN => n17);
   U21 : AND4_X1 port map( A1 => n180_port, A2 => n149, A3 => n166_port, A4 => 
                           n132, ZN => n18);
   U22 : AND2_X1 port map( A1 => R(3), A2 => n379, ZN => n19);
   U23 : BUF_X1 port map( A => n215_port, Z => n305);
   U24 : BUF_X1 port map( A => n339, Z => n334);
   U25 : BUF_X1 port map( A => n375, Z => n370);
   U26 : BUF_X1 port map( A => n375, Z => n369);
   U27 : BUF_X1 port map( A => n374, Z => n373);
   U28 : BUF_X1 port map( A => n374, Z => n372);
   U29 : BUF_X1 port map( A => n374, Z => n371);
   U30 : BUF_X1 port map( A => n333, Z => n338);
   U31 : BUF_X1 port map( A => n353, Z => n374);
   U32 : BUF_X1 port map( A => n56_port, Z => n331);
   U33 : BUF_X1 port map( A => n56_port, Z => n332);
   U34 : BUF_X1 port map( A => n525, Z => n351);
   U35 : BUF_X1 port map( A => n294, Z => n286);
   U36 : BUF_X1 port map( A => n294, Z => n287);
   U37 : BUF_X1 port map( A => R(0), Z => n294);
   U38 : BUF_X1 port map( A => n310, Z => n312);
   U39 : BUF_X1 port map( A => n305, Z => n308);
   U40 : BUF_X1 port map( A => n305, Z => n306);
   U41 : BUF_X1 port map( A => n93_port, Z => n298);
   U42 : BUF_X1 port map( A => n93_port, Z => n299);
   U43 : BUF_X1 port map( A => n93_port, Z => n300);
   U44 : BUF_X1 port map( A => n305, Z => n307);
   U45 : BUF_X1 port map( A => n318, Z => n320);
   U46 : BUF_X1 port map( A => n338, Z => n335);
   U47 : BUF_X1 port map( A => n92_port, Z => n295);
   U48 : BUF_X1 port map( A => n99_port, Z => n303);
   U49 : BUF_X1 port map( A => n99_port, Z => n301);
   U50 : BUF_X1 port map( A => n92_port, Z => n296);
   U51 : BUF_X1 port map( A => n92_port, Z => n297);
   U52 : BUF_X1 port map( A => n99_port, Z => n302);
   U53 : BUF_X1 port map( A => n304, Z => n309);
   U54 : BUF_X1 port map( A => n215_port, Z => n304);
   U55 : BUF_X1 port map( A => n344, Z => n341);
   U56 : BUF_X1 port map( A => n344, Z => n342);
   U57 : BUF_X1 port map( A => n338, Z => n336);
   U58 : BUF_X1 port map( A => n373, Z => n354);
   U59 : BUF_X1 port map( A => n373, Z => n355);
   U60 : BUF_X1 port map( A => n373, Z => n356);
   U61 : BUF_X1 port map( A => n372, Z => n357);
   U62 : BUF_X1 port map( A => n372, Z => n358);
   U63 : BUF_X1 port map( A => n372, Z => n359);
   U64 : BUF_X1 port map( A => n371, Z => n360);
   U65 : BUF_X1 port map( A => n371, Z => n361);
   U66 : BUF_X1 port map( A => n371, Z => n362);
   U67 : BUF_X1 port map( A => n370, Z => n363);
   U68 : BUF_X1 port map( A => n370, Z => n364);
   U69 : BUF_X1 port map( A => n370, Z => n365);
   U70 : BUF_X1 port map( A => n369, Z => n366);
   U71 : BUF_X1 port map( A => n369, Z => n367);
   U72 : BUF_X1 port map( A => n369, Z => n368);
   U73 : BUF_X1 port map( A => n338, Z => n337);
   U74 : BUF_X1 port map( A => n333, Z => n339);
   U75 : NAND2_X1 port map( A1 => n284, A2 => n285, ZN => n96_port);
   U76 : BUF_X1 port map( A => n286, Z => n293);
   U77 : BUF_X1 port map( A => n287, Z => n290);
   U78 : BUF_X1 port map( A => n286, Z => n291);
   U79 : BUF_X1 port map( A => n345, Z => n340);
   U80 : BUF_X1 port map( A => n19, Z => n345);
   U81 : BUF_X1 port map( A => n19, Z => n344);
   U82 : BUF_X1 port map( A => n287, Z => n289);
   U83 : BUF_X1 port map( A => n286, Z => n292);
   U84 : BUF_X1 port map( A => n352, Z => n346);
   U85 : BUF_X1 port map( A => n352, Z => n347);
   U86 : BUF_X1 port map( A => n351, Z => n348);
   U87 : BUF_X1 port map( A => n351, Z => n349);
   U88 : INV_X1 port map( A => n331, ZN => n329);
   U89 : INV_X1 port map( A => n331, ZN => n330);
   U90 : BUF_X1 port map( A => n332, Z => n327);
   U91 : BUF_X1 port map( A => n332, Z => n326);
   U92 : BUF_X1 port map( A => n332, Z => n328);
   U93 : BUF_X1 port map( A => n351, Z => n350);
   U94 : BUF_X1 port map( A => n287, Z => n288);
   U95 : AND2_X1 port map( A1 => R(3), A2 => R(4), ZN => n20);
   U96 : AND3_X1 port map( A1 => n230, A2 => n231, A3 => n232, ZN => n21);
   U97 : AND4_X1 port map( A1 => n188_port, A2 => n189_port, A3 => n190_port, 
                           A4 => n191_port, ZN => n22);
   U98 : AND4_X1 port map( A1 => n184_port, A2 => n185_port, A3 => n186_port, 
                           A4 => n187_port, ZN => n23);
   U99 : AND3_X1 port map( A1 => n220_port, A2 => n221_port, A3 => n222, ZN => 
                           n24);
   U100 : AND3_X1 port map( A1 => n224, A2 => n225, A3 => n226, ZN => n25);
   U101 : AND4_X1 port map( A1 => n212_port, A2 => n181_port, A3 => n198_port, 
                           A4 => n167_port, ZN => n26);
   U102 : AND4_X1 port map( A1 => n220_port, A2 => n185_port, A3 => n202_port, 
                           A4 => n171_port, ZN => n27);
   U103 : AND4_X1 port map( A1 => n224, A2 => n189_port, A3 => n206_port, A4 =>
                           n175_port, ZN => n28_port);
   U104 : AND4_X1 port map( A1 => n230, A2 => n193_port, A3 => n210_port, A4 =>
                           n179_port, ZN => n29);
   U105 : AND4_X1 port map( A1 => n196_port, A2 => n197_port, A3 => n198_port, 
                           A4 => n199_port, ZN => n30);
   U106 : AND4_X1 port map( A1 => n192_port, A2 => n193_port, A3 => n194_port, 
                           A4 => n195_port, ZN => n31);
   U107 : AND3_X1 port map( A1 => n247, A2 => n199_port, A3 => n269, ZN => n32)
                           ;
   U108 : AND3_X1 port map( A1 => n235, A2 => n195_port, A3 => n266, ZN => n33)
                           ;
   U109 : AND3_X1 port map( A1 => n212_port, A2 => n213_port, A3 => n214_port, 
                           ZN => n34);
   U110 : AND4_X1 port map( A1 => n243, A2 => n197_port, A3 => n218_port, A4 =>
                           n183_port, ZN => n35_port);
   U111 : AND4_X1 port map( A1 => n200_port, A2 => n201_port, A3 => n202_port, 
                           A4 => n203_port, ZN => n36);
   U112 : AND4_X1 port map( A1 => n204_port, A2 => n205_port, A3 => n206_port, 
                           A4 => n207_port, ZN => n37_port);
   U113 : AND4_X1 port map( A1 => n208_port, A2 => n209_port, A3 => n210_port, 
                           A4 => n211_port, ZN => n38_port);
   U114 : INV_X1 port map( A => n229, ZN => n488);
   U115 : AND4_X1 port map( A1 => n184_port, A2 => n153, A3 => n170_port, A4 =>
                           n139, ZN => n39_port);
   U116 : AND4_X1 port map( A1 => n188_port, A2 => n157, A3 => n174_port, A4 =>
                           n143, ZN => n40_port);
   U117 : AND4_X1 port map( A1 => n164_port, A2 => n165_port, A3 => n166_port, 
                           A4 => n167_port, ZN => n41_port);
   U118 : AND4_X1 port map( A1 => n192_port, A2 => n161_port, A3 => n178_port, 
                           A4 => n147, ZN => n42_port);
   U119 : AND4_X1 port map( A1 => n168_port, A2 => n169_port, A3 => n170_port, 
                           A4 => n171_port, ZN => n43_port);
   U120 : AND4_X1 port map( A1 => n196_port, A2 => n165_port, A3 => n182_port, 
                           A4 => n151, ZN => n44);
   U121 : AND4_X1 port map( A1 => n172_port, A2 => n173_port, A3 => n174_port, 
                           A4 => n175_port, ZN => n45);
   U122 : AND4_X1 port map( A1 => n200_port, A2 => n169_port, A3 => n186_port, 
                           A4 => n155, ZN => n46);
   U123 : AND4_X1 port map( A1 => n176_port, A2 => n177_port, A3 => n178_port, 
                           A4 => n179_port, ZN => n47);
   U124 : AND4_X1 port map( A1 => n204_port, A2 => n173_port, A3 => n190_port, 
                           A4 => n159_port, ZN => n48);
   U125 : AND4_X1 port map( A1 => n180_port, A2 => n181_port, A3 => n182_port, 
                           A4 => n183_port, ZN => n49);
   U126 : AND4_X1 port map( A1 => n208_port, A2 => n177_port, A3 => n194_port, 
                           A4 => n163_port, ZN => n50);
   U127 : AND3_X1 port map( A1 => n140, A2 => n97_port, A3 => n254, ZN => n51);
   U128 : AND3_X1 port map( A1 => n144, A2 => n105, A3 => n256, ZN => n52);
   U129 : AND3_X1 port map( A1 => n116_port, A2 => n117, A3 => n118, ZN => 
                           n53_port);
   U130 : AND3_X1 port map( A1 => n148, A2 => n111_port, A3 => n258, ZN => 
                           n54_port);
   U131 : AND3_X1 port map( A1 => n121, A2 => n122, A3 => n123, ZN => n55_port)
                           ;
   U132 : BUF_X1 port map( A => n525, Z => n352);
   U133 : BUF_X1 port map( A => n353, Z => n375);
   U134 : NOR2_X1 port map( A1 => n3, A2 => n264, ZN => n262);
   U135 : OAI211_X1 port map( C1 => out_mask_32_port, C2 => n96_port, A => 
                           n201_port, B => n187_port, ZN => n264);
   U136 : NOR2_X1 port map( A1 => n4, A2 => n265, ZN => n263);
   U137 : OAI211_X1 port map( C1 => out_mask_33_port, C2 => n96_port, A => 
                           n205_port, B => n191_port, ZN => n265);
   U138 : NOR2_X1 port map( A1 => n239, A2 => n238, ZN => n229);
   U139 : AND2_X1 port map( A1 => data_in(31), A2 => n238, ZN => n56_port);
   U140 : NAND2_X1 port map( A1 => n239, A2 => data_in(31), ZN => n219_port);
   U141 : AND3_X1 port map( A1 => n152, A2 => n120, A3 => n260, ZN => n57_port)
                           ;
   U142 : AND3_X1 port map( A1 => n126, A2 => n127, A3 => n128, ZN => n58_port)
                           ;
   U143 : AND3_X1 port map( A1 => n131, A2 => n132, A3 => n133, ZN => n59_port)
                           ;
   U144 : BUF_X1 port map( A => N28, Z => n353);
   U145 : AND2_X1 port map( A1 => n418, A2 => n417, ZN => n60_port);
   U146 : AND2_X1 port map( A1 => n421, A2 => n420, ZN => n61);
   U147 : AND2_X1 port map( A1 => n409, A2 => n408, ZN => n62);
   U148 : AND2_X1 port map( A1 => n406, A2 => n405, ZN => n63);
   U149 : AND2_X1 port map( A1 => n431, A2 => n430, ZN => n64);
   U150 : AND2_X1 port map( A1 => n434, A2 => n433, ZN => n65);
   U151 : AND2_X1 port map( A1 => n437, A2 => n436, ZN => n66);
   U152 : AND2_X1 port map( A1 => n427, A2 => n426, ZN => n67);
   U153 : AND2_X1 port map( A1 => n424, A2 => n423, ZN => n68_port);
   U154 : AND2_X1 port map( A1 => n440, A2 => n439, ZN => n69_port);
   U155 : AND2_X1 port map( A1 => n415, A2 => n414, ZN => n70_port);
   U156 : AND2_X1 port map( A1 => n412, A2 => n411, ZN => n71_port);
   U157 : NOR2_X1 port map( A1 => n598, A2 => conf(1), ZN => n239);
   U158 : OR2_X1 port map( A1 => conf(0), A2 => conf(1), ZN => n400);
   U159 : AND2_X1 port map( A1 => n500, A2 => n499, ZN => n72_port);
   U160 : AND2_X1 port map( A1 => n496, A2 => n495, ZN => n73_port);
   U161 : AND2_X1 port map( A1 => n492, A2 => n491, ZN => n74_port);
   U162 : AND2_X1 port map( A1 => n486, A2 => n485, ZN => n75_port);
   U163 : AND2_X1 port map( A1 => n481, A2 => n480, ZN => n76_port);
   U164 : AND2_X1 port map( A1 => n476, A2 => n475, ZN => n77_port);
   U165 : AND2_X1 port map( A1 => n471, A2 => n470, ZN => n78_port);
   U166 : AND2_X1 port map( A1 => n466, A2 => n465, ZN => n79_port);
   U167 : AND2_X1 port map( A1 => n461, A2 => n460, ZN => n80_port);
   U168 : AND2_X1 port map( A1 => n456, A2 => n455, ZN => n81_port);
   U169 : AND2_X1 port map( A1 => n452, A2 => n451, ZN => n82_port);
   U170 : AND2_X1 port map( A1 => n449, A2 => n448, ZN => n83_port);
   U171 : AND2_X1 port map( A1 => n446, A2 => n445, ZN => n84);
   U172 : AND2_X1 port map( A1 => n443, A2 => n442, ZN => n85_port);
   U173 : AND2_X1 port map( A1 => conf(1), A2 => n598, ZN => n238);
   U174 : INV_X1 port map( A => conf(0), ZN => n598);
   U175 : MUX2_X1 port map( A => n86_port, B => n87_port, S => n288, Z => N190)
                           ;
   U176 : OAI221_X1 port map( B1 => n88_port, B2 => n72_port, C1 => n89_port, 
                           C2 => n90_port, A => n91_port, ZN => n86_port);
   U177 : AOI22_X1 port map( A1 => out_mask_4_port, A2 => n297, B1 => 
                           out_mask_0_port, B2 => n300, ZN => n91_port);
   U178 : MUX2_X1 port map( A => n87_port, B => n94_port, S => n288, Z => N191)
                           ;
   U179 : INV_X1 port map( A => n95_port, ZN => n87_port);
   U180 : OAI211_X1 port map( C1 => out_mask_1_port, C2 => n96_port, A => 
                           n97_port, B => n98_port, ZN => n95_port);
   U181 : AOI21_X1 port map( B1 => n303, B2 => n100, A => n101, ZN => n98_port)
                           ;
   U182 : INV_X1 port map( A => n102, ZN => n101);
   U183 : MUX2_X1 port map( A => n94_port, B => n103, S => n288, Z => N192);
   U184 : INV_X1 port map( A => n104, ZN => n94_port);
   U185 : OAI211_X1 port map( C1 => out_mask_2_port, C2 => n96_port, A => n105,
                           B => n106, ZN => n104);
   U186 : AOI21_X1 port map( B1 => n303, B2 => n107, A => n108_port, ZN => n106
                           );
   U187 : INV_X1 port map( A => n109_port, ZN => n108_port);
   U188 : MUX2_X1 port map( A => n103, B => n53_port, S => n288, Z => N193);
   U189 : INV_X1 port map( A => n110_port, ZN => n103);
   U190 : OAI211_X1 port map( C1 => out_mask_3_port, C2 => n96_port, A => 
                           n111_port, B => n112_port, ZN => n110_port);
   U191 : AOI21_X1 port map( B1 => n303, B2 => n113_port, A => n114_port, ZN =>
                           n112_port);
   U192 : INV_X1 port map( A => n115_port, ZN => n114_port);
   U193 : MUX2_X1 port map( A => n53_port, B => n55_port, S => n289, Z => N194)
                           ;
   U194 : AOI21_X1 port map( B1 => n300, B2 => n107, A => n119, ZN => n118);
   U195 : INV_X1 port map( A => n120, ZN => n119);
   U196 : MUX2_X1 port map( A => n55_port, B => n58_port, S => n289, Z => N195)
                           ;
   U197 : AOI21_X1 port map( B1 => n300, B2 => n113_port, A => n124, ZN => n123
                           );
   U198 : INV_X1 port map( A => n125, ZN => n124);
   U199 : MUX2_X1 port map( A => n58_port, B => n59_port, S => n289, Z => N196)
                           ;
   U200 : AOI21_X1 port map( B1 => n300, B2 => n72_port, A => n129, ZN => n128)
                           ;
   U201 : INV_X1 port map( A => n130, ZN => n129);
   U202 : MUX2_X1 port map( A => n59_port, B => n11, S => n289, Z => N197);
   U203 : AOI21_X1 port map( B1 => n300, B2 => n73_port, A => n134, ZN => n133)
                           ;
   U204 : INV_X1 port map( A => n135, ZN => n134);
   U205 : MUX2_X1 port map( A => n11, B => n5, S => n289, Z => N198);
   U206 : MUX2_X1 port map( A => n5, B => n12, S => n289, Z => N199);
   U207 : MUX2_X1 port map( A => n12, B => n6, S => n289, Z => N200);
   U208 : MUX2_X1 port map( A => n6, B => n13, S => n289, Z => N201);
   U209 : MUX2_X1 port map( A => n13, B => n7, S => n289, Z => N202);
   U210 : MUX2_X1 port map( A => n7, B => n14, S => n289, Z => N203);
   U211 : MUX2_X1 port map( A => n14, B => n41_port, S => n289, Z => N204);
   U212 : MUX2_X1 port map( A => n41_port, B => n43_port, S => n289, Z => N205)
                           ;
   U213 : MUX2_X1 port map( A => n43_port, B => n45, S => n290, Z => N206);
   U214 : MUX2_X1 port map( A => n45, B => n47, S => n290, Z => N207);
   U215 : MUX2_X1 port map( A => n47, B => n49, S => n290, Z => N208);
   U216 : MUX2_X1 port map( A => n49, B => n23, S => n290, Z => N209);
   U217 : MUX2_X1 port map( A => n23, B => n22, S => n290, Z => N210);
   U218 : MUX2_X1 port map( A => n22, B => n31, S => n290, Z => N211);
   U219 : MUX2_X1 port map( A => n31, B => n30, S => n290, Z => N212);
   U220 : MUX2_X1 port map( A => n30, B => n36, S => n290, Z => N213);
   U221 : MUX2_X1 port map( A => n36, B => n37_port, S => n290, Z => N214);
   U222 : MUX2_X1 port map( A => n37_port, B => n38_port, S => n290, Z => N215)
                           ;
   U223 : MUX2_X1 port map( A => n38_port, B => n34, S => n290, Z => N216);
   U224 : MUX2_X1 port map( A => n34, B => n24, S => n290, Z => N217);
   U225 : AOI21_X1 port map( B1 => n309, B2 => n216_port, A => n217_port, ZN =>
                           n214_port);
   U226 : INV_X1 port map( A => n218_port, ZN => n217_port);
   U227 : MUX2_X1 port map( A => n24, B => n25, S => n291, Z => N218);
   U228 : AOI21_X1 port map( B1 => n309, B2 => n223, A => n3, ZN => n222);
   U229 : MUX2_X1 port map( A => n25, B => n21, S => n291, Z => N219);
   U230 : AOI21_X1 port map( B1 => n309, B2 => n227, A => n4, ZN => n226);
   U231 : MUX2_X1 port map( A => n21, B => n228, S => n291, Z => N220);
   U232 : AOI21_X1 port map( B1 => n309, B2 => n233, A => n234, ZN => n232);
   U233 : INV_X1 port map( A => n235, ZN => n234);
   U234 : MUX2_X1 port map( A => n228, B => n236, S => n291, Z => N221);
   U235 : OAI221_X1 port map( B1 => n237, B2 => n233, C1 => n96_port, C2 => 
                           n240, A => n241, ZN => n236);
   U236 : AOI22_X1 port map( A1 => out_mask_38_port, A2 => n309, B1 => 
                           out_mask_34_port, B2 => n303, ZN => n241);
   U237 : INV_X1 port map( A => n242, ZN => n228);
   U238 : OAI211_X1 port map( C1 => out_mask_35_port, C2 => n237, A => n243, B 
                           => n244, ZN => n242);
   U239 : AOI21_X1 port map( B1 => n309, B2 => n245, A => n246, ZN => n244);
   U240 : INV_X1 port map( A => n247, ZN => n246);
   U241 : MUX2_X1 port map( A => n248, B => n249, S => n291, Z => N158);
   U242 : OAI221_X1 port map( B1 => n237, B2 => n100, C1 => n96_port, C2 => 
                           n73_port, A => n250, ZN => n249);
   U243 : AOI22_X1 port map( A1 => out_mask_1_port, A2 => n309, B1 => 
                           out_mask_5_port, B2 => n303, ZN => n250);
   U244 : MUX2_X1 port map( A => n51, B => n248, S => n291, Z => N159);
   U245 : INV_X1 port map( A => n251, ZN => n248);
   U246 : OAI211_X1 port map( C1 => out_mask_4_port, C2 => n237, A => n136, B 
                           => n252, ZN => n251);
   U247 : AOI21_X1 port map( B1 => n309, B2 => n90_port, A => n253, ZN => n252)
                           ;
   U248 : INV_X1 port map( A => n116_port, ZN => n253);
   U249 : NAND2_X1 port map( A1 => n303, A2 => n72_port, ZN => n116_port);
   U250 : INV_X1 port map( A => out_mask_2_port, ZN => n90_port);
   U251 : NAND2_X1 port map( A1 => n300, A2 => n74_port, ZN => n136);
   U252 : MUX2_X1 port map( A => n52, B => n51, S => n291, Z => N160);
   U253 : AOI21_X1 port map( B1 => n309, B2 => n100, A => n255, ZN => n254);
   U254 : INV_X1 port map( A => n121, ZN => n255);
   U255 : NAND2_X1 port map( A1 => n303, A2 => n73_port, ZN => n121);
   U256 : INV_X1 port map( A => out_mask_3_port, ZN => n100);
   U257 : NAND2_X1 port map( A1 => n297, A2 => n113_port, ZN => n97_port);
   U258 : NAND2_X1 port map( A1 => n300, A2 => n75_port, ZN => n140);
   U259 : MUX2_X1 port map( A => n54_port, B => n52, S => n291, Z => N161);
   U260 : AOI21_X1 port map( B1 => n309, B2 => n107, A => n257, ZN => n256);
   U261 : INV_X1 port map( A => n126, ZN => n257);
   U262 : NAND2_X1 port map( A1 => n303, A2 => n74_port, ZN => n126);
   U263 : INV_X1 port map( A => out_mask_4_port, ZN => n107);
   U264 : NAND2_X1 port map( A1 => n297, A2 => n72_port, ZN => n105);
   U265 : NAND2_X1 port map( A1 => n300, A2 => n76_port, ZN => n144);
   U266 : MUX2_X1 port map( A => n57_port, B => n54_port, S => n291, Z => N162)
                           ;
   U267 : AOI21_X1 port map( B1 => n309, B2 => n113_port, A => n259, ZN => n258
                           );
   U268 : INV_X1 port map( A => n131, ZN => n259);
   U269 : NAND2_X1 port map( A1 => n302, A2 => n75_port, ZN => n131);
   U270 : INV_X1 port map( A => out_mask_5_port, ZN => n113_port);
   U271 : NAND2_X1 port map( A1 => n297, A2 => n73_port, ZN => n111_port);
   U272 : NAND2_X1 port map( A1 => n299, A2 => n77_port, ZN => n148);
   U273 : MUX2_X1 port map( A => n15, B => n57_port, S => n291, Z => N163);
   U274 : AOI21_X1 port map( B1 => n309, B2 => n72_port, A => n261, ZN => n260)
                           ;
   U275 : INV_X1 port map( A => n138, ZN => n261);
   U276 : NAND2_X1 port map( A1 => n302, A2 => n76_port, ZN => n138);
   U277 : NAND2_X1 port map( A1 => n297, A2 => n74_port, ZN => n120);
   U278 : NAND2_X1 port map( A1 => n299, A2 => n78_port, ZN => n152);
   U279 : MUX2_X1 port map( A => n8, B => n15, S => n291, Z => N164);
   U280 : NAND2_X1 port map( A1 => n308, A2 => n73_port, ZN => n102);
   U281 : NAND2_X1 port map( A1 => n302, A2 => n77_port, ZN => n142);
   U282 : NAND2_X1 port map( A1 => n297, A2 => n75_port, ZN => n125);
   U283 : NAND2_X1 port map( A1 => n299, A2 => n79_port, ZN => n156);
   U284 : MUX2_X1 port map( A => n16, B => n8, S => n291, Z => N165);
   U285 : NAND2_X1 port map( A1 => n308, A2 => n74_port, ZN => n109_port);
   U286 : NAND2_X1 port map( A1 => n302, A2 => n78_port, ZN => n146);
   U287 : NAND2_X1 port map( A1 => n297, A2 => n76_port, ZN => n130);
   U288 : NAND2_X1 port map( A1 => n299, A2 => n80_port, ZN => n160_port);
   U289 : MUX2_X1 port map( A => n9, B => n16, S => n292, Z => N166);
   U290 : NAND2_X1 port map( A1 => n308, A2 => n75_port, ZN => n115_port);
   U291 : NAND2_X1 port map( A1 => n302, A2 => n79_port, ZN => n150);
   U292 : NAND2_X1 port map( A1 => n297, A2 => n77_port, ZN => n135);
   U293 : NAND2_X1 port map( A1 => n299, A2 => n81_port, ZN => n164_port);
   U294 : MUX2_X1 port map( A => n17, B => n9, S => n292, Z => N167);
   U295 : NAND2_X1 port map( A1 => n308, A2 => n76_port, ZN => n117);
   U296 : NAND2_X1 port map( A1 => n302, A2 => n80_port, ZN => n154);
   U297 : NAND2_X1 port map( A1 => n296, A2 => n78_port, ZN => n137);
   U298 : NAND2_X1 port map( A1 => n299, A2 => n82_port, ZN => n168_port);
   U299 : MUX2_X1 port map( A => n10, B => n17, S => n292, Z => N168);
   U300 : NAND2_X1 port map( A1 => n308, A2 => n77_port, ZN => n122);
   U301 : NAND2_X1 port map( A1 => n302, A2 => n81_port, ZN => n158_port);
   U302 : NAND2_X1 port map( A1 => n297, A2 => n79_port, ZN => n141);
   U303 : NAND2_X1 port map( A1 => n299, A2 => n83_port, ZN => n172_port);
   U304 : MUX2_X1 port map( A => n18, B => n10, S => n292, Z => N169);
   U305 : NAND2_X1 port map( A1 => n308, A2 => n78_port, ZN => n127);
   U306 : NAND2_X1 port map( A1 => n302, A2 => n82_port, ZN => n162_port);
   U307 : NAND2_X1 port map( A1 => n297, A2 => n80_port, ZN => n145);
   U308 : NAND2_X1 port map( A1 => n299, A2 => n84, ZN => n176_port);
   U309 : MUX2_X1 port map( A => n39_port, B => n18, S => n292, Z => N170);
   U310 : NAND2_X1 port map( A1 => n308, A2 => n79_port, ZN => n132);
   U311 : NAND2_X1 port map( A1 => n302, A2 => n83_port, ZN => n166_port);
   U312 : NAND2_X1 port map( A1 => n296, A2 => n81_port, ZN => n149);
   U313 : NAND2_X1 port map( A1 => n299, A2 => n85_port, ZN => n180_port);
   U314 : MUX2_X1 port map( A => n40_port, B => n39_port, S => n292, Z => N171)
                           ;
   U315 : NAND2_X1 port map( A1 => n308, A2 => n80_port, ZN => n139);
   U316 : NAND2_X1 port map( A1 => n302, A2 => n84, ZN => n170_port);
   U317 : NAND2_X1 port map( A1 => n296, A2 => n82_port, ZN => n153);
   U318 : NAND2_X1 port map( A1 => n299, A2 => n69_port, ZN => n184_port);
   U319 : MUX2_X1 port map( A => n42_port, B => n40_port, S => n292, Z => N172)
                           ;
   U320 : NAND2_X1 port map( A1 => n308, A2 => n81_port, ZN => n143);
   U321 : NAND2_X1 port map( A1 => n302, A2 => n85_port, ZN => n174_port);
   U322 : NAND2_X1 port map( A1 => n296, A2 => n83_port, ZN => n157);
   U323 : NAND2_X1 port map( A1 => n299, A2 => n66, ZN => n188_port);
   U324 : MUX2_X1 port map( A => n44, B => n42_port, S => n292, Z => N173);
   U325 : NAND2_X1 port map( A1 => n308, A2 => n82_port, ZN => n147);
   U326 : NAND2_X1 port map( A1 => n301, A2 => n69_port, ZN => n178_port);
   U327 : NAND2_X1 port map( A1 => n296, A2 => n84, ZN => n161_port);
   U328 : NAND2_X1 port map( A1 => n298, A2 => n65, ZN => n192_port);
   U329 : MUX2_X1 port map( A => n46, B => n44, S => n292, Z => N174);
   U330 : NAND2_X1 port map( A1 => n307, A2 => n83_port, ZN => n151);
   U331 : NAND2_X1 port map( A1 => n301, A2 => n66, ZN => n182_port);
   U332 : NAND2_X1 port map( A1 => n296, A2 => n85_port, ZN => n165_port);
   U333 : NAND2_X1 port map( A1 => n298, A2 => n64, ZN => n196_port);
   U334 : MUX2_X1 port map( A => n48, B => n46, S => n292, Z => N175);
   U335 : NAND2_X1 port map( A1 => n307, A2 => n84, ZN => n155);
   U336 : NAND2_X1 port map( A1 => n301, A2 => n65, ZN => n186_port);
   U337 : NAND2_X1 port map( A1 => n296, A2 => n69_port, ZN => n169_port);
   U338 : NAND2_X1 port map( A1 => n298, A2 => n67, ZN => n200_port);
   U339 : MUX2_X1 port map( A => n50, B => n48, S => n292, Z => N176);
   U340 : NAND2_X1 port map( A1 => n307, A2 => n85_port, ZN => n159_port);
   U341 : NAND2_X1 port map( A1 => n301, A2 => n64, ZN => n190_port);
   U342 : NAND2_X1 port map( A1 => n296, A2 => n66, ZN => n173_port);
   U343 : NAND2_X1 port map( A1 => n298, A2 => n68_port, ZN => n204_port);
   U344 : MUX2_X1 port map( A => n26, B => n50, S => n292, Z => N177);
   U345 : NAND2_X1 port map( A1 => n307, A2 => n69_port, ZN => n163_port);
   U346 : NAND2_X1 port map( A1 => n301, A2 => n67, ZN => n194_port);
   U347 : NAND2_X1 port map( A1 => n296, A2 => n65, ZN => n177_port);
   U348 : NAND2_X1 port map( A1 => n299, A2 => n61, ZN => n208_port);
   U349 : MUX2_X1 port map( A => n27, B => n26, S => n293, Z => N178);
   U350 : NAND2_X1 port map( A1 => n307, A2 => n66, ZN => n167_port);
   U351 : NAND2_X1 port map( A1 => n301, A2 => n68_port, ZN => n198_port);
   U352 : NAND2_X1 port map( A1 => n296, A2 => n64, ZN => n181_port);
   U353 : NAND2_X1 port map( A1 => n298, A2 => n60_port, ZN => n212_port);
   U354 : MUX2_X1 port map( A => n28_port, B => n27, S => n293, Z => N179);
   U355 : NAND2_X1 port map( A1 => n307, A2 => n65, ZN => n171_port);
   U356 : NAND2_X1 port map( A1 => n301, A2 => n61, ZN => n202_port);
   U357 : NAND2_X1 port map( A1 => n296, A2 => n67, ZN => n185_port);
   U358 : NAND2_X1 port map( A1 => n298, A2 => n70_port, ZN => n220_port);
   U359 : MUX2_X1 port map( A => n29, B => n28_port, S => n293, Z => N180);
   U360 : NAND2_X1 port map( A1 => n307, A2 => n64, ZN => n175_port);
   U361 : NAND2_X1 port map( A1 => n301, A2 => n60_port, ZN => n206_port);
   U362 : NAND2_X1 port map( A1 => n296, A2 => n68_port, ZN => n189_port);
   U363 : NAND2_X1 port map( A1 => n298, A2 => n71_port, ZN => n224);
   U364 : MUX2_X1 port map( A => n35_port, B => n29, S => n293, Z => N181);
   U365 : NAND2_X1 port map( A1 => n307, A2 => n67, ZN => n179_port);
   U366 : NAND2_X1 port map( A1 => n302, A2 => n70_port, ZN => n210_port);
   U367 : NAND2_X1 port map( A1 => n295, A2 => n61, ZN => n193_port);
   U368 : NAND2_X1 port map( A1 => n298, A2 => n62, ZN => n230);
   U369 : MUX2_X1 port map( A => n262, B => n35_port, S => n293, Z => N182);
   U370 : NAND2_X1 port map( A1 => n307, A2 => n68_port, ZN => n183_port);
   U371 : NAND2_X1 port map( A1 => n301, A2 => n71_port, ZN => n218_port);
   U372 : NAND2_X1 port map( A1 => n295, A2 => n60_port, ZN => n197_port);
   U373 : NAND2_X1 port map( A1 => n300, A2 => n63, ZN => n243);
   U374 : MUX2_X1 port map( A => n263, B => n262, S => n293, Z => N183);
   U375 : NAND2_X1 port map( A1 => n307, A2 => n61, ZN => n187_port);
   U376 : NAND2_X1 port map( A1 => n295, A2 => n70_port, ZN => n201_port);
   U377 : MUX2_X1 port map( A => n33, B => n263, S => n293, Z => N184);
   U378 : NAND2_X1 port map( A1 => n307, A2 => n60_port, ZN => n191_port);
   U379 : NAND2_X1 port map( A1 => n295, A2 => n71_port, ZN => n205_port);
   U380 : MUX2_X1 port map( A => n32, B => n33, S => n293, Z => N185);
   U381 : AOI21_X1 port map( B1 => n300, B2 => n223, A => n267, ZN => n266);
   U382 : INV_X1 port map( A => n209_port, ZN => n267);
   U383 : NAND2_X1 port map( A1 => n295, A2 => n62, ZN => n209_port);
   U384 : NAND2_X1 port map( A1 => n307, A2 => n70_port, ZN => n195_port);
   U385 : NAND2_X1 port map( A1 => n301, A2 => n240, ZN => n235);
   U386 : MUX2_X1 port map( A => n268, B => n32, S => n293, Z => N186);
   U387 : AOI21_X1 port map( B1 => n300, B2 => n227, A => n270, ZN => n269);
   U388 : INV_X1 port map( A => n213_port, ZN => n270);
   U389 : NAND2_X1 port map( A1 => n295, A2 => n63, ZN => n213_port);
   U390 : NAND2_X1 port map( A1 => n306, A2 => n71_port, ZN => n199_port);
   U391 : NAND2_X1 port map( A1 => n303, A2 => n216_port, ZN => n247);
   U392 : MUX2_X1 port map( A => n271, B => n268, S => n293, Z => N187);
   U393 : INV_X1 port map( A => n272, ZN => n268);
   U394 : OAI211_X1 port map( C1 => out_mask_36_port, C2 => n96_port, A => 
                           n221_port, B => n273, ZN => n272);
   U395 : AOI21_X1 port map( B1 => n303, B2 => n223, A => n274, ZN => n273);
   U396 : INV_X1 port map( A => n203_port, ZN => n274);
   U397 : NAND2_X1 port map( A1 => n306, A2 => n62, ZN => n203_port);
   U398 : NAND2_X1 port map( A1 => n295, A2 => n240, ZN => n221_port);
   U399 : MUX2_X1 port map( A => n275, B => n271, S => n293, Z => N188);
   U400 : INV_X1 port map( A => n276, ZN => n271);
   U401 : OAI211_X1 port map( C1 => out_mask_37_port, C2 => n96_port, A => n225
                           , B => n277, ZN => n276);
   U402 : AOI21_X1 port map( B1 => n303, B2 => n227, A => n278, ZN => n277);
   U403 : INV_X1 port map( A => n207_port, ZN => n278);
   U404 : NAND2_X1 port map( A1 => n308, A2 => n63, ZN => n207_port);
   U405 : INV_X1 port map( A => out_mask_35_port, ZN => n227);
   U406 : NAND2_X1 port map( A1 => n295, A2 => n216_port, ZN => n225);
   U407 : MUX2_X1 port map( A => n279, B => n275, S => n293, Z => N189);
   U408 : INV_X1 port map( A => n280, ZN => n275);
   U409 : OAI211_X1 port map( C1 => out_mask_38_port, C2 => n96_port, A => n231
                           , B => n281, ZN => n280);
   U410 : AOI21_X1 port map( B1 => n303, B2 => n233, A => n282, ZN => n281);
   U411 : INV_X1 port map( A => n211_port, ZN => n282);
   U412 : NAND2_X1 port map( A1 => n308, A2 => n240, ZN => n211_port);
   U413 : INV_X1 port map( A => out_mask_32_port, ZN => n240);
   U414 : INV_X1 port map( A => n88_port, ZN => n215_port);
   U415 : INV_X1 port map( A => out_mask_36_port, ZN => n233);
   U416 : INV_X1 port map( A => n89_port, ZN => n99_port);
   U417 : NAND2_X1 port map( A1 => n297, A2 => n223, ZN => n231);
   U418 : INV_X1 port map( A => out_mask_34_port, ZN => n223);
   U419 : OAI221_X1 port map( B1 => n88_port, B2 => n216_port, C1 => n89_port, 
                           C2 => n245, A => n283, ZN => n279);
   U420 : AOI22_X1 port map( A1 => out_mask_35_port, A2 => n297, B1 => 
                           out_mask_39_port, B2 => n300, ZN => n283);
   U421 : INV_X1 port map( A => n96_port, ZN => n93_port);
   U422 : INV_X1 port map( A => n237, ZN => n92_port);
   U423 : NAND2_X1 port map( A1 => R(2), A2 => n284, ZN => n237);
   U424 : INV_X1 port map( A => R(1), ZN => n284);
   U425 : INV_X1 port map( A => out_mask_37_port, ZN => n245);
   U426 : NAND2_X1 port map( A1 => R(1), A2 => n285, ZN => n89_port);
   U427 : INV_X1 port map( A => R(2), ZN => n285);
   U428 : INV_X1 port map( A => out_mask_33_port, ZN => n216_port);
   U429 : NAND2_X1 port map( A1 => R(1), A2 => R(2), ZN => n88_port);
   U430 : CLKBUF_X1 port map( A => n315, Z => n310);
   U431 : BUF_X1 port map( A => n2, Z => n311);
   U432 : BUF_X1 port map( A => n310, Z => n313);
   U433 : BUF_X1 port map( A => n310, Z => n314);
   U434 : BUF_X1 port map( A => n311, Z => n315);
   U435 : BUF_X1 port map( A => n311, Z => n316);
   U436 : CLKBUF_X1 port map( A => n311, Z => n317);
   U437 : CLKBUF_X1 port map( A => n323, Z => n318);
   U438 : BUF_X1 port map( A => n1, Z => n319);
   U439 : BUF_X1 port map( A => n318, Z => n321);
   U440 : BUF_X1 port map( A => n318, Z => n322);
   U441 : BUF_X1 port map( A => n319, Z => n323);
   U442 : BUF_X1 port map( A => n319, Z => n324);
   U443 : CLKBUF_X1 port map( A => n319, Z => n325);
   U444 : BUF_X1 port map( A => n344, Z => n343);
   U445 : NAND2_X1 port map( A1 => n229, A2 => n400, ZN => N28);
   U446 : INV_X1 port map( A => n400, ZN => n525);
   U447 : NAND2_X1 port map( A1 => n350, A2 => data_in(15), ZN => n428);
   U448 : NAND2_X1 port map( A1 => n330, A2 => n428, ZN => N60);
   U449 : NAND2_X1 port map( A1 => n350, A2 => data_in(7), ZN => n453);
   U450 : NAND2_X1 port map( A1 => n453, A2 => n329, ZN => n541);
   U451 : INV_X1 port map( A => data_in(31), ZN => n376);
   U452 : OAI21_X1 port map( B1 => n400, B2 => n376, A => n329, ZN => n542);
   U453 : INV_X1 port map( A => data_in(23), ZN => n377);
   U454 : OAI21_X1 port map( B1 => n377, B2 => n400, A => n329, ZN => n550);
   U455 : INV_X1 port map( A => R(3), ZN => n378);
   U456 : AOI22_X1 port map( A1 => mask_2_39_port, A2 => n324, B1 => 
                           mask_3_39_port, B2 => n334, ZN => n381);
   U457 : INV_X1 port map( A => R(4), ZN => n379);
   U458 : AOI22_X1 port map( A1 => mask_0_39_port, A2 => n316, B1 => 
                           mask_1_39_port, B2 => n340, ZN => n380);
   U459 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => out_mask_39_port);
   U460 : NAND2_X1 port map( A1 => n350, A2 => data_in(14), ZN => n432);
   U461 : NAND2_X1 port map( A1 => n330, A2 => n432, ZN => N59);
   U462 : NAND2_X1 port map( A1 => n350, A2 => data_in(6), ZN => n458);
   U463 : NAND2_X1 port map( A1 => n329, A2 => n458, ZN => N43);
   U464 : INV_X1 port map( A => data_in(30), ZN => n382);
   U465 : OAI21_X1 port map( B1 => n382, B2 => n400, A => n329, ZN => n543);
   U466 : NAND2_X1 port map( A1 => n350, A2 => data_in(22), ZN => n407);
   U467 : NAND2_X1 port map( A1 => n330, A2 => n407, ZN => N83);
   U468 : AOI22_X1 port map( A1 => mask_2_38_port, A2 => n324, B1 => 
                           mask_3_38_port, B2 => n334, ZN => n384);
   U469 : AOI22_X1 port map( A1 => mask_0_38_port, A2 => n317, B1 => 
                           mask_1_38_port, B2 => n340, ZN => n383);
   U470 : NAND2_X1 port map( A1 => n384, A2 => n383, ZN => out_mask_38_port);
   U471 : NAND2_X1 port map( A1 => n350, A2 => data_in(13), ZN => n435);
   U472 : NAND2_X1 port map( A1 => n329, A2 => n435, ZN => N58);
   U473 : NAND2_X1 port map( A1 => n349, A2 => data_in(5), ZN => n463);
   U474 : NAND2_X1 port map( A1 => n330, A2 => n463, ZN => N42);
   U475 : INV_X1 port map( A => data_in(29), ZN => n385);
   U476 : OAI21_X1 port map( B1 => n385, B2 => n400, A => n329, ZN => n544);
   U477 : NAND2_X1 port map( A1 => n349, A2 => data_in(21), ZN => n410);
   U478 : NAND2_X1 port map( A1 => n329, A2 => n410, ZN => N82);
   U479 : AOI22_X1 port map( A1 => mask_2_37_port, A2 => n322, B1 => 
                           mask_3_37_port, B2 => n334, ZN => n387);
   U480 : AOI22_X1 port map( A1 => mask_0_37_port, A2 => n314, B1 => 
                           mask_1_37_port, B2 => n340, ZN => n386);
   U481 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => out_mask_37_port);
   U482 : NAND2_X1 port map( A1 => n349, A2 => data_in(12), ZN => n438);
   U483 : NAND2_X1 port map( A1 => n330, A2 => n438, ZN => N57);
   U484 : NAND2_X1 port map( A1 => n349, A2 => data_in(4), ZN => n468);
   U485 : NAND2_X1 port map( A1 => n329, A2 => n468, ZN => N41);
   U486 : INV_X1 port map( A => data_in(28), ZN => n388);
   U487 : OAI21_X1 port map( B1 => n388, B2 => n400, A => n329, ZN => n545);
   U488 : NAND2_X1 port map( A1 => n349, A2 => data_in(20), ZN => n413);
   U489 : NAND2_X1 port map( A1 => n330, A2 => n413, ZN => N81);
   U490 : AOI22_X1 port map( A1 => mask_2_36_port, A2 => n321, B1 => 
                           mask_3_36_port, B2 => n334, ZN => n390);
   U491 : AOI22_X1 port map( A1 => mask_0_36_port, A2 => n313, B1 => 
                           mask_1_36_port, B2 => n340, ZN => n389);
   U492 : NAND2_X1 port map( A1 => n390, A2 => n389, ZN => out_mask_36_port);
   U493 : NAND2_X1 port map( A1 => n349, A2 => data_in(11), ZN => n441);
   U494 : NAND2_X1 port map( A1 => n330, A2 => n441, ZN => N56);
   U495 : NAND2_X1 port map( A1 => n349, A2 => data_in(3), ZN => n473);
   U496 : NAND2_X1 port map( A1 => n330, A2 => n473, ZN => N40);
   U497 : INV_X1 port map( A => data_in(27), ZN => n391);
   U498 : OAI21_X1 port map( B1 => n391, B2 => n400, A => n329, ZN => n546);
   U499 : NAND2_X1 port map( A1 => n349, A2 => data_in(19), ZN => n416);
   U500 : NAND2_X1 port map( A1 => n330, A2 => n416, ZN => N80);
   U501 : AOI22_X1 port map( A1 => mask_2_35_port, A2 => n322, B1 => 
                           mask_3_35_port, B2 => n334, ZN => n393);
   U502 : AOI22_X1 port map( A1 => mask_0_35_port, A2 => n314, B1 => 
                           mask_1_35_port, B2 => n340, ZN => n392);
   U503 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => out_mask_35_port);
   U504 : NAND2_X1 port map( A1 => n349, A2 => data_in(10), ZN => n444);
   U505 : NAND2_X1 port map( A1 => n330, A2 => n444, ZN => N55);
   U506 : NAND2_X1 port map( A1 => n349, A2 => data_in(2), ZN => n478);
   U507 : NAND2_X1 port map( A1 => n330, A2 => n478, ZN => N39);
   U508 : INV_X1 port map( A => data_in(26), ZN => n394);
   U509 : OAI21_X1 port map( B1 => n394, B2 => n400, A => n329, ZN => n547);
   U510 : NAND2_X1 port map( A1 => n349, A2 => data_in(18), ZN => n419);
   U511 : NAND2_X1 port map( A1 => n330, A2 => n419, ZN => N79);
   U512 : AOI22_X1 port map( A1 => mask_2_34_port, A2 => n319, B1 => 
                           mask_3_34_port, B2 => n334, ZN => n396);
   U513 : AOI22_X1 port map( A1 => mask_0_34_port, A2 => n310, B1 => 
                           mask_1_34_port, B2 => n340, ZN => n395);
   U514 : NAND2_X1 port map( A1 => n396, A2 => n395, ZN => out_mask_34_port);
   U515 : NAND2_X1 port map( A1 => n349, A2 => data_in(9), ZN => n447);
   U516 : NAND2_X1 port map( A1 => n330, A2 => n447, ZN => N54);
   U517 : NAND2_X1 port map( A1 => n349, A2 => data_in(1), ZN => n483);
   U518 : NAND2_X1 port map( A1 => n330, A2 => n483, ZN => N38);
   U519 : INV_X1 port map( A => data_in(25), ZN => n397);
   U520 : OAI21_X1 port map( B1 => n397, B2 => n400, A => n329, ZN => n548);
   U521 : NAND2_X1 port map( A1 => n348, A2 => data_in(17), ZN => n422);
   U522 : NAND2_X1 port map( A1 => n330, A2 => n422, ZN => N78);
   U523 : AOI22_X1 port map( A1 => mask_2_33_port, A2 => n324, B1 => 
                           mask_3_33_port, B2 => n334, ZN => n399);
   U524 : AOI22_X1 port map( A1 => mask_0_33_port, A2 => n316, B1 => 
                           mask_1_33_port, B2 => n340, ZN => n398);
   U525 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => out_mask_33_port);
   U526 : NAND2_X1 port map( A1 => n348, A2 => data_in(8), ZN => n450);
   U527 : NAND2_X1 port map( A1 => n330, A2 => n450, ZN => N53);
   U528 : NAND2_X1 port map( A1 => n348, A2 => data_in(0), ZN => n489);
   U529 : NAND2_X1 port map( A1 => n489, A2 => n329, ZN => N37);
   U530 : INV_X1 port map( A => data_in(24), ZN => n401);
   U531 : OAI21_X1 port map( B1 => n401, B2 => n400, A => n329, ZN => n549);
   U532 : NAND2_X1 port map( A1 => n348, A2 => data_in(16), ZN => n425);
   U533 : NAND2_X1 port map( A1 => n330, A2 => n425, ZN => N77);
   U534 : AOI22_X1 port map( A1 => mask_2_32_port, A2 => n323, B1 => 
                           mask_3_32_port, B2 => n334, ZN => n403);
   U535 : AOI22_X1 port map( A1 => mask_0_32_port, A2 => n315, B1 => 
                           mask_1_32_port, B2 => n340, ZN => n402);
   U536 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => out_mask_32_port);
   U537 : INV_X1 port map( A => n550, ZN => n404);
   U538 : NAND2_X1 port map( A1 => n219_port, A2 => n404, ZN => N116);
   U539 : AOI22_X1 port map( A1 => mask_2_31_port, A2 => n319, B1 => 
                           mask_3_31_port, B2 => n334, ZN => n406);
   U540 : AOI22_X1 port map( A1 => mask_0_31_port, A2 => n311, B1 => 
                           mask_1_31_port, B2 => n340, ZN => n405);
   U541 : NAND2_X1 port map( A1 => data_in(30), A2 => n488, ZN => n457);
   U542 : NAND2_X1 port map( A1 => n457, A2 => n407, ZN => N115);
   U543 : AOI22_X1 port map( A1 => mask_2_30_port, A2 => n325, B1 => 
                           mask_3_30_port, B2 => n334, ZN => n409);
   U544 : AOI22_X1 port map( A1 => mask_0_30_port, A2 => n317, B1 => 
                           mask_1_30_port, B2 => n340, ZN => n408);
   U545 : NAND2_X1 port map( A1 => data_in(29), A2 => n488, ZN => n462);
   U546 : NAND2_X1 port map( A1 => n462, A2 => n410, ZN => N114);
   U547 : AOI22_X1 port map( A1 => mask_2_29_port, A2 => n322, B1 => 
                           mask_3_29_port, B2 => n334, ZN => n412);
   U548 : AOI22_X1 port map( A1 => mask_0_29_port, A2 => n314, B1 => 
                           mask_1_29_port, B2 => n340, ZN => n411);
   U549 : NAND2_X1 port map( A1 => data_in(28), A2 => n488, ZN => n467);
   U550 : NAND2_X1 port map( A1 => n467, A2 => n413, ZN => N113);
   U551 : AOI22_X1 port map( A1 => mask_2_28_port, A2 => n320, B1 => 
                           mask_3_28_port, B2 => n334, ZN => n415);
   U552 : AOI22_X1 port map( A1 => mask_0_28_port, A2 => n312, B1 => 
                           mask_1_28_port, B2 => n340, ZN => n414);
   U553 : NAND2_X1 port map( A1 => data_in(27), A2 => n488, ZN => n472);
   U554 : NAND2_X1 port map( A1 => n472, A2 => n416, ZN => N112);
   U555 : AOI22_X1 port map( A1 => mask_2_27_port, A2 => n1, B1 => 
                           mask_3_27_port, B2 => n335, ZN => n418);
   U556 : AOI22_X1 port map( A1 => mask_0_27_port, A2 => n2, B1 => 
                           mask_1_27_port, B2 => n341, ZN => n417);
   U557 : NAND2_X1 port map( A1 => data_in(26), A2 => n488, ZN => n477);
   U558 : NAND2_X1 port map( A1 => n477, A2 => n419, ZN => N111);
   U559 : AOI22_X1 port map( A1 => mask_2_26_port, A2 => n321, B1 => 
                           mask_3_26_port, B2 => n335, ZN => n421);
   U560 : AOI22_X1 port map( A1 => mask_0_26_port, A2 => n313, B1 => 
                           mask_1_26_port, B2 => n341, ZN => n420);
   U561 : NAND2_X1 port map( A1 => data_in(25), A2 => n488, ZN => n482);
   U562 : NAND2_X1 port map( A1 => n482, A2 => n422, ZN => N110);
   U563 : AOI22_X1 port map( A1 => mask_2_25_port, A2 => n325, B1 => 
                           mask_3_25_port, B2 => n335, ZN => n424);
   U564 : AOI22_X1 port map( A1 => mask_0_25_port, A2 => n317, B1 => 
                           mask_1_25_port, B2 => n341, ZN => n423);
   U565 : NAND2_X1 port map( A1 => data_in(24), A2 => n488, ZN => n487);
   U566 : NAND2_X1 port map( A1 => n487, A2 => n425, ZN => N109);
   U567 : AOI22_X1 port map( A1 => mask_2_24_port, A2 => n324, B1 => 
                           mask_3_24_port, B2 => n335, ZN => n427);
   U568 : AOI22_X1 port map( A1 => mask_0_24_port, A2 => n316, B1 => 
                           mask_1_24_port, B2 => n341, ZN => n426);
   U569 : NAND2_X1 port map( A1 => data_in(23), A2 => n488, ZN => n454);
   U570 : NAND2_X1 port map( A1 => n454, A2 => n428, ZN => N108);
   U571 : INV_X1 port map( A => n541, ZN => n429);
   U572 : NAND2_X1 port map( A1 => n219_port, A2 => n429, ZN => N76);
   U573 : AOI22_X1 port map( A1 => mask_2_23_port, A2 => n1, B1 => 
                           mask_3_23_port, B2 => n335, ZN => n431);
   U574 : AOI22_X1 port map( A1 => mask_0_23_port, A2 => n2, B1 => 
                           mask_1_23_port, B2 => n341, ZN => n430);
   U575 : NAND2_X1 port map( A1 => data_in(22), A2 => n488, ZN => n459);
   U576 : NAND2_X1 port map( A1 => n459, A2 => n432, ZN => n551);
   U577 : NAND2_X1 port map( A1 => n457, A2 => n458, ZN => N75);
   U578 : AOI22_X1 port map( A1 => mask_2_22_port, A2 => n324, B1 => 
                           mask_3_22_port, B2 => n335, ZN => n434);
   U579 : AOI22_X1 port map( A1 => mask_0_22_port, A2 => n316, B1 => 
                           mask_1_22_port, B2 => n341, ZN => n433);
   U580 : NAND2_X1 port map( A1 => data_in(21), A2 => n488, ZN => n464);
   U581 : NAND2_X1 port map( A1 => n464, A2 => n435, ZN => n552);
   U582 : NAND2_X1 port map( A1 => n462, A2 => n463, ZN => N74);
   U583 : AOI22_X1 port map( A1 => mask_2_21_port, A2 => n323, B1 => 
                           mask_3_21_port, B2 => n335, ZN => n437);
   U584 : AOI22_X1 port map( A1 => mask_0_21_port, A2 => n315, B1 => 
                           mask_1_21_port, B2 => n341, ZN => n436);
   U585 : NAND2_X1 port map( A1 => data_in(20), A2 => n488, ZN => n469);
   U586 : NAND2_X1 port map( A1 => n469, A2 => n438, ZN => n553);
   U587 : NAND2_X1 port map( A1 => n467, A2 => n468, ZN => N73);
   U588 : AOI22_X1 port map( A1 => mask_2_20_port, A2 => n321, B1 => 
                           mask_3_20_port, B2 => n335, ZN => n440);
   U589 : AOI22_X1 port map( A1 => mask_0_20_port, A2 => n313, B1 => 
                           mask_1_20_port, B2 => n341, ZN => n439);
   U590 : NAND2_X1 port map( A1 => data_in(19), A2 => n488, ZN => n474);
   U591 : NAND2_X1 port map( A1 => n474, A2 => n441, ZN => n554);
   U592 : NAND2_X1 port map( A1 => n472, A2 => n473, ZN => N72);
   U593 : AOI22_X1 port map( A1 => mask_2_19_port, A2 => n322, B1 => 
                           mask_3_19_port, B2 => n335, ZN => n443);
   U594 : AOI22_X1 port map( A1 => mask_0_19_port, A2 => n314, B1 => 
                           mask_1_19_port, B2 => n341, ZN => n442);
   U595 : NAND2_X1 port map( A1 => data_in(18), A2 => n488, ZN => n479);
   U596 : NAND2_X1 port map( A1 => n479, A2 => n444, ZN => n555);
   U597 : NAND2_X1 port map( A1 => n477, A2 => n478, ZN => N71);
   U598 : AOI22_X1 port map( A1 => mask_2_18_port, A2 => n321, B1 => 
                           mask_3_18_port, B2 => n335, ZN => n446);
   U599 : AOI22_X1 port map( A1 => mask_0_18_port, A2 => n313, B1 => 
                           mask_1_18_port, B2 => n341, ZN => n445);
   U600 : NAND2_X1 port map( A1 => data_in(17), A2 => n488, ZN => n484);
   U601 : NAND2_X1 port map( A1 => n484, A2 => n447, ZN => n556);
   U602 : NAND2_X1 port map( A1 => n482, A2 => n483, ZN => N70);
   U603 : AOI22_X1 port map( A1 => mask_2_17_port, A2 => n320, B1 => 
                           mask_3_17_port, B2 => n335, ZN => n449);
   U604 : AOI22_X1 port map( A1 => mask_0_17_port, A2 => n312, B1 => 
                           mask_1_17_port, B2 => n341, ZN => n448);
   U605 : NAND2_X1 port map( A1 => data_in(16), A2 => n488, ZN => n490);
   U606 : NAND2_X1 port map( A1 => n490, A2 => n450, ZN => n557);
   U607 : NAND2_X1 port map( A1 => n487, A2 => n489, ZN => N69);
   U608 : AOI22_X1 port map( A1 => mask_2_16_port, A2 => n1, B1 => 
                           mask_3_16_port, B2 => n335, ZN => n452);
   U609 : AOI22_X1 port map( A1 => mask_0_16_port, A2 => n2, B1 => 
                           mask_1_16_port, B2 => n341, ZN => n451);
   U610 : NAND2_X1 port map( A1 => n219_port, A2 => n329, ZN => N35);
   U611 : NAND2_X1 port map( A1 => data_in(15), A2 => n488, ZN => n494);
   U612 : NAND2_X1 port map( A1 => n494, A2 => n453, ZN => n558);
   U613 : INV_X1 port map( A => n454, ZN => n533);
   U614 : AOI22_X1 port map( A1 => mask_2_15_port, A2 => n324, B1 => 
                           mask_3_15_port, B2 => n336, ZN => n456);
   U615 : AOI22_X1 port map( A1 => mask_0_15_port, A2 => n317, B1 => 
                           mask_1_15_port, B2 => n342, ZN => n455);
   U616 : INV_X1 port map( A => n457, ZN => n540);
   U617 : NAND2_X1 port map( A1 => data_in(14), A2 => n488, ZN => n498);
   U618 : NAND2_X1 port map( A1 => n498, A2 => n458, ZN => N99);
   U619 : INV_X1 port map( A => n459, ZN => n532);
   U620 : AOI22_X1 port map( A1 => mask_2_14_port, A2 => n319, B1 => 
                           mask_3_14_port, B2 => n336, ZN => n461);
   U621 : AOI22_X1 port map( A1 => mask_0_14_port, A2 => n311, B1 => 
                           mask_1_14_port, B2 => n342, ZN => n460);
   U622 : INV_X1 port map( A => n462, ZN => n539);
   U623 : NAND2_X1 port map( A1 => data_in(13), A2 => n488, ZN => n502);
   U624 : NAND2_X1 port map( A1 => n502, A2 => n463, ZN => N98);
   U625 : INV_X1 port map( A => n464, ZN => n531);
   U626 : AOI22_X1 port map( A1 => mask_2_13_port, A2 => n318, B1 => 
                           mask_3_13_port, B2 => n336, ZN => n466);
   U627 : AOI22_X1 port map( A1 => mask_0_13_port, A2 => n310, B1 => 
                           mask_1_13_port, B2 => n342, ZN => n465);
   U628 : INV_X1 port map( A => n467, ZN => n538);
   U629 : NAND2_X1 port map( A1 => data_in(12), A2 => n488, ZN => n506);
   U630 : NAND2_X1 port map( A1 => n506, A2 => n468, ZN => N97);
   U631 : INV_X1 port map( A => n469, ZN => n530);
   U632 : AOI22_X1 port map( A1 => mask_2_12_port, A2 => n325, B1 => 
                           mask_3_12_port, B2 => n336, ZN => n471);
   U633 : AOI22_X1 port map( A1 => mask_0_12_port, A2 => n317, B1 => 
                           mask_1_12_port, B2 => n342, ZN => n470);
   U634 : INV_X1 port map( A => n472, ZN => n537);
   U635 : NAND2_X1 port map( A1 => data_in(11), A2 => n488, ZN => n510);
   U636 : NAND2_X1 port map( A1 => n510, A2 => n473, ZN => N96);
   U637 : INV_X1 port map( A => n474, ZN => n529);
   U638 : AOI22_X1 port map( A1 => mask_2_11_port, A2 => n320, B1 => 
                           mask_3_11_port, B2 => n336, ZN => n476);
   U639 : AOI22_X1 port map( A1 => mask_0_11_port, A2 => n312, B1 => 
                           mask_1_11_port, B2 => n342, ZN => n475);
   U640 : INV_X1 port map( A => n477, ZN => n536);
   U641 : NAND2_X1 port map( A1 => data_in(10), A2 => n488, ZN => n514);
   U642 : NAND2_X1 port map( A1 => n514, A2 => n478, ZN => N95);
   U643 : INV_X1 port map( A => n479, ZN => n528);
   U644 : AOI22_X1 port map( A1 => mask_2_10_port, A2 => n323, B1 => 
                           mask_3_10_port, B2 => n336, ZN => n481);
   U645 : AOI22_X1 port map( A1 => mask_0_10_port, A2 => n315, B1 => 
                           mask_1_10_port, B2 => n342, ZN => n480);
   U646 : INV_X1 port map( A => n482, ZN => n535);
   U647 : NAND2_X1 port map( A1 => data_in(9), A2 => n488, ZN => n518);
   U648 : NAND2_X1 port map( A1 => n518, A2 => n483, ZN => N94);
   U649 : INV_X1 port map( A => n484, ZN => n527);
   U650 : AOI22_X1 port map( A1 => mask_2_9_port, A2 => n325, B1 => 
                           mask_3_9_port, B2 => n336, ZN => n486);
   U651 : AOI22_X1 port map( A1 => mask_0_9_port, A2 => n317, B1 => 
                           mask_1_9_port, B2 => n342, ZN => n485);
   U652 : INV_X1 port map( A => n487, ZN => n534);
   U653 : NAND2_X1 port map( A1 => data_in(8), A2 => n488, ZN => n522);
   U654 : NAND2_X1 port map( A1 => n522, A2 => n489, ZN => N93);
   U655 : INV_X1 port map( A => n490, ZN => n526);
   U656 : AOI22_X1 port map( A1 => mask_2_8_port, A2 => n1, B1 => mask_3_8_port
                           , B2 => n336, ZN => n492);
   U657 : AOI22_X1 port map( A1 => mask_0_8_port, A2 => n2, B1 => mask_1_8_port
                           , B2 => n342, ZN => n491);
   U658 : INV_X1 port map( A => data_in(7), ZN => n493);
   U659 : NOR2_X1 port map( A1 => n229, A2 => n493, ZN => N92);
   U660 : INV_X1 port map( A => n494, ZN => N68);
   U661 : AOI22_X1 port map( A1 => mask_2_7_port, A2 => n320, B1 => 
                           mask_3_7_port, B2 => n336, ZN => n496);
   U662 : AOI22_X1 port map( A1 => mask_0_7_port, A2 => n312, B1 => 
                           mask_1_7_port, B2 => n342, ZN => n495);
   U663 : INV_X1 port map( A => data_in(6), ZN => n497);
   U664 : NOR2_X1 port map( A1 => n229, A2 => n497, ZN => N91);
   U665 : INV_X1 port map( A => n498, ZN => n559);
   U666 : AOI22_X1 port map( A1 => mask_2_6_port, A2 => n323, B1 => 
                           mask_3_6_port, B2 => n336, ZN => n500);
   U667 : AOI22_X1 port map( A1 => mask_0_6_port, A2 => n315, B1 => 
                           mask_1_6_port, B2 => n342, ZN => n499);
   U668 : INV_X1 port map( A => data_in(5), ZN => n501);
   U669 : NOR2_X1 port map( A1 => n229, A2 => n501, ZN => N90);
   U670 : INV_X1 port map( A => n502, ZN => n560);
   U671 : AOI22_X1 port map( A1 => mask_2_5_port, A2 => n323, B1 => 
                           mask_3_5_port, B2 => n336, ZN => n504);
   U672 : AOI22_X1 port map( A1 => mask_0_5_port, A2 => n315, B1 => 
                           mask_1_5_port, B2 => n342, ZN => n503);
   U673 : NAND2_X1 port map( A1 => n504, A2 => n503, ZN => out_mask_5_port);
   U674 : INV_X1 port map( A => data_in(4), ZN => n505);
   U675 : NOR2_X1 port map( A1 => n229, A2 => n505, ZN => N89);
   U676 : INV_X1 port map( A => n506, ZN => n561);
   U677 : AOI22_X1 port map( A1 => mask_2_4_port, A2 => n325, B1 => 
                           mask_3_4_port, B2 => n336, ZN => n508);
   U678 : AOI22_X1 port map( A1 => mask_0_4_port, A2 => n316, B1 => 
                           mask_1_4_port, B2 => n342, ZN => n507);
   U679 : NAND2_X1 port map( A1 => n508, A2 => n507, ZN => out_mask_4_port);
   U680 : INV_X1 port map( A => data_in(3), ZN => n509);
   U681 : NOR2_X1 port map( A1 => n229, A2 => n509, ZN => N88);
   U682 : INV_X1 port map( A => n510, ZN => n562);
   U683 : AOI22_X1 port map( A1 => mask_2_3_port, A2 => n325, B1 => 
                           mask_3_3_port, B2 => n337, ZN => n512);
   U684 : AOI22_X1 port map( A1 => mask_0_3_port, A2 => n316, B1 => 
                           mask_1_3_port, B2 => n343, ZN => n511);
   U685 : NAND2_X1 port map( A1 => n512, A2 => n511, ZN => out_mask_3_port);
   U686 : INV_X1 port map( A => data_in(2), ZN => n513);
   U687 : NOR2_X1 port map( A1 => n229, A2 => n513, ZN => N87);
   U688 : INV_X1 port map( A => n514, ZN => n563);
   U689 : AOI22_X1 port map( A1 => mask_2_2_port, A2 => n1, B1 => mask_3_2_port
                           , B2 => n337, ZN => n516);
   U690 : AOI22_X1 port map( A1 => mask_0_2_port, A2 => n2, B1 => mask_1_2_port
                           , B2 => n343, ZN => n515);
   U691 : NAND2_X1 port map( A1 => n516, A2 => n515, ZN => out_mask_2_port);
   U692 : INV_X1 port map( A => data_in(1), ZN => n517);
   U693 : NOR2_X1 port map( A1 => n229, A2 => n517, ZN => N86);
   U694 : INV_X1 port map( A => n518, ZN => n564);
   U695 : AOI22_X1 port map( A1 => mask_2_1_port, A2 => n318, B1 => 
                           mask_3_1_port, B2 => n337, ZN => n520);
   U696 : AOI22_X1 port map( A1 => mask_0_1_port, A2 => n311, B1 => 
                           mask_1_1_port, B2 => n343, ZN => n519);
   U697 : NAND2_X1 port map( A1 => n520, A2 => n519, ZN => out_mask_1_port);
   U698 : INV_X1 port map( A => data_in(0), ZN => n521);
   U699 : NOR2_X1 port map( A1 => n229, A2 => n521, ZN => N85);
   U700 : INV_X1 port map( A => n522, ZN => n565);
   U701 : AOI22_X1 port map( A1 => mask_2_0_port, A2 => n320, B1 => 
                           mask_3_0_port, B2 => n337, ZN => n524);
   U702 : AOI22_X1 port map( A1 => mask_0_0_port, A2 => n312, B1 => 
                           mask_1_0_port, B2 => n343, ZN => n523);
   U703 : NAND2_X1 port map( A1 => n524, A2 => n523, ZN => out_mask_0_port);
   U704 : MUX2_X1 port map( A => N190, B => N158, S => n348, Z => data_out(0));
   U705 : MUX2_X1 port map( A => N191, B => N159, S => n348, Z => data_out(1));
   U706 : MUX2_X1 port map( A => N192, B => N160, S => n348, Z => data_out(2));
   U707 : MUX2_X1 port map( A => N193, B => N161, S => n348, Z => data_out(3));
   U708 : MUX2_X1 port map( A => N194, B => N162, S => n348, Z => data_out(4));
   U709 : MUX2_X1 port map( A => N195, B => N163, S => n348, Z => data_out(5));
   U710 : MUX2_X1 port map( A => N196, B => N164, S => n348, Z => data_out(6));
   U711 : MUX2_X1 port map( A => N197, B => N165, S => n348, Z => data_out(7));
   U712 : MUX2_X1 port map( A => N198, B => N166, S => n347, Z => data_out(8));
   U713 : MUX2_X1 port map( A => N199, B => N167, S => n347, Z => data_out(9));
   U714 : MUX2_X1 port map( A => N200, B => N168, S => n347, Z => data_out(10))
                           ;
   U715 : MUX2_X1 port map( A => N201, B => N169, S => n347, Z => data_out(11))
                           ;
   U716 : MUX2_X1 port map( A => N202, B => N170, S => n347, Z => data_out(12))
                           ;
   U717 : MUX2_X1 port map( A => N203, B => N171, S => n347, Z => data_out(13))
                           ;
   U718 : MUX2_X1 port map( A => N204, B => N172, S => n347, Z => data_out(14))
                           ;
   U719 : MUX2_X1 port map( A => N205, B => N173, S => n347, Z => data_out(15))
                           ;
   U720 : MUX2_X1 port map( A => N206, B => N174, S => n347, Z => data_out(16))
                           ;
   U721 : MUX2_X1 port map( A => N207, B => N175, S => n347, Z => data_out(17))
                           ;
   U722 : MUX2_X1 port map( A => N208, B => N176, S => n347, Z => data_out(18))
                           ;
   U723 : MUX2_X1 port map( A => N209, B => N177, S => n347, Z => data_out(19))
                           ;
   U724 : MUX2_X1 port map( A => N210, B => N178, S => n346, Z => data_out(20))
                           ;
   U725 : MUX2_X1 port map( A => N211, B => N179, S => n346, Z => data_out(21))
                           ;
   U726 : MUX2_X1 port map( A => N212, B => N180, S => n346, Z => data_out(22))
                           ;
   U727 : MUX2_X1 port map( A => N213, B => N181, S => n346, Z => data_out(23))
                           ;
   U728 : MUX2_X1 port map( A => N214, B => N182, S => n346, Z => data_out(24))
                           ;
   U729 : MUX2_X1 port map( A => N215, B => N183, S => n346, Z => data_out(25))
                           ;
   U730 : MUX2_X1 port map( A => N216, B => N184, S => n346, Z => data_out(26))
                           ;
   U731 : MUX2_X1 port map( A => N217, B => N185, S => n346, Z => data_out(27))
                           ;
   U732 : MUX2_X1 port map( A => N218, B => N186, S => n346, Z => data_out(28))
                           ;
   U733 : MUX2_X1 port map( A => N219, B => N187, S => n346, Z => data_out(29))
                           ;
   U734 : MUX2_X1 port map( A => N220, B => N188, S => n346, Z => data_out(30))
                           ;
   U735 : MUX2_X1 port map( A => N221, B => N189, S => n346, Z => data_out(31))
                           ;

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal C_internal, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, carry_1_port, carry_0_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38 : std_logic;

begin
   
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => n30, 
                           B(30) => n32, B(29) => n31, B(28) => n29, B(27) => 
                           n28, B(26) => n27, B(25) => n25, B(24) => n26, B(23)
                           => n12, B(22) => n23, B(21) => n11, B(20) => n22, 
                           B(19) => n8, B(18) => n20, B(17) => n15, B(16) => 
                           n10, B(15) => n17, B(14) => n13, B(13) => n24, B(12)
                           => n14, B(11) => n18, B(10) => n19, B(9) => n21, 
                           B(8) => n9, B(7) => n7, B(6) => n16, B(5) => n6, 
                           B(4) => n3, B(3) => n1, B(2) => n5, B(1) => n4, B(0)
                           => n2, Cin => C_internal, Co(8) => Cout, Co(7) => 
                           carry_7_port, Co(6) => carry_6_port, Co(5) => 
                           carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => n30, B(30) => n32, 
                           B(29) => n31, B(28) => n29, B(27) => n28, B(26) => 
                           n27, B(25) => n25, B(24) => n26, B(23) => n12, B(22)
                           => n23, B(21) => n11, B(20) => n22, B(19) => n8, 
                           B(18) => n20, B(17) => n15, B(16) => n10, B(15) => 
                           n17, B(14) => n13, B(13) => n24, B(12) => n14, B(11)
                           => n18, B(10) => n19, B(9) => n21, B(8) => n9, B(7) 
                           => n7, B(6) => n16, B(5) => n6, B(4) => n3, B(3) => 
                           n1, B(2) => n5, B(1) => n4, B(0) => n2, Ci(7) => 
                           carry_7_port, Ci(6) => carry_6_port, Ci(5) => 
                           carry_5_port, Ci(4) => carry_4_port, Ci(3) => 
                           carry_3_port, Ci(2) => carry_2_port, Ci(1) => 
                           carry_1_port, Ci(0) => carry_0_port, S(31) => S(31),
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U4 : XNOR2_X1 port map( A => n34, B => B(3), ZN => n1);
   U5 : BUF_X1 port map( A => n38, Z => n37);
   U6 : CLKBUF_X1 port map( A => n38, Z => n36);
   U7 : CLKBUF_X1 port map( A => n38, Z => n35);
   U8 : CLKBUF_X1 port map( A => n38, Z => n33);
   U9 : BUF_X1 port map( A => n38, Z => n34);
   U10 : XNOR2_X1 port map( A => n38, B => B(0), ZN => n2);
   U11 : XNOR2_X1 port map( A => n37, B => B(4), ZN => n3);
   U12 : XNOR2_X1 port map( A => n36, B => B(1), ZN => n4);
   U13 : XNOR2_X1 port map( A => n35, B => B(2), ZN => n5);
   U14 : XNOR2_X1 port map( A => n36, B => B(5), ZN => n6);
   U15 : XNOR2_X1 port map( A => n33, B => B(7), ZN => n7);
   U16 : XNOR2_X1 port map( A => n37, B => B(19), ZN => n8);
   U17 : XNOR2_X1 port map( A => n37, B => B(8), ZN => n9);
   U18 : XNOR2_X1 port map( A => n36, B => B(16), ZN => n10);
   U19 : XNOR2_X1 port map( A => n33, B => B(21), ZN => n11);
   U20 : XNOR2_X1 port map( A => n35, B => B(23), ZN => n12);
   U21 : XNOR2_X1 port map( A => n34, B => B(14), ZN => n13);
   U22 : XNOR2_X1 port map( A => n33, B => B(12), ZN => n14);
   U23 : XNOR2_X1 port map( A => n34, B => B(17), ZN => n15);
   U24 : XNOR2_X1 port map( A => n35, B => B(6), ZN => n16);
   U25 : XNOR2_X1 port map( A => n36, B => B(15), ZN => n17);
   U26 : XNOR2_X1 port map( A => n34, B => B(11), ZN => n18);
   U27 : XNOR2_X1 port map( A => n33, B => B(10), ZN => n19);
   U28 : XNOR2_X1 port map( A => n36, B => B(18), ZN => n20);
   U29 : XNOR2_X1 port map( A => n35, B => B(9), ZN => n21);
   U30 : XNOR2_X1 port map( A => n35, B => B(20), ZN => n22);
   U31 : XNOR2_X1 port map( A => n37, B => B(22), ZN => n23);
   U32 : XNOR2_X1 port map( A => n37, B => B(13), ZN => n24);
   U33 : XNOR2_X1 port map( A => n33, B => B(25), ZN => n25);
   U34 : XNOR2_X1 port map( A => n36, B => B(24), ZN => n26);
   U35 : XNOR2_X1 port map( A => n35, B => B(26), ZN => n27);
   U36 : XNOR2_X1 port map( A => n34, B => B(27), ZN => n28);
   U37 : XNOR2_X1 port map( A => n37, B => B(28), ZN => n29);
   U38 : XNOR2_X1 port map( A => n34, B => B(31), ZN => n30);
   U39 : XNOR2_X1 port map( A => n33, B => B(29), ZN => n31);
   U40 : XNOR2_X1 port map( A => n36, B => B(30), ZN => n32);
   U41 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);
   U42 : INV_X1 port map( A => ADD_SUB, ZN => n38);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_0;

architecture SYN_Behavioral of AND2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_NBIT32_NREG32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_NBIT32_NREG32;

architecture SYN_BEHAVIORAL of RF_NBIT32_NREG32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N128, N129, N130, N131, N132, 
      N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, 
      N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, 
      N157, N158, N159, N193, N194, N195, N196, N197, N198, N199, N200, N201, 
      N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, 
      N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, 
      N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, 
      N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, 
      N250, N251, N252, N253, N254, N255, N256, N259, N260, N261, N262, N263, 
      N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, 
      N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, 
      N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, 
      N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, 
      N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, 
      N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, 
      N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, 
      N348, N349, N350, N351, N352, N353, n1, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n2, n3, 
      n4, n5, n6, n7, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128_port, n129_port, n130_port, 
      n131_port, n132_port, n133_port, n134_port, n135_port, n136_port, 
      n137_port, n138_port, n139_port, n140_port, n141_port, n142_port, 
      n143_port, n144_port, n145_port, n146_port, n147_port, n148_port, 
      n149_port, n150_port, n151_port, n152_port, n153_port, n154_port, 
      n155_port, n156_port, n157_port, n158_port, n159_port, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193_port, n194_port, n195_port, 
      n196_port, n197_port, n198_port, n199_port, n200_port, n201_port, 
      n202_port, n203_port, n204_port, n205_port, n206_port, n207_port, 
      n208_port, n209_port, n210_port, n211_port, n212_port, n213_port, 
      n214_port, n215_port, n216_port, n217_port, n218_port, n219_port, 
      n220_port, n221_port, n222_port, n223_port, n224_port, n225_port, 
      n226_port, n227_port, n228_port, n229_port, n230_port, n231_port, 
      n232_port, n233_port, n234_port, n235_port, n236_port, n237_port, 
      n238_port, n239_port, n240_port, n241_port, n242_port, n243_port, 
      n244_port, n245_port, n246_port, n247_port, n248_port, n249_port, 
      n250_port, n251_port, n252_port, n253_port, n254_port, n255_port, 
      n256_port, n257, n258, n259_port, n260_port, n261_port, n262_port, 
      n263_port, n264_port, n265_port, n266_port, n267_port, n268_port, 
      n269_port, n270_port, n271_port, n272_port, n273_port, n274_port, 
      n275_port, n276_port, n277_port, n278_port, n279_port, n280_port, 
      n281_port, n282_port, n283_port, n284_port, n285_port, n286_port, 
      n287_port, n288_port, n289_port, n290_port, n291_port, n292_port, 
      n293_port, n294_port, n295_port, n296_port, n297_port, n298_port, 
      n299_port, n300_port, n301_port, n302_port, n303_port, n304_port, 
      n305_port, n306_port, n307_port, n308_port, n309_port, n310_port, 
      n311_port, n312_port, n313_port, n314_port, n315_port, n316_port, 
      n317_port, n318_port, n319_port, n320_port, n321_port, n322_port, 
      n323_port, n324_port, n325_port, n326_port, n327_port, n328_port, 
      n329_port, n330_port, n331_port, n332_port, n333_port, n334_port, 
      n335_port, n336_port, n337_port, n338_port, n339_port, n340_port, 
      n341_port, n342_port, n343_port, n344_port, n345_port, n346_port, 
      n347_port, n348_port, n349_port, n350_port, n351_port, n352_port, 
      n353_port, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
      n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
      n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
      n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
      n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
      n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796 : std_logic;

begin
   
   OUT1_reg_31_inst : DLH_X1 port map( G => CLK, D => N256, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => CLK, D => N255, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => CLK, D => N254, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => CLK, D => N253, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => CLK, D => N252, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => CLK, D => N251, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => CLK, D => N250, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => CLK, D => N249, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => CLK, D => N248, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => CLK, D => N247, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => CLK, D => N246, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => CLK, D => N245, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => CLK, D => N244, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => CLK, D => N243, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => CLK, D => N242, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => CLK, D => N241, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => CLK, D => N240, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => CLK, D => N239, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => CLK, D => N238, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => CLK, D => N237, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => CLK, D => N236, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => CLK, D => N235, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => CLK, D => N234, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => CLK, D => N233, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => CLK, D => N232, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => CLK, D => N231, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => CLK, D => N230, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => CLK, D => N229, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => CLK, D => N228, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => CLK, D => N227, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => CLK, D => N226, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => CLK, D => N225, Q => OUT1(0));
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => N353, D => n1698, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => N353, D => n1701, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => N353, D => n1704, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => N353, D => n1707, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N353, D => n1710, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => N353, D => n1713, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => N353, D => n1716, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => N353, D => n1719, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => N353, D => n1723, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => N353, D => n1727, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => N353, D => n1731, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => N353, D => n1735, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => N353, D => n1739, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => N353, D => n1743, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => N353, D => n1747, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N353, D => n1751, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => N353, D => n1755, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N353, D => n1759, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N353, D => n1763, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => N353, D => n1767, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => N353, D => n1771, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => N353, D => n1775, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => N353, D => n1779, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => N353, D => n1783, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => N352, D => n1698, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => N352, D => n1701, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => N352, D => n1704, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => N352, D => n1707, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => N352, D => n1710, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => N352, D => n1713, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => N352, D => n1716, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => N352, D => n1719, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => N352, D => n1723, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => N352, D => n1727, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => N352, D => n1731, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => N352, D => n1735, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => N352, D => n1739, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => N352, D => n1743, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N352, D => n1747, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => N352, D => n1751, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N352, D => n1755, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N352, D => n1759, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N352, D => n1763, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => N352, D => n1767, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => N352, D => n1771, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => N352, D => n1775, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => N352, D => n1779, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => N352, D => n1783, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => N351, D => n1698, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => N351, D => n1701, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => N351, D => n1704, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => N351, D => n1707, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => N351, D => n1710, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => N351, D => n1713, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => N351, D => n1716, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => N351, D => n1719, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => N351, D => n1723, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => N351, D => n1727, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => N351, D => n1731, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => N351, D => n1735, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => N351, D => n1739, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => N351, D => n1743, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N351, D => n1747, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => N351, D => n1751, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N351, D => n1755, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N351, D => n1759, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N351, D => n1763, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => N351, D => n1767, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => N351, D => n1771, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => N351, D => n1775, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => N351, D => n1779, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => N351, D => n1783, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => N350, D => n1698, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => N350, D => n1701, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => N350, D => n1704, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => N350, D => n1707, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => N350, D => n1710, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => N350, D => n1713, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => N350, D => n1716, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => N350, D => n1719, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => N350, D => n1723, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => N350, D => n1727, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => N350, D => n1731, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => N350, D => n1735, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => N350, D => n1739, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => N350, D => n1743, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N350, D => n1747, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => N350, D => n1751, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N350, D => n1755, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N350, D => n1759, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N350, D => n1763, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => N350, D => n1767, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => N350, D => n1771, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => N350, D => n1775, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => N350, D => n1779, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => N350, D => n1783, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => N349, D => n1698, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => N349, D => n1701, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => N349, D => n1704, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => N349, D => n1707, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => N349, D => n1710, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => N349, D => n1713, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => N349, D => n1716, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => N349, D => n1719, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => N349, D => n1723, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => N349, D => n1727, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => N349, D => n1731, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => N349, D => n1735, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => N349, D => n1739, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => N349, D => n1743, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N349, D => n1747, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => N349, D => n1751, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N349, D => n1755, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N349, D => n1759, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N349, D => n1763, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => N349, D => n1767, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => N349, D => n1771, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => N349, D => n1775, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => N349, D => n1779, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => N349, D => n1783, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => N348, D => n1698, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => N348, D => n1701, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => N348, D => n1704, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => N348, D => n1707, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => N348, D => n1710, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => N348, D => n1713, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => N348, D => n1716, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => N348, D => n1719, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => N348, D => n1723, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => N348, D => n1727, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => N348, D => n1731, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => N348, D => n1735, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => N348, D => n1739, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => N348, D => n1743, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N348, D => n1747, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => N348, D => n1751, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N348, D => n1755, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N348, D => n1759, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N348, D => n1763, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => N348, D => n1767, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => N348, D => n1771, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => N348, D => n1775, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => N348, D => n1779, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => N348, D => n1783, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => N347, D => n1698, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => N347, D => n1701, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => N347, D => n1704, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => N347, D => n1707, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => N347, D => n1710, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => N347, D => n1713, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => N347, D => n1716, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => N347, D => n1719, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => N347, D => n1723, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => N347, D => n1727, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => N347, D => n1731, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => N347, D => n1735, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => N347, D => n1739, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => N347, D => n1743, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N347, D => n1747, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => N347, D => n1751, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N347, D => n1755, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N347, D => n1759, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N347, D => n1763, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => N347, D => n1767, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => N347, D => n1771, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => N347, D => n1775, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => N347, D => n1779, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => N347, D => n1783, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => N346, D => n1698, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => N346, D => n1701, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => N346, D => n1704, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => N346, D => n1707, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => N346, D => n1710, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => N346, D => n1713, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => N346, D => n1716, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => N346, D => n1719, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => N346, D => n1723, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => N346, D => n1727, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => N346, D => n1731, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => N346, D => n1735, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => N346, D => n1739, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => N346, D => n1743, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => N346, D => n1747, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => N346, D => n1751, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N346, D => n1755, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N346, D => n1759, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N346, D => n1763, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => N346, D => n1767, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => N346, D => n1771, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => N346, D => n1775, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => N346, D => n1779, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N346, D => n1783, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => N345, D => n1698, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => N345, D => n1701, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => N345, D => n1704, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => N345, D => n1707, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => N345, D => n1710, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => N345, D => n1713, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => N345, D => n1716, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => N345, D => n1719, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => N345, D => n1723, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => N345, D => n1727, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => N345, D => n1731, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => N345, D => n1735, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => N345, D => n1739, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => N345, D => n1743, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N345, D => n1747, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => N345, D => n1751, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N345, D => n1755, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N345, D => n1759, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N345, D => n1763, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => N345, D => n1767, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => N345, D => n1771, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => N345, D => n1775, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => N345, D => n1779, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => N345, D => n1783, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => N344, D => n1698, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => N344, D => n1701, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => N344, D => n1704, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => N344, D => n1707, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => N344, D => n1710, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => N344, D => n1713, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => N344, D => n1716, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => N344, D => n1719, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => N344, D => n1723, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => N344, D => n1727, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => N344, D => n1731, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => N344, D => n1735, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => N344, D => n1739, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N344, D => n1743, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => N344, D => n1747, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N344, D => n1751, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => N344, D => n1755, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => N344, D => n1759, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N344, D => n1763, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => N344, D => n1767, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => N344, D => n1771, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => N344, D => n1775, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => N344, D => n1779, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N344, D => n1783, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => N343, D => n1698, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => N343, D => n1701, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => N343, D => n1704, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => N343, D => n1707, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => N343, D => n1710, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => N343, D => n1713, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => N343, D => n1716, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => N343, D => n1719, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => N343, D => n1723, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => N343, D => n1727, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => N343, D => n1731, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => N343, D => n1735, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => N343, D => n1739, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => N343, D => n1743, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N343, D => n1747, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => N343, D => n1751, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N343, D => n1755, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N343, D => n1759, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N343, D => n1763, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => N343, D => n1767, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => N343, D => n1771, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => N343, D => n1775, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => N343, D => n1779, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => N343, D => n1783, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => N342, D => n1699, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => N342, D => n1702, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => N342, D => n1705, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => N342, D => n1708, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => N342, D => n1711, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => N342, D => n1714, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => N342, D => n1717, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => N342, D => n1720, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => N342, D => n1724, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => N342, D => n1728, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => N342, D => n1732, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => N342, D => n1736, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => N342, D => n1740, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => N342, D => n1744, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N342, D => n1748, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => N342, D => n1752, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N342, D => n1756, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N342, D => n1760, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N342, D => n1764, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => N342, D => n1768, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => N342, D => n1772, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => N342, D => n1776, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => N342, D => n1780, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => N342, D => n1784, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => N341, D => n1699, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => N341, D => n1702, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => N341, D => n1705, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => N341, D => n1708, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => N341, D => n1711, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => N341, D => n1714, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => N341, D => n1717, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => N341, D => n1720, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => N341, D => n1724, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => N341, D => n1728, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => N341, D => n1732, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => N341, D => n1736, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => N341, D => n1740, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => N341, D => n1744, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N341, D => n1748, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => N341, D => n1752, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N341, D => n1756, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N341, D => n1760, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N341, D => n1764, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => N341, D => n1768, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => N341, D => n1772, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => N341, D => n1776, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => N341, D => n1780, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => N341, D => n1784, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => N340, D => n1699, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => N340, D => n1702, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => N340, D => n1705, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => N340, D => n1708, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => N340, D => n1711, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => N340, D => n1714, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => N340, D => n1717, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => N340, D => n1720, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => N340, D => n1724, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => N340, D => n1728, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => N340, D => n1732, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => N340, D => n1736, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => N340, D => n1740, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => N340, D => n1744, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N340, D => n1748, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => N340, D => n1752, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N340, D => n1756, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N340, D => n1760, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N340, D => n1764, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => N340, D => n1768, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => N340, D => n1772, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => N340, D => n1776, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => N340, D => n1780, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => N340, D => n1784, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => N339, D => n1699, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => N339, D => n1702, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => N339, D => n1705, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => N339, D => n1708, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => N339, D => n1711, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => N339, D => n1714, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => N339, D => n1717, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => N339, D => n1720, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => N339, D => n1724, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => N339, D => n1728, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => N339, D => n1732, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => N339, D => n1736, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => N339, D => n1740, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => N339, D => n1744, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N339, D => n1748, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => N339, D => n1752, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N339, D => n1756, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N339, D => n1760, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N339, D => n1764, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => N339, D => n1768, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => N339, D => n1772, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => N339, D => n1776, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => N339, D => n1780, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => N339, D => n1784, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => N338, D => n1699, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => N338, D => n1702, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => N338, D => n1705, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => N338, D => n1708, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => N338, D => n1711, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => N338, D => n1714, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => N338, D => n1717, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => N338, D => n1720, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => N338, D => n1724, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => N338, D => n1728, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => N338, D => n1732, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => N338, D => n1736, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => N338, D => n1740, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => N338, D => n1744, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N338, D => n1748, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => N338, D => n1752, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N338, D => n1756, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N338, D => n1760, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N338, D => n1764, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => N338, D => n1768, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => N338, D => n1772, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => N338, D => n1776, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => N338, D => n1780, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => N338, D => n1784, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => N337, D => n1699, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => N337, D => n1702, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => N337, D => n1705, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => N337, D => n1708, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => N337, D => n1711, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => N337, D => n1714, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => N337, D => n1717, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => N337, D => n1720, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => N337, D => n1724, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => N337, D => n1728, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => N337, D => n1732, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => N337, D => n1736, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => N337, D => n1740, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => N337, D => n1744, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N337, D => n1748, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => N337, D => n1752, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N337, D => n1756, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N337, D => n1760, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N337, D => n1764, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => N337, D => n1768, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => N337, D => n1772, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => N337, D => n1776, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => N337, D => n1780, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => N337, D => n1784, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => N336, D => n1699, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => N336, D => n1702, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => N336, D => n1705, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => N336, D => n1708, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => N336, D => n1711, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => N336, D => n1714, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => N336, D => n1717, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => N336, D => n1720, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => N336, D => n1724, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => N336, D => n1728, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => N336, D => n1732, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => N336, D => n1736, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => N336, D => n1740, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => N336, D => n1744, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N336, D => n1748, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => N336, D => n1752, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N336, D => n1756, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N336, D => n1760, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N336, D => n1764, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => N336, D => n1768, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => N336, D => n1772, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => N336, D => n1776, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => N336, D => n1780, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => N336, D => n1784, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => N335, D => n1699, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => N335, D => n1702, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => N335, D => n1705, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => N335, D => n1708, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => N335, D => n1711, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => N335, D => n1714, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => N335, D => n1717, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => N335, D => n1720, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => N335, D => n1724, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => N335, D => n1728, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => N335, D => n1732, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => N335, D => n1736, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => N335, D => n1740, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => N335, D => n1744, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N335, D => n1748, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => N335, D => n1752, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N335, D => n1756, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N335, D => n1760, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N335, D => n1764, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => N335, D => n1768, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => N335, D => n1772, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => N335, D => n1776, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => N335, D => n1780, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => N335, D => n1784, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => N334, D => n1699, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => N334, D => n1702, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => N334, D => n1705, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => N334, D => n1708, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => N334, D => n1711, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => N334, D => n1714, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => N334, D => n1717, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => N334, D => n1720, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => N334, D => n1724, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => N334, D => n1728, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => N334, D => n1732, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => N334, D => n1736, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => N334, D => n1740, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => N334, D => n1744, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N334, D => n1748, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => N334, D => n1752, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N334, D => n1756, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N334, D => n1760, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N334, D => n1764, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => N334, D => n1768, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => N334, D => n1772, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => N334, D => n1776, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => N334, D => n1780, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => N334, D => n1784, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => N333, D => n1699, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => N333, D => n1702, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => N333, D => n1705, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => N333, D => n1708, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => N333, D => n1711, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => N333, D => n1714, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => N333, D => n1717, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => N333, D => n1720, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => N333, D => n1724, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => N333, D => n1728, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => N333, D => n1732, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => N333, D => n1736, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => N333, D => n1740, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => N333, D => n1744, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N333, D => n1748, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => N333, D => n1752, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N333, D => n1756, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N333, D => n1760, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N333, D => n1764, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => N333, D => n1768, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => N333, D => n1772, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => N333, D => n1776, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => N333, D => n1780, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => N333, D => n1784, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => N332, D => n1699, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => N332, D => n1702, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => N332, D => n1705, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => N332, D => n1708, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => N332, D => n1711, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => N332, D => n1714, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => N332, D => n1717, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => N332, D => n1720, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => N332, D => n1724, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => N332, D => n1728, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => N332, D => n1732, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => N332, D => n1736, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => N332, D => n1740, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => N332, D => n1744, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N332, D => n1748, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => N332, D => n1752, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N332, D => n1756, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N332, D => n1760, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N332, D => n1764, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => N332, D => n1768, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => N332, D => n1772, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => N332, D => n1776, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => N332, D => n1780, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => N332, D => n1784, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => N331, D => n1721, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => N331, D => n1725, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => N331, D => n1729, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => N331, D => n1733, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => N331, D => n1737, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => N331, D => n1741, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => N331, D => n1745, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N331, D => n1749, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => N331, D => n1753, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N331, D => n1757, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N331, D => n1761, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N331, D => n1765, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => N331, D => n1769, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => N331, D => n1773, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => N331, D => n1777, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => N331, D => n1781, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => N331, D => n1785, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => N330, D => n1721, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => N330, D => n1725, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => N330, D => n1729, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => N330, D => n1733, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => N330, D => n1737, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => N330, D => n1741, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N330, D => n1745, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N330, D => n1749, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => N330, D => n1753, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N330, D => n1757, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N330, D => n1761, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => N330, D => n1765, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => N330, D => n1769, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => N330, D => n1773, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => N330, D => n1777, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => N330, D => n1781, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => N330, D => n1785, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => N329, D => n1721, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => N329, D => n1725, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => N329, D => n1729, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => N329, D => n1733, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => N329, D => n1737, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => N329, D => n1741, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => N329, D => n1745, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N329, D => n1749, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => N329, D => n1753, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N329, D => n1757, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N329, D => n1761, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N329, D => n1765, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => N329, D => n1769, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => N329, D => n1773, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => N329, D => n1777, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => N329, D => n1781, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => N329, D => n1785, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => N328, D => n1721, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => N328, D => n1725, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => N328, D => n1729, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => N328, D => n1733, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => N328, D => n1737, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => N328, D => n1741, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => N328, D => n1745, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N328, D => n1749, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => N328, D => n1753, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N328, D => n1757, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N328, D => n1761, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N328, D => n1765, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => N328, D => n1769, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => N328, D => n1773, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => N328, D => n1777, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => N328, D => n1781, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => N328, D => n1785, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => N327, D => n1721, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => N327, D => n1725, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => N327, D => n1729, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => N327, D => n1733, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => N327, D => n1737, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => N327, D => n1741, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => N327, D => n1745, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N327, D => n1749, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => N327, D => n1753, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N327, D => n1757, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N327, D => n1761, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N327, D => n1765, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => N327, D => n1769, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => N327, D => n1773, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => N327, D => n1777, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => N327, D => n1781, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => N327, D => n1785, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => N326, D => n1721, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => N326, D => n1725, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => N326, D => n1729, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => N326, D => n1733, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => N326, D => n1737, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => N326, D => n1741, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => N326, D => n1745, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N326, D => n1749, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => N326, D => n1753, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N326, D => n1757, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N326, D => n1761, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N326, D => n1765, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => N326, D => n1769, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => N326, D => n1773, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => N326, D => n1777, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => N326, D => n1781, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => N326, D => n1785, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => N325, D => n1721, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => N325, D => n1725, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => N325, D => n1729, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => N325, D => n1733, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => N325, D => n1737, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => N325, D => n1741, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => N325, D => n1745, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N325, D => n1749, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => N325, D => n1753, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N325, D => n1757, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N325, D => n1761, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N325, D => n1765, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => N325, D => n1769, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => N325, D => n1773, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => N325, D => n1777, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => N325, D => n1781, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => N325, D => n1785, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => N324, D => n1721, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => N324, D => n1725, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => N324, D => n1729, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => N324, D => n1733, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => N324, D => n1737, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => N324, D => n1741, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => N324, D => n1745, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N324, D => n1749, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => N324, D => n1753, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N324, D => n1757, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N324, D => n1761, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N324, D => n1765, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => N324, D => n1769, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => N324, D => n1773, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => N324, D => n1777, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => N324, D => n1781, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => N324, D => n1785, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N323, D => n1757, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N323, D => n1761, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N323, D => n1765, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => N323, D => n1769, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => N323, D => n1773, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => N323, D => n1777, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => N323, D => n1781, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => N323, D => n1785, Q => 
                           REGISTERS_31_0_port);
   OUT2_reg_31_inst : DLH_X1 port map( G => CLK, D => N322, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => CLK, D => N321, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => CLK, D => N320, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => CLK, D => N319, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => CLK, D => N318, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => CLK, D => N317, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => CLK, D => N316, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => CLK, D => N315, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => CLK, D => N314, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => CLK, D => N313, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => CLK, D => N312, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => CLK, D => N311, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => CLK, D => N310, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => CLK, D => N309, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => CLK, D => N308, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => CLK, D => N307, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => CLK, D => N306, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => CLK, D => N305, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => CLK, D => N304, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => CLK, D => N303, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => CLK, D => N302, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => CLK, D => N301, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => CLK, D => N300, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => CLK, D => N299, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => CLK, D => N298, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => CLK, D => N297, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => CLK, D => N296, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => CLK, D => N295, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => CLK, D => N294, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => CLK, D => N293, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => CLK, D => N292, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => CLK, D => N291, Q => OUT2(0));
   U35 : OAI21_X2 port map( B1 => n9, B2 => n10, A => n8, ZN => N353);
   U36 : OAI21_X2 port map( B1 => n9, B2 => n11, A => n8, ZN => N352);
   U37 : OAI21_X2 port map( B1 => n9, B2 => n12, A => n8, ZN => N351);
   U38 : OAI21_X2 port map( B1 => n9, B2 => n13, A => n8, ZN => N350);
   U39 : OAI21_X2 port map( B1 => n9, B2 => n14, A => n8, ZN => N349);
   U40 : OAI21_X2 port map( B1 => n9, B2 => n15, A => n8, ZN => N348);
   U41 : OAI21_X2 port map( B1 => n9, B2 => n16, A => n8, ZN => N347);
   U42 : OAI21_X2 port map( B1 => n18, B2 => n19, A => n8, ZN => N346);
   U43 : OAI21_X2 port map( B1 => n10, B2 => n18, A => n8, ZN => N345);
   U44 : OAI21_X2 port map( B1 => n11, B2 => n18, A => n8, ZN => N344);
   U45 : OAI21_X2 port map( B1 => n12, B2 => n18, A => n8, ZN => N343);
   U46 : OAI21_X2 port map( B1 => n13, B2 => n18, A => n8, ZN => N342);
   U47 : OAI21_X2 port map( B1 => n14, B2 => n18, A => n8, ZN => N341);
   U48 : OAI21_X2 port map( B1 => n15, B2 => n18, A => n8, ZN => N340);
   U49 : OAI21_X2 port map( B1 => n16, B2 => n18, A => n8, ZN => N339);
   U50 : OAI21_X2 port map( B1 => n19, B2 => n20, A => n8, ZN => N338);
   U51 : OAI21_X2 port map( B1 => n10, B2 => n20, A => n8, ZN => N337);
   U52 : OAI21_X2 port map( B1 => n11, B2 => n20, A => n8, ZN => N336);
   U53 : OAI21_X2 port map( B1 => n12, B2 => n20, A => n8, ZN => N335);
   U54 : OAI21_X2 port map( B1 => n13, B2 => n20, A => n8, ZN => N334);
   U55 : OAI21_X2 port map( B1 => n14, B2 => n20, A => n8, ZN => N333);
   U56 : OAI21_X2 port map( B1 => n15, B2 => n20, A => n8, ZN => N332);
   U57 : OAI21_X2 port map( B1 => n16, B2 => n20, A => n8, ZN => N331);
   U58 : OAI21_X2 port map( B1 => n19, B2 => n21, A => n8, ZN => N330);
   U59 : OAI21_X2 port map( B1 => n10, B2 => n21, A => n8, ZN => N329);
   U60 : OAI21_X2 port map( B1 => n11, B2 => n21, A => n8, ZN => N328);
   U61 : OAI21_X2 port map( B1 => n12, B2 => n21, A => n8, ZN => N327);
   U62 : OAI21_X2 port map( B1 => n13, B2 => n21, A => n8, ZN => N326);
   U63 : OAI21_X2 port map( B1 => n14, B2 => n21, A => n8, ZN => N325);
   U64 : OAI21_X2 port map( B1 => n15, B2 => n21, A => n8, ZN => N324);
   U65 : OAI21_X2 port map( B1 => n16, B2 => n21, A => n8, ZN => N323);
   U66 : NAND2_X2 port map( A1 => n1787, A2 => n1, ZN => n8);
   U177 : NAND3_X1 port map( A1 => n1793, A2 => n1792, A3 => n17, ZN => n9);
   U178 : NAND3_X1 port map( A1 => n17, A2 => n1792, A3 => ADD_WR(3), ZN => n18
                           );
   U179 : NAND3_X1 port map( A1 => n17, A2 => n1793, A3 => ADD_WR(4), ZN => n20
                           );
   U180 : NAND3_X1 port map( A1 => n1795, A2 => n1794, A3 => n1796, ZN => n19);
   U181 : NAND3_X1 port map( A1 => n1795, A2 => n1794, A3 => ADD_WR(0), ZN => 
                           n10);
   U182 : NAND3_X1 port map( A1 => n1796, A2 => n1794, A3 => ADD_WR(1), ZN => 
                           n11);
   U183 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1794, A3 => ADD_WR(1), ZN 
                           => n12);
   U184 : NAND3_X1 port map( A1 => n1796, A2 => n1795, A3 => ADD_WR(2), ZN => 
                           n13);
   U185 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1795, A3 => ADD_WR(2), ZN 
                           => n14);
   U186 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n1796, A3 => ADD_WR(2), ZN 
                           => n15);
   U187 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n17, A3 => ADD_WR(4), ZN =>
                           n21);
   U188 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n16);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => N323, D => N159, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => N324, D => N159, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => N325, D => N159, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => N326, D => N159, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => N327, D => N159, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => N328, D => N159, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => N329, D => N159, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => N330, D => N159, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => N331, D => N159, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => N323, D => N136, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => N323, D => N135, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => N323, D => N134, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => N323, D => N133, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => N323, D => N132, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => N323, D => N131, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => N324, D => N136, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => N324, D => N135, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => N324, D => N134, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => N324, D => N133, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => N324, D => N132, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => N324, D => N131, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => N325, D => N136, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => N325, D => N135, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => N325, D => N134, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => N325, D => N133, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => N325, D => N132, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => N325, D => N131, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => N326, D => N136, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => N326, D => N135, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => N326, D => N134, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => N326, D => N133, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => N326, D => N132, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => N326, D => N131, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => N327, D => N136, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => N327, D => N135, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => N327, D => N134, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => N327, D => N133, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => N327, D => N132, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => N327, D => N131, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => N328, D => N136, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => N328, D => N135, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => N328, D => N134, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => N328, D => N133, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => N328, D => N132, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => N328, D => N131, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => N329, D => N136, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => N329, D => N135, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => N329, D => N134, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => N329, D => N133, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => N329, D => N132, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => N329, D => N131, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => N330, D => N136, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => N330, D => N135, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => N330, D => N134, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => N330, D => N133, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => N330, D => N132, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => N330, D => N131, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => N331, D => N136, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => N331, D => N135, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => N331, D => N134, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => N331, D => N133, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => N331, D => N132, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => N331, D => N131, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => N323, D => N137, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => N324, D => N137, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => N325, D => N137, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => N326, D => N137, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => N327, D => N137, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => N328, D => N137, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => N329, D => N137, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => N330, D => N137, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => N331, D => N137, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => N332, D => N159, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => N333, D => N159, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => N334, D => N159, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => N335, D => N159, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => N336, D => N159, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => N337, D => N159, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => N338, D => N159, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => N339, D => N159, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => N340, D => N159, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => N341, D => N159, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => N342, D => N159, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => N343, D => N159, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => N344, D => N159, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => N345, D => N159, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => N346, D => N159, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => N347, D => N159, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => N348, D => N159, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => N349, D => N159, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => N350, D => N159, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => N351, D => N159, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => N352, D => N159, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => N353, D => N159, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => N332, D => N136, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => N332, D => N135, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => N332, D => N134, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => N332, D => N133, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => N332, D => N132, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => N332, D => N131, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => N333, D => N136, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => N333, D => N135, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => N333, D => N134, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => N333, D => N133, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => N333, D => N132, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => N333, D => N131, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => N334, D => N136, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => N334, D => N135, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => N334, D => N134, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => N334, D => N133, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => N334, D => N132, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => N334, D => N131, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => N335, D => N136, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => N335, D => N135, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => N335, D => N134, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => N335, D => N133, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => N335, D => N132, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => N335, D => N131, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => N336, D => N136, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => N336, D => N135, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => N336, D => N134, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => N336, D => N133, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => N336, D => N132, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => N336, D => N131, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => N337, D => N136, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => N337, D => N135, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => N337, D => N134, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => N337, D => N133, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => N337, D => N132, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => N337, D => N131, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => N338, D => N136, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => N338, D => N135, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => N338, D => N134, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => N338, D => N133, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => N338, D => N132, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => N338, D => N131, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => N339, D => N136, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => N339, D => N135, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => N339, D => N134, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => N339, D => N133, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => N339, D => N132, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => N339, D => N131, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => N340, D => N136, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => N340, D => N135, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => N340, D => N134, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => N340, D => N133, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => N340, D => N132, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => N340, D => N131, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => N341, D => N136, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => N341, D => N135, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => N341, D => N134, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => N341, D => N133, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => N341, D => N132, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => N341, D => N131, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => N342, D => N136, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => N342, D => N135, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => N342, D => N134, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => N342, D => N133, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => N342, D => N132, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => N342, D => N131, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => N343, D => N136, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => N343, D => N135, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => N343, D => N134, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => N343, D => N133, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => N343, D => N132, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => N343, D => N131, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => N344, D => N136, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => N344, D => N135, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => N344, D => N134, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => N344, D => N133, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => N344, D => N132, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => N344, D => N131, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => N345, D => N136, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => N345, D => N135, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => N345, D => N134, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => N345, D => N133, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => N345, D => N132, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => N345, D => N131, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => N346, D => N136, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => N346, D => N135, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => N346, D => N134, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => N346, D => N133, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => N346, D => N132, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => N346, D => N131, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => N347, D => N136, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => N347, D => N135, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => N347, D => N134, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => N347, D => N133, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => N347, D => N132, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => N347, D => N131, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => N348, D => N136, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => N348, D => N135, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => N348, D => N134, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => N348, D => N133, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => N348, D => N132, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => N348, D => N131, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => N349, D => N136, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => N349, D => N135, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => N349, D => N134, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => N349, D => N133, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => N349, D => N132, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => N349, D => N131, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => N350, D => N136, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => N350, D => N135, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => N350, D => N134, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => N350, D => N133, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => N350, D => N132, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => N350, D => N131, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => N351, D => N136, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => N351, D => N135, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => N351, D => N134, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => N351, D => N133, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => N351, D => N132, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => N351, D => N131, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => N352, D => N136, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => N352, D => N135, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => N352, D => N134, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => N352, D => N133, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => N352, D => N132, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => N352, D => N131, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => N353, D => N136, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => N353, D => N135, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => N353, D => N134, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => N353, D => N133, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => N353, D => N132, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => N353, D => N131, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => N332, D => N137, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => N333, D => N137, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => N334, D => N137, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => N335, D => N137, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => N336, D => N137, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => N337, D => N137, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => N338, D => N137, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => N339, D => N137, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => N340, D => N137, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => N341, D => N137, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => N342, D => N137, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => N343, D => N137, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => N344, D => N137, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => N345, D => N137, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => N346, D => N137, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => N347, D => N137, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => N348, D => N137, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => N349, D => N137, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => N350, D => N137, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => N351, D => N137, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => N352, D => N137, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => N353, D => N137, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => N323, D => N158, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => N323, D => N157, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => N323, D => N156, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => N323, D => N155, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => N323, D => N154, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => N323, D => N153, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => N323, D => N152, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => N324, D => N158, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => N324, D => N157, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => N324, D => N156, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => N324, D => N155, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => N324, D => N154, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => N324, D => N153, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => N324, D => N152, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => N325, D => N158, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => N325, D => N157, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => N325, D => N156, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => N325, D => N155, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => N325, D => N154, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => N325, D => N153, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => N325, D => N152, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => N326, D => N158, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => N326, D => N157, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => N326, D => N156, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => N326, D => N155, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => N326, D => N154, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => N326, D => N153, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => N326, D => N152, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => N327, D => N158, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => N327, D => N157, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => N327, D => N156, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => N327, D => N155, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => N327, D => N154, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => N327, D => N153, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => N327, D => N152, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => N328, D => N158, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => N328, D => N157, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => N328, D => N156, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => N328, D => N155, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => N328, D => N154, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => N328, D => N153, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => N328, D => N152, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => N329, D => N158, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => N329, D => N157, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => N329, D => N156, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => N329, D => N155, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => N329, D => N154, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => N329, D => N153, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => N329, D => N152, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => N330, D => N158, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => N330, D => N157, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => N330, D => N156, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => N330, D => N155, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => N330, D => N154, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => N330, D => N153, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => N330, D => N152, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => N331, D => N158, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => N331, D => N157, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => N331, D => N156, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => N331, D => N155, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => N331, D => N154, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => N331, D => N153, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => N331, D => N152, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => N323, D => N151, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => N323, D => N150, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => N323, D => N149, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => N323, D => N148, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => N323, D => N147, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => N323, D => N146, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => N323, D => N145, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N323, D => N144, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => N323, D => N143, Q => 
                           REGISTERS_31_15_port);
   U3 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n863, ZN => n2);
   U4 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n35, ZN => n3);
   U5 : AND2_X1 port map( A1 => n862, A2 => ADD_RD2(0), ZN => n4);
   U6 : AND2_X1 port map( A1 => n865, A2 => ADD_RD2(0), ZN => n5);
   U7 : AND2_X1 port map( A1 => n864, A2 => ADD_RD2(0), ZN => n6);
   U8 : AND2_X1 port map( A1 => n34, A2 => ADD_RD1(0), ZN => n7);
   U9 : AND2_X1 port map( A1 => n37, A2 => ADD_RD1(0), ZN => n28);
   U10 : AND2_X1 port map( A1 => n36, A2 => ADD_RD1(0), ZN => n29);
   U11 : AND2_X1 port map( A1 => n34, A2 => n716, ZN => n30);
   U12 : AND2_X1 port map( A1 => n862, A2 => n1544, ZN => n31);
   U13 : AND2_X1 port map( A1 => n35, A2 => n716, ZN => n32);
   U14 : AND2_X1 port map( A1 => n863, A2 => n1544, ZN => n33);
   U15 : BUF_X1 port map( A => n1787, Z => n1791);
   U16 : BUF_X1 port map( A => n1634, Z => n1636);
   U17 : BUF_X1 port map( A => n1617, Z => n1619);
   U18 : BUF_X1 port map( A => n1634, Z => n1637);
   U19 : BUF_X1 port map( A => n1617, Z => n1620);
   U20 : BUF_X1 port map( A => n806, Z => n808);
   U21 : BUF_X1 port map( A => n789, Z => n791);
   U22 : BUF_X1 port map( A => n806, Z => n809);
   U23 : BUF_X1 port map( A => n789, Z => n792);
   U24 : BUF_X1 port map( A => n31, Z => n1634);
   U25 : BUF_X1 port map( A => n33, Z => n1617);
   U26 : BUF_X1 port map( A => n30, Z => n806);
   U27 : BUF_X1 port map( A => n32, Z => n789);
   U28 : BUF_X1 port map( A => n1600, Z => n1602);
   U29 : BUF_X1 port map( A => n1583, Z => n1585);
   U30 : BUF_X1 port map( A => n1566, Z => n1568);
   U31 : BUF_X1 port map( A => n1549, Z => n1551);
   U32 : BUF_X1 port map( A => n1662, Z => n1664);
   U33 : BUF_X1 port map( A => n1600, Z => n1603);
   U34 : BUF_X1 port map( A => n1583, Z => n1586);
   U67 : BUF_X1 port map( A => n1566, Z => n1569);
   U68 : BUF_X1 port map( A => n1549, Z => n1552);
   U69 : BUF_X1 port map( A => n1662, Z => n1665);
   U70 : BUF_X1 port map( A => n1650, Z => n1653);
   U71 : BUF_X1 port map( A => n772, Z => n774);
   U72 : BUF_X1 port map( A => n755, Z => n757);
   U73 : BUF_X1 port map( A => n738, Z => n740);
   U74 : BUF_X1 port map( A => n721, Z => n723);
   U75 : BUF_X1 port map( A => n834, Z => n836);
   U76 : BUF_X1 port map( A => n772, Z => n775);
   U77 : BUF_X1 port map( A => n755, Z => n758);
   U78 : BUF_X1 port map( A => n738, Z => n741);
   U79 : BUF_X1 port map( A => n721, Z => n724);
   U80 : BUF_X1 port map( A => n834, Z => n837);
   U81 : BUF_X1 port map( A => n822, Z => n825);
   U82 : BUF_X1 port map( A => n1650, Z => n1652);
   U83 : BUF_X1 port map( A => n822, Z => n824);
   U84 : BUF_X1 port map( A => n1633, Z => n1638);
   U85 : BUF_X1 port map( A => n1616, Z => n1621);
   U86 : BUF_X1 port map( A => n805, Z => n810);
   U87 : BUF_X1 port map( A => n788, Z => n793);
   U88 : BUF_X1 port map( A => N128, Z => n1786);
   U89 : BUF_X1 port map( A => N129, Z => n1782);
   U90 : BUF_X1 port map( A => N130, Z => n1778);
   U91 : BUF_X1 port map( A => N138, Z => n1774);
   U92 : BUF_X1 port map( A => N139, Z => n1770);
   U93 : BUF_X1 port map( A => N140, Z => n1766);
   U94 : BUF_X1 port map( A => N141, Z => n1762);
   U95 : BUF_X1 port map( A => N142, Z => n1758);
   U96 : BUF_X1 port map( A => N143, Z => n1754);
   U97 : BUF_X1 port map( A => N144, Z => n1750);
   U98 : BUF_X1 port map( A => N145, Z => n1746);
   U99 : BUF_X1 port map( A => N146, Z => n1742);
   U100 : BUF_X1 port map( A => N147, Z => n1738);
   U101 : BUF_X1 port map( A => N148, Z => n1734);
   U102 : BUF_X1 port map( A => N149, Z => n1730);
   U103 : BUF_X1 port map( A => N150, Z => n1726);
   U104 : BUF_X1 port map( A => N151, Z => n1722);
   U105 : BUF_X1 port map( A => N152, Z => n1718);
   U106 : BUF_X1 port map( A => N153, Z => n1715);
   U107 : BUF_X1 port map( A => N154, Z => n1712);
   U108 : BUF_X1 port map( A => N155, Z => n1709);
   U109 : BUF_X1 port map( A => N156, Z => n1706);
   U110 : BUF_X1 port map( A => N157, Z => n1703);
   U111 : BUF_X1 port map( A => N158, Z => n1700);
   U112 : BUF_X1 port map( A => n2, Z => n1549);
   U113 : BUF_X1 port map( A => n6, Z => n1600);
   U114 : BUF_X1 port map( A => n5, Z => n1583);
   U115 : BUF_X1 port map( A => n4, Z => n1566);
   U116 : BUF_X1 port map( A => n29, Z => n772);
   U117 : BUF_X1 port map( A => n28, Z => n755);
   U118 : BUF_X1 port map( A => n7, Z => n738);
   U119 : BUF_X1 port map( A => n3, Z => n721);
   U120 : BUF_X1 port map( A => n1530, Z => n1662);
   U121 : BUF_X1 port map( A => n1529, Z => n1650);
   U122 : BUF_X1 port map( A => n702, Z => n834);
   U123 : BUF_X1 port map( A => n701, Z => n822);
   U124 : BUF_X1 port map( A => n1599, Z => n1604);
   U125 : BUF_X1 port map( A => n1582, Z => n1587);
   U126 : BUF_X1 port map( A => n1565, Z => n1570);
   U127 : BUF_X1 port map( A => n1548, Z => n1553);
   U128 : BUF_X1 port map( A => n771, Z => n776);
   U129 : BUF_X1 port map( A => n754, Z => n759);
   U130 : BUF_X1 port map( A => n737, Z => n742);
   U131 : BUF_X1 port map( A => n720, Z => n725);
   U132 : BUF_X1 port map( A => n712, Z => n854);
   U133 : BUF_X1 port map( A => n714, Z => n858);
   U134 : BUF_X1 port map( A => n710, Z => n850);
   U135 : BUF_X1 port map( A => n708, Z => n846);
   U136 : BUF_X1 port map( A => n1538, Z => n1678);
   U137 : BUF_X1 port map( A => n1536, Z => n1674);
   U138 : BUF_X1 port map( A => n1540, Z => n1682);
   U139 : BUF_X1 port map( A => n1542, Z => n1686);
   U140 : BUF_X1 port map( A => n22, Z => n1697);
   U141 : BUF_X1 port map( A => n25, Z => n1693);
   U142 : BUF_X1 port map( A => n1636, Z => n1647);
   U143 : BUF_X1 port map( A => n1636, Z => n1646);
   U144 : BUF_X1 port map( A => n1636, Z => n1645);
   U145 : BUF_X1 port map( A => n1637, Z => n1644);
   U146 : BUF_X1 port map( A => n1637, Z => n1643);
   U147 : BUF_X1 port map( A => n1637, Z => n1642);
   U148 : BUF_X1 port map( A => n808, Z => n819);
   U149 : BUF_X1 port map( A => n808, Z => n818);
   U150 : BUF_X1 port map( A => n808, Z => n817);
   U151 : BUF_X1 port map( A => n809, Z => n816);
   U152 : BUF_X1 port map( A => n809, Z => n815);
   U153 : BUF_X1 port map( A => n809, Z => n814);
   U154 : BUF_X1 port map( A => n1635, Z => n1649);
   U155 : BUF_X1 port map( A => n1635, Z => n1648);
   U156 : BUF_X1 port map( A => n807, Z => n821);
   U157 : BUF_X1 port map( A => n807, Z => n820);
   U158 : BUF_X1 port map( A => n1619, Z => n1630);
   U159 : BUF_X1 port map( A => n1619, Z => n1629);
   U160 : BUF_X1 port map( A => n1619, Z => n1628);
   U161 : BUF_X1 port map( A => n1620, Z => n1627);
   U162 : BUF_X1 port map( A => n1620, Z => n1626);
   U163 : BUF_X1 port map( A => n1620, Z => n1625);
   U164 : BUF_X1 port map( A => n791, Z => n802);
   U165 : BUF_X1 port map( A => n791, Z => n801);
   U166 : BUF_X1 port map( A => n791, Z => n800);
   U167 : BUF_X1 port map( A => n792, Z => n799);
   U168 : BUF_X1 port map( A => n792, Z => n798);
   U169 : BUF_X1 port map( A => n792, Z => n797);
   U170 : BUF_X1 port map( A => n1618, Z => n1632);
   U171 : BUF_X1 port map( A => n1618, Z => n1631);
   U172 : BUF_X1 port map( A => n790, Z => n804);
   U173 : BUF_X1 port map( A => n790, Z => n803);
   U174 : INV_X1 port map( A => n1791, ZN => n1788);
   U175 : INV_X1 port map( A => n1791, ZN => n1789);
   U176 : INV_X1 port map( A => n1791, ZN => n1790);
   U189 : BUF_X1 port map( A => n1634, Z => n1635);
   U190 : BUF_X1 port map( A => n1617, Z => n1618);
   U191 : BUF_X1 port map( A => n806, Z => n807);
   U192 : BUF_X1 port map( A => n789, Z => n790);
   U193 : BUF_X1 port map( A => n1652, Z => n1659);
   U194 : BUF_X1 port map( A => n824, Z => n831);
   U195 : BUF_X1 port map( A => n1651, Z => n1661);
   U196 : BUF_X1 port map( A => n1651, Z => n1660);
   U197 : BUF_X1 port map( A => n823, Z => n833);
   U198 : BUF_X1 port map( A => n823, Z => n832);
   U199 : BUF_X1 port map( A => n1652, Z => n1658);
   U200 : BUF_X1 port map( A => n1653, Z => n1655);
   U201 : BUF_X1 port map( A => n824, Z => n830);
   U202 : BUF_X1 port map( A => n825, Z => n827);
   U203 : BUF_X1 port map( A => n1652, Z => n1657);
   U204 : BUF_X1 port map( A => n1653, Z => n1656);
   U205 : BUF_X1 port map( A => n824, Z => n829);
   U206 : BUF_X1 port map( A => n825, Z => n828);
   U207 : BUF_X1 port map( A => n1602, Z => n1613);
   U208 : BUF_X1 port map( A => n1568, Z => n1579);
   U209 : BUF_X1 port map( A => n1664, Z => n1671);
   U210 : BUF_X1 port map( A => n1602, Z => n1612);
   U211 : BUF_X1 port map( A => n1568, Z => n1578);
   U212 : BUF_X1 port map( A => n1602, Z => n1611);
   U213 : BUF_X1 port map( A => n1568, Z => n1577);
   U214 : BUF_X1 port map( A => n1664, Z => n1670);
   U215 : BUF_X1 port map( A => n1603, Z => n1610);
   U216 : BUF_X1 port map( A => n1569, Z => n1576);
   U217 : BUF_X1 port map( A => n1664, Z => n1669);
   U218 : BUF_X1 port map( A => n1603, Z => n1609);
   U219 : BUF_X1 port map( A => n1569, Z => n1575);
   U220 : BUF_X1 port map( A => n1665, Z => n1668);
   U221 : BUF_X1 port map( A => n1603, Z => n1608);
   U222 : BUF_X1 port map( A => n1569, Z => n1574);
   U223 : BUF_X1 port map( A => n1665, Z => n1667);
   U224 : BUF_X1 port map( A => n1665, Z => n1666);
   U225 : BUF_X1 port map( A => n774, Z => n785);
   U226 : BUF_X1 port map( A => n740, Z => n751);
   U227 : BUF_X1 port map( A => n836, Z => n843);
   U228 : BUF_X1 port map( A => n774, Z => n784);
   U229 : BUF_X1 port map( A => n740, Z => n750);
   U230 : BUF_X1 port map( A => n774, Z => n783);
   U231 : BUF_X1 port map( A => n740, Z => n749);
   U232 : BUF_X1 port map( A => n836, Z => n842);
   U233 : BUF_X1 port map( A => n775, Z => n782);
   U234 : BUF_X1 port map( A => n741, Z => n748);
   U235 : BUF_X1 port map( A => n836, Z => n841);
   U236 : BUF_X1 port map( A => n775, Z => n781);
   U237 : BUF_X1 port map( A => n741, Z => n747);
   U238 : BUF_X1 port map( A => n837, Z => n840);
   U239 : BUF_X1 port map( A => n775, Z => n780);
   U240 : BUF_X1 port map( A => n741, Z => n746);
   U241 : BUF_X1 port map( A => n837, Z => n839);
   U242 : BUF_X1 port map( A => n837, Z => n838);
   U243 : BUF_X1 port map( A => n1638, Z => n1641);
   U244 : BUF_X1 port map( A => n1638, Z => n1640);
   U245 : BUF_X1 port map( A => n810, Z => n813);
   U246 : BUF_X1 port map( A => n810, Z => n812);
   U247 : BUF_X1 port map( A => n1601, Z => n1615);
   U248 : BUF_X1 port map( A => n1567, Z => n1581);
   U249 : BUF_X1 port map( A => n1663, Z => n1673);
   U250 : BUF_X1 port map( A => n1601, Z => n1614);
   U251 : BUF_X1 port map( A => n1567, Z => n1580);
   U252 : BUF_X1 port map( A => n1663, Z => n1672);
   U253 : BUF_X1 port map( A => n773, Z => n787);
   U254 : BUF_X1 port map( A => n739, Z => n753);
   U255 : BUF_X1 port map( A => n835, Z => n845);
   U256 : BUF_X1 port map( A => n773, Z => n786);
   U257 : BUF_X1 port map( A => n739, Z => n752);
   U258 : BUF_X1 port map( A => n835, Z => n844);
   U259 : BUF_X1 port map( A => n1585, Z => n1596);
   U260 : BUF_X1 port map( A => n1551, Z => n1562);
   U261 : BUF_X1 port map( A => n1585, Z => n1595);
   U262 : BUF_X1 port map( A => n1551, Z => n1561);
   U263 : BUF_X1 port map( A => n1585, Z => n1594);
   U264 : BUF_X1 port map( A => n1551, Z => n1560);
   U265 : BUF_X1 port map( A => n1586, Z => n1593);
   U266 : BUF_X1 port map( A => n1552, Z => n1559);
   U267 : BUF_X1 port map( A => n1586, Z => n1592);
   U268 : BUF_X1 port map( A => n1552, Z => n1558);
   U269 : BUF_X1 port map( A => n1586, Z => n1591);
   U270 : BUF_X1 port map( A => n1552, Z => n1557);
   U271 : BUF_X1 port map( A => n1621, Z => n1624);
   U272 : BUF_X1 port map( A => n1621, Z => n1623);
   U273 : BUF_X1 port map( A => n757, Z => n768);
   U274 : BUF_X1 port map( A => n723, Z => n734);
   U275 : BUF_X1 port map( A => n757, Z => n767);
   U276 : BUF_X1 port map( A => n723, Z => n733);
   U277 : BUF_X1 port map( A => n757, Z => n766);
   U278 : BUF_X1 port map( A => n723, Z => n732);
   U279 : BUF_X1 port map( A => n758, Z => n765);
   U280 : BUF_X1 port map( A => n724, Z => n731);
   U281 : BUF_X1 port map( A => n758, Z => n764);
   U282 : BUF_X1 port map( A => n724, Z => n730);
   U283 : BUF_X1 port map( A => n758, Z => n763);
   U284 : BUF_X1 port map( A => n724, Z => n729);
   U285 : BUF_X1 port map( A => n793, Z => n796);
   U286 : BUF_X1 port map( A => n793, Z => n795);
   U287 : BUF_X1 port map( A => n1584, Z => n1598);
   U288 : BUF_X1 port map( A => n1550, Z => n1564);
   U289 : BUF_X1 port map( A => n1584, Z => n1597);
   U290 : BUF_X1 port map( A => n1550, Z => n1563);
   U291 : BUF_X1 port map( A => n756, Z => n770);
   U292 : BUF_X1 port map( A => n722, Z => n736);
   U293 : BUF_X1 port map( A => n756, Z => n769);
   U294 : BUF_X1 port map( A => n722, Z => n735);
   U295 : BUF_X1 port map( A => n1653, Z => n1654);
   U296 : BUF_X1 port map( A => n825, Z => n826);
   U297 : BUF_X1 port map( A => n1638, Z => n1639);
   U298 : BUF_X1 port map( A => n810, Z => n811);
   U299 : BUF_X1 port map( A => n1621, Z => n1622);
   U300 : BUF_X1 port map( A => n793, Z => n794);
   U301 : BUF_X1 port map( A => n1786, Z => n1785);
   U302 : BUF_X1 port map( A => n1782, Z => n1781);
   U303 : BUF_X1 port map( A => n1778, Z => n1777);
   U304 : BUF_X1 port map( A => n1774, Z => n1773);
   U305 : BUF_X1 port map( A => n1770, Z => n1769);
   U306 : BUF_X1 port map( A => n1766, Z => n1765);
   U307 : BUF_X1 port map( A => n1762, Z => n1761);
   U308 : BUF_X1 port map( A => n1758, Z => n1757);
   U309 : BUF_X1 port map( A => n1754, Z => n1753);
   U310 : BUF_X1 port map( A => n1750, Z => n1749);
   U311 : BUF_X1 port map( A => n1746, Z => n1745);
   U312 : BUF_X1 port map( A => n1742, Z => n1741);
   U313 : BUF_X1 port map( A => n1738, Z => n1737);
   U314 : BUF_X1 port map( A => n1734, Z => n1733);
   U315 : BUF_X1 port map( A => n1730, Z => n1729);
   U316 : BUF_X1 port map( A => n1726, Z => n1725);
   U317 : BUF_X1 port map( A => n1722, Z => n1721);
   U318 : BUF_X1 port map( A => n1786, Z => n1784);
   U319 : BUF_X1 port map( A => n1782, Z => n1780);
   U320 : BUF_X1 port map( A => n1778, Z => n1776);
   U321 : BUF_X1 port map( A => n1774, Z => n1772);
   U322 : BUF_X1 port map( A => n1770, Z => n1768);
   U323 : BUF_X1 port map( A => n1766, Z => n1764);
   U324 : BUF_X1 port map( A => n1762, Z => n1760);
   U325 : BUF_X1 port map( A => n1758, Z => n1756);
   U326 : BUF_X1 port map( A => n1754, Z => n1752);
   U327 : BUF_X1 port map( A => n1750, Z => n1748);
   U328 : BUF_X1 port map( A => n1746, Z => n1744);
   U329 : BUF_X1 port map( A => n1742, Z => n1740);
   U330 : BUF_X1 port map( A => n1738, Z => n1736);
   U331 : BUF_X1 port map( A => n1734, Z => n1732);
   U332 : BUF_X1 port map( A => n1730, Z => n1728);
   U333 : BUF_X1 port map( A => n1726, Z => n1724);
   U334 : BUF_X1 port map( A => n1722, Z => n1720);
   U335 : BUF_X1 port map( A => n1718, Z => n1717);
   U336 : BUF_X1 port map( A => n1715, Z => n1714);
   U337 : BUF_X1 port map( A => n1712, Z => n1711);
   U338 : BUF_X1 port map( A => n1709, Z => n1708);
   U339 : BUF_X1 port map( A => n1706, Z => n1705);
   U340 : BUF_X1 port map( A => n1703, Z => n1702);
   U341 : BUF_X1 port map( A => n1700, Z => n1699);
   U342 : BUF_X1 port map( A => n1786, Z => n1783);
   U343 : BUF_X1 port map( A => n1782, Z => n1779);
   U344 : BUF_X1 port map( A => n1778, Z => n1775);
   U345 : BUF_X1 port map( A => n1774, Z => n1771);
   U346 : BUF_X1 port map( A => n1770, Z => n1767);
   U347 : BUF_X1 port map( A => n1766, Z => n1763);
   U348 : BUF_X1 port map( A => n1762, Z => n1759);
   U349 : BUF_X1 port map( A => n1758, Z => n1755);
   U350 : BUF_X1 port map( A => n1754, Z => n1751);
   U351 : BUF_X1 port map( A => n1750, Z => n1747);
   U352 : BUF_X1 port map( A => n1746, Z => n1743);
   U353 : BUF_X1 port map( A => n1742, Z => n1739);
   U354 : BUF_X1 port map( A => n1738, Z => n1735);
   U355 : BUF_X1 port map( A => n1734, Z => n1731);
   U356 : BUF_X1 port map( A => n1730, Z => n1727);
   U357 : BUF_X1 port map( A => n1726, Z => n1723);
   U358 : BUF_X1 port map( A => n1722, Z => n1719);
   U359 : BUF_X1 port map( A => n1718, Z => n1716);
   U360 : BUF_X1 port map( A => n1715, Z => n1713);
   U361 : BUF_X1 port map( A => n1712, Z => n1710);
   U362 : BUF_X1 port map( A => n1709, Z => n1707);
   U363 : BUF_X1 port map( A => n1706, Z => n1704);
   U364 : BUF_X1 port map( A => n1703, Z => n1701);
   U365 : BUF_X1 port map( A => n1700, Z => n1698);
   U366 : BUF_X1 port map( A => n31, Z => n1633);
   U367 : BUF_X1 port map( A => n33, Z => n1616);
   U368 : BUF_X1 port map( A => n30, Z => n805);
   U369 : BUF_X1 port map( A => n32, Z => n788);
   U370 : BUF_X1 port map( A => RESET, Z => n1787);
   U371 : BUF_X1 port map( A => n1662, Z => n1663);
   U372 : BUF_X1 port map( A => n1650, Z => n1651);
   U373 : BUF_X1 port map( A => n834, Z => n835);
   U374 : BUF_X1 port map( A => n822, Z => n823);
   U375 : BUF_X1 port map( A => n1600, Z => n1601);
   U376 : BUF_X1 port map( A => n1583, Z => n1584);
   U377 : BUF_X1 port map( A => n1566, Z => n1567);
   U378 : BUF_X1 port map( A => n1549, Z => n1550);
   U379 : BUF_X1 port map( A => n772, Z => n773);
   U380 : BUF_X1 port map( A => n755, Z => n756);
   U381 : BUF_X1 port map( A => n738, Z => n739);
   U382 : BUF_X1 port map( A => n721, Z => n722);
   U383 : BUF_X1 port map( A => n1604, Z => n1607);
   U384 : BUF_X1 port map( A => n1570, Z => n1573);
   U385 : BUF_X1 port map( A => n1604, Z => n1606);
   U386 : BUF_X1 port map( A => n1570, Z => n1572);
   U387 : BUF_X1 port map( A => n776, Z => n779);
   U388 : BUF_X1 port map( A => n742, Z => n745);
   U389 : BUF_X1 port map( A => n776, Z => n778);
   U390 : BUF_X1 port map( A => n742, Z => n744);
   U391 : BUF_X1 port map( A => n1587, Z => n1590);
   U392 : BUF_X1 port map( A => n1553, Z => n1556);
   U393 : BUF_X1 port map( A => n1587, Z => n1589);
   U394 : BUF_X1 port map( A => n1553, Z => n1555);
   U395 : BUF_X1 port map( A => n759, Z => n762);
   U396 : BUF_X1 port map( A => n725, Z => n728);
   U397 : BUF_X1 port map( A => n759, Z => n761);
   U398 : BUF_X1 port map( A => n725, Z => n727);
   U399 : BUF_X1 port map( A => n1604, Z => n1605);
   U400 : BUF_X1 port map( A => n1570, Z => n1571);
   U401 : BUF_X1 port map( A => n776, Z => n777);
   U402 : BUF_X1 port map( A => n742, Z => n743);
   U403 : BUF_X1 port map( A => n1587, Z => n1588);
   U404 : BUF_X1 port map( A => n1553, Z => n1554);
   U405 : BUF_X1 port map( A => n759, Z => n760);
   U406 : BUF_X1 port map( A => n725, Z => n726);
   U407 : AND2_X1 port map( A1 => DATAIN(9), A2 => n1788, ZN => N137);
   U408 : AND2_X1 port map( A1 => DATAIN(3), A2 => n1788, ZN => N131);
   U409 : AND2_X1 port map( A1 => DATAIN(4), A2 => n1788, ZN => N132);
   U410 : AND2_X1 port map( A1 => DATAIN(5), A2 => n1788, ZN => N133);
   U411 : AND2_X1 port map( A1 => DATAIN(6), A2 => n1788, ZN => N134);
   U412 : AND2_X1 port map( A1 => DATAIN(7), A2 => n1788, ZN => N135);
   U413 : AND2_X1 port map( A1 => DATAIN(8), A2 => n1788, ZN => N136);
   U414 : AND2_X1 port map( A1 => DATAIN(31), A2 => n1790, ZN => N159);
   U415 : AND2_X1 port map( A1 => DATAIN(0), A2 => n1788, ZN => N128);
   U416 : AND2_X1 port map( A1 => DATAIN(1), A2 => n1788, ZN => N129);
   U417 : AND2_X1 port map( A1 => DATAIN(2), A2 => n1788, ZN => N130);
   U418 : AND2_X1 port map( A1 => DATAIN(10), A2 => n1788, ZN => N138);
   U419 : AND2_X1 port map( A1 => DATAIN(11), A2 => n1788, ZN => N139);
   U420 : AND2_X1 port map( A1 => DATAIN(12), A2 => n1789, ZN => N140);
   U421 : AND2_X1 port map( A1 => DATAIN(13), A2 => n1789, ZN => N141);
   U422 : AND2_X1 port map( A1 => DATAIN(14), A2 => n1789, ZN => N142);
   U423 : AND2_X1 port map( A1 => DATAIN(15), A2 => n1789, ZN => N143);
   U424 : AND2_X1 port map( A1 => DATAIN(16), A2 => n1789, ZN => N144);
   U425 : AND2_X1 port map( A1 => DATAIN(17), A2 => n1789, ZN => N145);
   U426 : AND2_X1 port map( A1 => DATAIN(18), A2 => n1789, ZN => N146);
   U427 : AND2_X1 port map( A1 => DATAIN(19), A2 => n1789, ZN => N147);
   U428 : AND2_X1 port map( A1 => DATAIN(20), A2 => n1789, ZN => N148);
   U429 : AND2_X1 port map( A1 => DATAIN(21), A2 => n1789, ZN => N149);
   U430 : AND2_X1 port map( A1 => DATAIN(22), A2 => n1789, ZN => N150);
   U431 : AND2_X1 port map( A1 => DATAIN(23), A2 => n1789, ZN => N151);
   U432 : AND2_X1 port map( A1 => DATAIN(24), A2 => n1790, ZN => N152);
   U433 : AND2_X1 port map( A1 => DATAIN(25), A2 => n1790, ZN => N153);
   U434 : AND2_X1 port map( A1 => DATAIN(26), A2 => n1790, ZN => N154);
   U435 : AND2_X1 port map( A1 => DATAIN(27), A2 => n1790, ZN => N155);
   U436 : AND2_X1 port map( A1 => DATAIN(28), A2 => n1790, ZN => N156);
   U437 : AND2_X1 port map( A1 => DATAIN(29), A2 => n1790, ZN => N157);
   U438 : AND2_X1 port map( A1 => DATAIN(30), A2 => n1790, ZN => N158);
   U439 : BUF_X1 port map( A => n6, Z => n1599);
   U440 : BUF_X1 port map( A => n5, Z => n1582);
   U441 : BUF_X1 port map( A => n4, Z => n1565);
   U442 : BUF_X1 port map( A => n2, Z => n1548);
   U443 : BUF_X1 port map( A => n29, Z => n771);
   U444 : BUF_X1 port map( A => n28, Z => n754);
   U445 : BUF_X1 port map( A => n7, Z => n737);
   U446 : BUF_X1 port map( A => n3, Z => n720);
   U447 : AND2_X1 port map( A1 => N290, A2 => n1696, ZN => N291);
   U448 : AND2_X1 port map( A1 => N289, A2 => n1696, ZN => N292);
   U449 : AND2_X1 port map( A1 => N288, A2 => n1696, ZN => N293);
   U450 : AND2_X1 port map( A1 => N287, A2 => n1696, ZN => N294);
   U451 : AND2_X1 port map( A1 => N286, A2 => n1696, ZN => N295);
   U452 : AND2_X1 port map( A1 => N285, A2 => n1696, ZN => N296);
   U453 : AND2_X1 port map( A1 => N284, A2 => n1696, ZN => N297);
   U454 : AND2_X1 port map( A1 => N283, A2 => n1696, ZN => N298);
   U455 : AND2_X1 port map( A1 => N282, A2 => n1695, ZN => N299);
   U456 : AND2_X1 port map( A1 => N281, A2 => n1695, ZN => N300);
   U457 : AND2_X1 port map( A1 => N280, A2 => n1695, ZN => N301);
   U458 : AND2_X1 port map( A1 => N279, A2 => n1695, ZN => N302);
   U459 : AND2_X1 port map( A1 => N278, A2 => n1695, ZN => N303);
   U460 : AND2_X1 port map( A1 => N277, A2 => n1695, ZN => N304);
   U461 : AND2_X1 port map( A1 => N276, A2 => n1695, ZN => N305);
   U462 : AND2_X1 port map( A1 => N275, A2 => n1695, ZN => N306);
   U463 : AND2_X1 port map( A1 => N274, A2 => n1695, ZN => N307);
   U464 : AND2_X1 port map( A1 => N273, A2 => n1695, ZN => N308);
   U465 : AND2_X1 port map( A1 => N272, A2 => n1695, ZN => N309);
   U466 : AND2_X1 port map( A1 => N271, A2 => n1695, ZN => N310);
   U467 : AND2_X1 port map( A1 => N270, A2 => n1694, ZN => N311);
   U468 : AND2_X1 port map( A1 => N269, A2 => n1694, ZN => N312);
   U469 : AND2_X1 port map( A1 => N268, A2 => n1694, ZN => N313);
   U470 : AND2_X1 port map( A1 => N267, A2 => n1694, ZN => N314);
   U471 : AND2_X1 port map( A1 => N266, A2 => n1694, ZN => N315);
   U472 : AND2_X1 port map( A1 => N265, A2 => n1694, ZN => N316);
   U473 : AND2_X1 port map( A1 => N264, A2 => n1694, ZN => N317);
   U474 : AND2_X1 port map( A1 => N263, A2 => n1694, ZN => N318);
   U475 : AND2_X1 port map( A1 => N262, A2 => n1694, ZN => N319);
   U476 : AND2_X1 port map( A1 => N261, A2 => n1694, ZN => N320);
   U477 : AND2_X1 port map( A1 => N260, A2 => n1694, ZN => N321);
   U478 : AND2_X1 port map( A1 => N259, A2 => n1694, ZN => N322);
   U479 : AND2_X1 port map( A1 => N224, A2 => n1692, ZN => N225);
   U480 : AND2_X1 port map( A1 => N223, A2 => n1692, ZN => N226);
   U481 : AND2_X1 port map( A1 => N222, A2 => n1692, ZN => N227);
   U482 : AND2_X1 port map( A1 => N221, A2 => n1692, ZN => N228);
   U483 : AND2_X1 port map( A1 => N220, A2 => n1692, ZN => N229);
   U484 : AND2_X1 port map( A1 => N219, A2 => n1692, ZN => N230);
   U485 : AND2_X1 port map( A1 => N218, A2 => n1692, ZN => N231);
   U486 : AND2_X1 port map( A1 => N217, A2 => n1692, ZN => N232);
   U487 : AND2_X1 port map( A1 => N216, A2 => n1691, ZN => N233);
   U488 : AND2_X1 port map( A1 => N215, A2 => n1691, ZN => N234);
   U489 : AND2_X1 port map( A1 => N214, A2 => n1691, ZN => N235);
   U490 : AND2_X1 port map( A1 => N213, A2 => n1691, ZN => N236);
   U491 : AND2_X1 port map( A1 => N212, A2 => n1691, ZN => N237);
   U492 : AND2_X1 port map( A1 => N211, A2 => n1691, ZN => N238);
   U493 : AND2_X1 port map( A1 => N210, A2 => n1691, ZN => N239);
   U494 : AND2_X1 port map( A1 => N209, A2 => n1691, ZN => N240);
   U495 : AND2_X1 port map( A1 => N208, A2 => n1691, ZN => N241);
   U496 : AND2_X1 port map( A1 => N207, A2 => n1691, ZN => N242);
   U497 : AND2_X1 port map( A1 => N206, A2 => n1691, ZN => N243);
   U498 : AND2_X1 port map( A1 => N205, A2 => n1691, ZN => N244);
   U499 : AND2_X1 port map( A1 => N204, A2 => n1690, ZN => N245);
   U500 : AND2_X1 port map( A1 => N203, A2 => n1690, ZN => N246);
   U501 : AND2_X1 port map( A1 => N202, A2 => n1690, ZN => N247);
   U502 : AND2_X1 port map( A1 => N201, A2 => n1690, ZN => N248);
   U503 : AND2_X1 port map( A1 => N200, A2 => n1690, ZN => N249);
   U504 : AND2_X1 port map( A1 => N199, A2 => n1690, ZN => N250);
   U505 : AND2_X1 port map( A1 => N198, A2 => n1690, ZN => N251);
   U506 : AND2_X1 port map( A1 => N197, A2 => n1690, ZN => N252);
   U507 : AND2_X1 port map( A1 => N196, A2 => n1690, ZN => N253);
   U508 : AND2_X1 port map( A1 => N195, A2 => n1690, ZN => N254);
   U509 : AND2_X1 port map( A1 => N194, A2 => n1690, ZN => N255);
   U510 : AND2_X1 port map( A1 => N193, A2 => n1690, ZN => N256);
   U511 : BUF_X1 port map( A => n1678, Z => n1681);
   U512 : BUF_X1 port map( A => n1678, Z => n1680);
   U513 : BUF_X1 port map( A => n850, Z => n853);
   U514 : BUF_X1 port map( A => n850, Z => n852);
   U515 : BUF_X1 port map( A => n1697, Z => n1695);
   U516 : BUF_X1 port map( A => n1697, Z => n1694);
   U517 : BUF_X1 port map( A => n1693, Z => n1691);
   U518 : BUF_X1 port map( A => n1693, Z => n1690);
   U519 : BUF_X1 port map( A => n1674, Z => n1677);
   U520 : BUF_X1 port map( A => n1674, Z => n1676);
   U521 : BUF_X1 port map( A => n846, Z => n849);
   U522 : BUF_X1 port map( A => n846, Z => n848);
   U523 : BUF_X1 port map( A => n1686, Z => n1689);
   U524 : BUF_X1 port map( A => n1686, Z => n1688);
   U525 : BUF_X1 port map( A => n858, Z => n861);
   U526 : BUF_X1 port map( A => n858, Z => n860);
   U527 : BUF_X1 port map( A => n1682, Z => n1685);
   U528 : BUF_X1 port map( A => n854, Z => n857);
   U529 : BUF_X1 port map( A => n1682, Z => n1684);
   U530 : BUF_X1 port map( A => n854, Z => n856);
   U531 : BUF_X1 port map( A => n1678, Z => n1679);
   U532 : BUF_X1 port map( A => n850, Z => n851);
   U533 : BUF_X1 port map( A => n1674, Z => n1675);
   U534 : BUF_X1 port map( A => n846, Z => n847);
   U535 : BUF_X1 port map( A => n1697, Z => n1696);
   U536 : BUF_X1 port map( A => n1693, Z => n1692);
   U537 : BUF_X1 port map( A => n1686, Z => n1687);
   U538 : BUF_X1 port map( A => n858, Z => n859);
   U539 : BUF_X1 port map( A => n1682, Z => n1683);
   U540 : BUF_X1 port map( A => n854, Z => n855);
   U541 : NAND2_X1 port map( A1 => REGISTERS_2_31_port, A2 => n1659, ZN => 
                           n1525);
   U542 : NAND2_X1 port map( A1 => REGISTERS_2_31_port, A2 => n831, ZN => n697)
                           ;
   U543 : NAND2_X1 port map( A1 => REGISTERS_2_0_port, A2 => n1661, ZN => n874)
                           ;
   U544 : NAND2_X1 port map( A1 => REGISTERS_2_1_port, A2 => n1661, ZN => n895)
                           ;
   U545 : NAND2_X1 port map( A1 => REGISTERS_2_2_port, A2 => n1661, ZN => n916)
                           ;
   U546 : NAND2_X1 port map( A1 => REGISTERS_2_3_port, A2 => n1661, ZN => n937)
                           ;
   U547 : NAND2_X1 port map( A1 => REGISTERS_2_4_port, A2 => n1661, ZN => n958)
                           ;
   U548 : NAND2_X1 port map( A1 => REGISTERS_2_5_port, A2 => n1661, ZN => n979)
                           ;
   U549 : NAND2_X1 port map( A1 => REGISTERS_2_6_port, A2 => n1661, ZN => n1000
                           );
   U550 : NAND2_X1 port map( A1 => REGISTERS_2_7_port, A2 => n1661, ZN => n1021
                           );
   U551 : NAND2_X1 port map( A1 => REGISTERS_2_8_port, A2 => n1661, ZN => n1042
                           );
   U552 : NAND2_X1 port map( A1 => REGISTERS_2_9_port, A2 => n1661, ZN => n1063
                           );
   U553 : NAND2_X1 port map( A1 => REGISTERS_2_10_port, A2 => n1661, ZN => 
                           n1084);
   U554 : NAND2_X1 port map( A1 => REGISTERS_2_11_port, A2 => n1661, ZN => 
                           n1105);
   U555 : NAND2_X1 port map( A1 => REGISTERS_2_12_port, A2 => n1660, ZN => 
                           n1126);
   U556 : NAND2_X1 port map( A1 => REGISTERS_2_13_port, A2 => n1660, ZN => 
                           n1147);
   U557 : NAND2_X1 port map( A1 => REGISTERS_2_14_port, A2 => n1660, ZN => 
                           n1168);
   U558 : NAND2_X1 port map( A1 => REGISTERS_2_15_port, A2 => n1660, ZN => 
                           n1189);
   U559 : NAND2_X1 port map( A1 => REGISTERS_2_16_port, A2 => n1660, ZN => 
                           n1210);
   U560 : NAND2_X1 port map( A1 => REGISTERS_2_17_port, A2 => n1660, ZN => 
                           n1231);
   U561 : NAND2_X1 port map( A1 => REGISTERS_2_18_port, A2 => n1660, ZN => 
                           n1252);
   U562 : NAND2_X1 port map( A1 => REGISTERS_2_19_port, A2 => n1660, ZN => 
                           n1273);
   U563 : NAND2_X1 port map( A1 => REGISTERS_2_20_port, A2 => n1660, ZN => 
                           n1294);
   U564 : NAND2_X1 port map( A1 => REGISTERS_2_21_port, A2 => n1660, ZN => 
                           n1315);
   U565 : NAND2_X1 port map( A1 => REGISTERS_2_22_port, A2 => n1660, ZN => 
                           n1336);
   U566 : NAND2_X1 port map( A1 => REGISTERS_2_23_port, A2 => n1660, ZN => 
                           n1357);
   U567 : NAND2_X1 port map( A1 => REGISTERS_2_24_port, A2 => n1659, ZN => 
                           n1378);
   U568 : NAND2_X1 port map( A1 => REGISTERS_2_25_port, A2 => n1659, ZN => 
                           n1399);
   U569 : NAND2_X1 port map( A1 => REGISTERS_2_26_port, A2 => n1659, ZN => 
                           n1420);
   U570 : NAND2_X1 port map( A1 => REGISTERS_2_27_port, A2 => n1659, ZN => 
                           n1441);
   U571 : NAND2_X1 port map( A1 => REGISTERS_2_28_port, A2 => n1659, ZN => 
                           n1462);
   U572 : NAND2_X1 port map( A1 => REGISTERS_2_29_port, A2 => n1659, ZN => 
                           n1483);
   U573 : NAND2_X1 port map( A1 => REGISTERS_2_30_port, A2 => n1659, ZN => 
                           n1504);
   U574 : NAND2_X1 port map( A1 => REGISTERS_2_0_port, A2 => n833, ZN => n46);
   U575 : NAND2_X1 port map( A1 => REGISTERS_2_1_port, A2 => n833, ZN => n67);
   U576 : NAND2_X1 port map( A1 => REGISTERS_2_2_port, A2 => n833, ZN => n88);
   U577 : NAND2_X1 port map( A1 => REGISTERS_2_3_port, A2 => n833, ZN => n109);
   U578 : NAND2_X1 port map( A1 => REGISTERS_2_4_port, A2 => n833, ZN => 
                           n130_port);
   U579 : NAND2_X1 port map( A1 => REGISTERS_2_5_port, A2 => n833, ZN => 
                           n151_port);
   U580 : NAND2_X1 port map( A1 => REGISTERS_2_6_port, A2 => n833, ZN => n172);
   U581 : NAND2_X1 port map( A1 => REGISTERS_2_7_port, A2 => n833, ZN => 
                           n193_port);
   U582 : NAND2_X1 port map( A1 => REGISTERS_2_8_port, A2 => n833, ZN => 
                           n214_port);
   U583 : NAND2_X1 port map( A1 => REGISTERS_2_9_port, A2 => n833, ZN => 
                           n235_port);
   U584 : NAND2_X1 port map( A1 => REGISTERS_2_10_port, A2 => n833, ZN => 
                           n256_port);
   U585 : NAND2_X1 port map( A1 => REGISTERS_2_11_port, A2 => n833, ZN => 
                           n277_port);
   U586 : NAND2_X1 port map( A1 => REGISTERS_2_12_port, A2 => n832, ZN => 
                           n298_port);
   U587 : NAND2_X1 port map( A1 => REGISTERS_2_13_port, A2 => n832, ZN => 
                           n319_port);
   U588 : NAND2_X1 port map( A1 => REGISTERS_2_14_port, A2 => n832, ZN => 
                           n340_port);
   U589 : NAND2_X1 port map( A1 => REGISTERS_2_15_port, A2 => n832, ZN => n361)
                           ;
   U590 : NAND2_X1 port map( A1 => REGISTERS_2_16_port, A2 => n832, ZN => n382)
                           ;
   U591 : NAND2_X1 port map( A1 => REGISTERS_2_17_port, A2 => n832, ZN => n403)
                           ;
   U592 : NAND2_X1 port map( A1 => REGISTERS_2_18_port, A2 => n832, ZN => n424)
                           ;
   U593 : NAND2_X1 port map( A1 => REGISTERS_2_19_port, A2 => n832, ZN => n445)
                           ;
   U594 : NAND2_X1 port map( A1 => REGISTERS_2_20_port, A2 => n832, ZN => n466)
                           ;
   U595 : NAND2_X1 port map( A1 => REGISTERS_2_21_port, A2 => n832, ZN => n487)
                           ;
   U596 : NAND2_X1 port map( A1 => REGISTERS_2_22_port, A2 => n832, ZN => n508)
                           ;
   U597 : NAND2_X1 port map( A1 => REGISTERS_2_23_port, A2 => n832, ZN => n529)
                           ;
   U598 : NAND2_X1 port map( A1 => REGISTERS_2_24_port, A2 => n831, ZN => n550)
                           ;
   U599 : NAND2_X1 port map( A1 => REGISTERS_2_25_port, A2 => n831, ZN => n571)
                           ;
   U600 : NAND2_X1 port map( A1 => REGISTERS_2_26_port, A2 => n831, ZN => n592)
                           ;
   U601 : NAND2_X1 port map( A1 => REGISTERS_2_27_port, A2 => n831, ZN => n613)
                           ;
   U602 : NAND2_X1 port map( A1 => REGISTERS_2_28_port, A2 => n831, ZN => n634)
                           ;
   U603 : NAND2_X1 port map( A1 => REGISTERS_2_29_port, A2 => n831, ZN => n655)
                           ;
   U604 : NAND2_X1 port map( A1 => REGISTERS_2_30_port, A2 => n831, ZN => n676)
                           ;
   U605 : INV_X1 port map( A => ADD_RD2(0), ZN => n1544);
   U606 : INV_X1 port map( A => ADD_RD2(3), ZN => n1547);
   U607 : INV_X1 port map( A => ADD_RD2(2), ZN => n1546);
   U608 : INV_X1 port map( A => ADD_RD1(0), ZN => n716);
   U609 : INV_X1 port map( A => ADD_RD2(1), ZN => n1545);
   U610 : AND3_X1 port map( A1 => ENABLE, A2 => n1, A3 => WR, ZN => n17);
   U611 : INV_X1 port map( A => ADD_RD1(1), ZN => n717);
   U612 : INV_X1 port map( A => ADD_RD1(3), ZN => n719);
   U613 : INV_X1 port map( A => ADD_RD1(2), ZN => n718);
   U614 : INV_X1 port map( A => ADD_WR(0), ZN => n1796);
   U615 : INV_X1 port map( A => ADD_WR(2), ZN => n1794);
   U616 : INV_X1 port map( A => ADD_WR(1), ZN => n1795);
   U617 : AND2_X1 port map( A1 => RD2, A2 => n23, ZN => n22);
   U618 : OR4_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => ADD_RD2(2)
                           , A4 => n24, ZN => n23);
   U619 : OR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), ZN => n24);
   U620 : AND2_X1 port map( A1 => RD1, A2 => n26, ZN => n25);
   U621 : OR4_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => ADD_RD1(2)
                           , A4 => n27, ZN => n26);
   U622 : OR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n27);
   U623 : INV_X1 port map( A => ADD_WR(4), ZN => n1792);
   U624 : INV_X1 port map( A => ADD_WR(3), ZN => n1793);
   U625 : INV_X1 port map( A => CLK, ZN => n1);
   U626 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n719, ZN => n714);
   U627 : NOR2_X1 port map( A1 => n718, A2 => ADD_RD1(1), ZN => n34);
   U628 : NOR2_X1 port map( A1 => n718, A2 => n717, ZN => n35);
   U629 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n753, B1 => 
                           REGISTERS_23_0_port, B2 => n736, ZN => n41);
   U630 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n36);
   U631 : NOR2_X1 port map( A1 => n717, A2 => ADD_RD1(2), ZN => n37);
   U632 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n787, B1 => 
                           REGISTERS_19_0_port, B2 => n770, ZN => n40);
   U633 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n821, B1 => 
                           REGISTERS_22_0_port, B2 => n804, ZN => n39);
   U634 : AND2_X1 port map( A1 => n36, A2 => n716, ZN => n702);
   U635 : AND2_X1 port map( A1 => n37, A2 => n716, ZN => n701);
   U636 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n845, B1 => 
                           REGISTERS_18_0_port, B2 => n831, ZN => n38);
   U637 : AND4_X1 port map( A1 => n41, A2 => n40, A3 => n39, A4 => n38, ZN => 
                           n58);
   U638 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n712);
   U639 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n753, B1 => 
                           REGISTERS_31_0_port, B2 => n736, ZN => n45);
   U640 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n787, B1 => 
                           REGISTERS_27_0_port, B2 => n770, ZN => n44);
   U641 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n821, B1 => 
                           REGISTERS_30_0_port, B2 => n804, ZN => n43);
   U642 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n845, B1 => 
                           REGISTERS_26_0_port, B2 => n831, ZN => n42);
   U643 : AND4_X1 port map( A1 => n45, A2 => n44, A3 => n43, A4 => n42, ZN => 
                           n57);
   U644 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n753, B1 => 
                           REGISTERS_7_0_port, B2 => n736, ZN => n49);
   U645 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n787, B1 => 
                           REGISTERS_3_0_port, B2 => n770, ZN => n48);
   U646 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n821, B1 => 
                           REGISTERS_6_0_port, B2 => n804, ZN => n47);
   U647 : NAND4_X1 port map( A1 => n49, A2 => n48, A3 => n47, A4 => n46, ZN => 
                           n55);
   U648 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n710);
   U649 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n753, B1 => 
                           REGISTERS_15_0_port, B2 => n736, ZN => n53);
   U650 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n787, B1 => 
                           REGISTERS_11_0_port, B2 => n770, ZN => n52);
   U651 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n821, B1 => 
                           REGISTERS_14_0_port, B2 => n804, ZN => n51);
   U652 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n845, B1 => 
                           REGISTERS_10_0_port, B2 => n831, ZN => n50);
   U653 : NAND4_X1 port map( A1 => n53, A2 => n52, A3 => n51, A4 => n50, ZN => 
                           n54);
   U654 : NOR2_X1 port map( A1 => n719, A2 => ADD_RD1(4), ZN => n708);
   U655 : AOI22_X1 port map( A1 => n55, A2 => n853, B1 => n54, B2 => n849, ZN 
                           => n56);
   U656 : OAI221_X1 port map( B1 => n861, B2 => n58, C1 => n855, C2 => n57, A 
                           => n56, ZN => N224);
   U657 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n753, B1 => 
                           REGISTERS_23_1_port, B2 => n736, ZN => n62);
   U658 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n787, B1 => 
                           REGISTERS_19_1_port, B2 => n770, ZN => n61);
   U659 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n821, B1 => 
                           REGISTERS_22_1_port, B2 => n804, ZN => n60);
   U660 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n845, B1 => 
                           REGISTERS_18_1_port, B2 => n831, ZN => n59);
   U661 : AND4_X1 port map( A1 => n62, A2 => n61, A3 => n60, A4 => n59, ZN => 
                           n79);
   U662 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n753, B1 => 
                           REGISTERS_31_1_port, B2 => n736, ZN => n66);
   U663 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n787, B1 => 
                           REGISTERS_27_1_port, B2 => n770, ZN => n65);
   U664 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n821, B1 => 
                           REGISTERS_30_1_port, B2 => n804, ZN => n64);
   U665 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n845, B1 => 
                           REGISTERS_26_1_port, B2 => n831, ZN => n63);
   U666 : AND4_X1 port map( A1 => n66, A2 => n65, A3 => n64, A4 => n63, ZN => 
                           n78);
   U667 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n753, B1 => 
                           REGISTERS_7_1_port, B2 => n736, ZN => n70);
   U668 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n787, B1 => 
                           REGISTERS_3_1_port, B2 => n770, ZN => n69);
   U669 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n821, B1 => 
                           REGISTERS_6_1_port, B2 => n804, ZN => n68);
   U670 : NAND4_X1 port map( A1 => n70, A2 => n69, A3 => n68, A4 => n67, ZN => 
                           n76);
   U671 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n753, B1 => 
                           REGISTERS_15_1_port, B2 => n736, ZN => n74);
   U672 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n787, B1 => 
                           REGISTERS_11_1_port, B2 => n770, ZN => n73);
   U673 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n821, B1 => 
                           REGISTERS_14_1_port, B2 => n804, ZN => n72);
   U674 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n845, B1 => 
                           REGISTERS_10_1_port, B2 => n831, ZN => n71);
   U675 : NAND4_X1 port map( A1 => n74, A2 => n73, A3 => n72, A4 => n71, ZN => 
                           n75);
   U676 : AOI22_X1 port map( A1 => n76, A2 => n853, B1 => n75, B2 => n849, ZN 
                           => n77);
   U677 : OAI221_X1 port map( B1 => n861, B2 => n79, C1 => n855, C2 => n78, A 
                           => n77, ZN => N223);
   U678 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n753, B1 => 
                           REGISTERS_23_2_port, B2 => n736, ZN => n83);
   U679 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n787, B1 => 
                           REGISTERS_19_2_port, B2 => n770, ZN => n82);
   U680 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n821, B1 => 
                           REGISTERS_22_2_port, B2 => n804, ZN => n81);
   U681 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n845, B1 => 
                           REGISTERS_18_2_port, B2 => n831, ZN => n80);
   U682 : AND4_X1 port map( A1 => n83, A2 => n82, A3 => n81, A4 => n80, ZN => 
                           n100);
   U683 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n753, B1 => 
                           REGISTERS_31_2_port, B2 => n736, ZN => n87);
   U684 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n787, B1 => 
                           REGISTERS_27_2_port, B2 => n770, ZN => n86);
   U685 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n821, B1 => 
                           REGISTERS_30_2_port, B2 => n804, ZN => n85);
   U686 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n845, B1 => 
                           REGISTERS_26_2_port, B2 => n830, ZN => n84);
   U687 : AND4_X1 port map( A1 => n87, A2 => n86, A3 => n85, A4 => n84, ZN => 
                           n99);
   U688 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n753, B1 => 
                           REGISTERS_7_2_port, B2 => n736, ZN => n91);
   U689 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n787, B1 => 
                           REGISTERS_3_2_port, B2 => n770, ZN => n90);
   U690 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n821, B1 => 
                           REGISTERS_6_2_port, B2 => n804, ZN => n89);
   U691 : NAND4_X1 port map( A1 => n91, A2 => n90, A3 => n89, A4 => n88, ZN => 
                           n97);
   U692 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n753, B1 => 
                           REGISTERS_15_2_port, B2 => n736, ZN => n95);
   U693 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n787, B1 => 
                           REGISTERS_11_2_port, B2 => n770, ZN => n94);
   U694 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n821, B1 => 
                           REGISTERS_14_2_port, B2 => n804, ZN => n93);
   U695 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n845, B1 => 
                           REGISTERS_10_2_port, B2 => n830, ZN => n92);
   U696 : NAND4_X1 port map( A1 => n95, A2 => n94, A3 => n93, A4 => n92, ZN => 
                           n96);
   U697 : AOI22_X1 port map( A1 => n97, A2 => n853, B1 => n96, B2 => n849, ZN 
                           => n98);
   U698 : OAI221_X1 port map( B1 => n861, B2 => n100, C1 => n855, C2 => n99, A 
                           => n98, ZN => N222);
   U699 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n752, B1 => 
                           REGISTERS_23_3_port, B2 => n735, ZN => n104);
   U700 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n786, B1 => 
                           REGISTERS_19_3_port, B2 => n769, ZN => n103);
   U701 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n820, B1 => 
                           REGISTERS_22_3_port, B2 => n803, ZN => n102);
   U702 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n845, B1 => 
                           REGISTERS_18_3_port, B2 => n830, ZN => n101);
   U703 : AND4_X1 port map( A1 => n104, A2 => n103, A3 => n102, A4 => n101, ZN 
                           => n121);
   U704 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n752, B1 => 
                           REGISTERS_31_3_port, B2 => n735, ZN => n108);
   U705 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n786, B1 => 
                           REGISTERS_27_3_port, B2 => n769, ZN => n107);
   U706 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n820, B1 => 
                           REGISTERS_30_3_port, B2 => n803, ZN => n106);
   U707 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n845, B1 => 
                           REGISTERS_26_3_port, B2 => n830, ZN => n105);
   U708 : AND4_X1 port map( A1 => n108, A2 => n107, A3 => n106, A4 => n105, ZN 
                           => n120);
   U709 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n752, B1 => 
                           REGISTERS_7_3_port, B2 => n735, ZN => n112);
   U710 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n786, B1 => 
                           REGISTERS_3_3_port, B2 => n769, ZN => n111);
   U711 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n820, B1 => 
                           REGISTERS_6_3_port, B2 => n803, ZN => n110);
   U712 : NAND4_X1 port map( A1 => n112, A2 => n111, A3 => n110, A4 => n109, ZN
                           => n118);
   U713 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n752, B1 => 
                           REGISTERS_15_3_port, B2 => n735, ZN => n116);
   U714 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n786, B1 => 
                           REGISTERS_11_3_port, B2 => n769, ZN => n115);
   U715 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n820, B1 => 
                           REGISTERS_14_3_port, B2 => n803, ZN => n114);
   U716 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n845, B1 => 
                           REGISTERS_10_3_port, B2 => n830, ZN => n113);
   U717 : NAND4_X1 port map( A1 => n116, A2 => n115, A3 => n114, A4 => n113, ZN
                           => n117);
   U718 : AOI22_X1 port map( A1 => n118, A2 => n853, B1 => n117, B2 => n849, ZN
                           => n119);
   U719 : OAI221_X1 port map( B1 => n861, B2 => n121, C1 => n855, C2 => n120, A
                           => n119, ZN => N221);
   U720 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n752, B1 => 
                           REGISTERS_23_4_port, B2 => n735, ZN => n125);
   U721 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n786, B1 => 
                           REGISTERS_19_4_port, B2 => n769, ZN => n124);
   U722 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n820, B1 => 
                           REGISTERS_22_4_port, B2 => n803, ZN => n123);
   U723 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n844, B1 => 
                           REGISTERS_18_4_port, B2 => n830, ZN => n122);
   U724 : AND4_X1 port map( A1 => n125, A2 => n124, A3 => n123, A4 => n122, ZN 
                           => n142_port);
   U725 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n752, B1 => 
                           REGISTERS_31_4_port, B2 => n735, ZN => n129_port);
   U726 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n786, B1 => 
                           REGISTERS_27_4_port, B2 => n769, ZN => n128_port);
   U727 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n820, B1 => 
                           REGISTERS_30_4_port, B2 => n803, ZN => n127);
   U728 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n844, B1 => 
                           REGISTERS_26_4_port, B2 => n830, ZN => n126);
   U729 : AND4_X1 port map( A1 => n129_port, A2 => n128_port, A3 => n127, A4 =>
                           n126, ZN => n141_port);
   U730 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n752, B1 => 
                           REGISTERS_7_4_port, B2 => n735, ZN => n133_port);
   U731 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n786, B1 => 
                           REGISTERS_3_4_port, B2 => n769, ZN => n132_port);
   U732 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n820, B1 => 
                           REGISTERS_6_4_port, B2 => n803, ZN => n131_port);
   U733 : NAND4_X1 port map( A1 => n133_port, A2 => n132_port, A3 => n131_port,
                           A4 => n130_port, ZN => n139_port);
   U734 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n752, B1 => 
                           REGISTERS_15_4_port, B2 => n735, ZN => n137_port);
   U735 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n786, B1 => 
                           REGISTERS_11_4_port, B2 => n769, ZN => n136_port);
   U736 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n820, B1 => 
                           REGISTERS_14_4_port, B2 => n803, ZN => n135_port);
   U737 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n844, B1 => 
                           REGISTERS_10_4_port, B2 => n830, ZN => n134_port);
   U738 : NAND4_X1 port map( A1 => n137_port, A2 => n136_port, A3 => n135_port,
                           A4 => n134_port, ZN => n138_port);
   U739 : AOI22_X1 port map( A1 => n139_port, A2 => n853, B1 => n138_port, B2 
                           => n849, ZN => n140_port);
   U740 : OAI221_X1 port map( B1 => n861, B2 => n142_port, C1 => n855, C2 => 
                           n141_port, A => n140_port, ZN => N220);
   U741 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n752, B1 => 
                           REGISTERS_23_5_port, B2 => n735, ZN => n146_port);
   U742 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n786, B1 => 
                           REGISTERS_19_5_port, B2 => n769, ZN => n145_port);
   U743 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n820, B1 => 
                           REGISTERS_22_5_port, B2 => n803, ZN => n144_port);
   U744 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n844, B1 => 
                           REGISTERS_18_5_port, B2 => n830, ZN => n143_port);
   U745 : AND4_X1 port map( A1 => n146_port, A2 => n145_port, A3 => n144_port, 
                           A4 => n143_port, ZN => n163);
   U746 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n752, B1 => 
                           REGISTERS_31_5_port, B2 => n735, ZN => n150_port);
   U747 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n786, B1 => 
                           REGISTERS_27_5_port, B2 => n769, ZN => n149_port);
   U748 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n820, B1 => 
                           REGISTERS_30_5_port, B2 => n803, ZN => n148_port);
   U749 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n844, B1 => 
                           REGISTERS_26_5_port, B2 => n830, ZN => n147_port);
   U750 : AND4_X1 port map( A1 => n150_port, A2 => n149_port, A3 => n148_port, 
                           A4 => n147_port, ZN => n162);
   U751 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n752, B1 => 
                           REGISTERS_7_5_port, B2 => n735, ZN => n154_port);
   U752 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n786, B1 => 
                           REGISTERS_3_5_port, B2 => n769, ZN => n153_port);
   U753 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n820, B1 => 
                           REGISTERS_6_5_port, B2 => n803, ZN => n152_port);
   U754 : NAND4_X1 port map( A1 => n154_port, A2 => n153_port, A3 => n152_port,
                           A4 => n151_port, ZN => n160);
   U755 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n752, B1 => 
                           REGISTERS_15_5_port, B2 => n735, ZN => n158_port);
   U756 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n786, B1 => 
                           REGISTERS_11_5_port, B2 => n769, ZN => n157_port);
   U757 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n820, B1 => 
                           REGISTERS_14_5_port, B2 => n803, ZN => n156_port);
   U758 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n844, B1 => 
                           REGISTERS_10_5_port, B2 => n830, ZN => n155_port);
   U759 : NAND4_X1 port map( A1 => n158_port, A2 => n157_port, A3 => n156_port,
                           A4 => n155_port, ZN => n159_port);
   U760 : AOI22_X1 port map( A1 => n160, A2 => n853, B1 => n159_port, B2 => 
                           n849, ZN => n161);
   U761 : OAI221_X1 port map( B1 => n861, B2 => n163, C1 => n855, C2 => n162, A
                           => n161, ZN => N219);
   U762 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n751, B1 => 
                           REGISTERS_23_6_port, B2 => n734, ZN => n167);
   U763 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n785, B1 => 
                           REGISTERS_19_6_port, B2 => n768, ZN => n166);
   U764 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n819, B1 => 
                           REGISTERS_22_6_port, B2 => n802, ZN => n165);
   U765 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n844, B1 => 
                           REGISTERS_18_6_port, B2 => n830, ZN => n164);
   U766 : AND4_X1 port map( A1 => n167, A2 => n166, A3 => n165, A4 => n164, ZN 
                           => n184);
   U767 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n751, B1 => 
                           REGISTERS_31_6_port, B2 => n734, ZN => n171);
   U768 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n785, B1 => 
                           REGISTERS_27_6_port, B2 => n768, ZN => n170);
   U769 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n819, B1 => 
                           REGISTERS_30_6_port, B2 => n802, ZN => n169);
   U770 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n844, B1 => 
                           REGISTERS_26_6_port, B2 => n830, ZN => n168);
   U771 : AND4_X1 port map( A1 => n171, A2 => n170, A3 => n169, A4 => n168, ZN 
                           => n183);
   U772 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n751, B1 => 
                           REGISTERS_7_6_port, B2 => n734, ZN => n175);
   U773 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n785, B1 => 
                           REGISTERS_3_6_port, B2 => n768, ZN => n174);
   U774 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n819, B1 => 
                           REGISTERS_6_6_port, B2 => n802, ZN => n173);
   U775 : NAND4_X1 port map( A1 => n175, A2 => n174, A3 => n173, A4 => n172, ZN
                           => n181);
   U776 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n751, B1 => 
                           REGISTERS_15_6_port, B2 => n734, ZN => n179);
   U777 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n785, B1 => 
                           REGISTERS_11_6_port, B2 => n768, ZN => n178);
   U778 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n819, B1 => 
                           REGISTERS_14_6_port, B2 => n802, ZN => n177);
   U779 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n844, B1 => 
                           REGISTERS_10_6_port, B2 => n830, ZN => n176);
   U780 : NAND4_X1 port map( A1 => n179, A2 => n178, A3 => n177, A4 => n176, ZN
                           => n180);
   U781 : AOI22_X1 port map( A1 => n181, A2 => n853, B1 => n180, B2 => n849, ZN
                           => n182);
   U782 : OAI221_X1 port map( B1 => n861, B2 => n184, C1 => n855, C2 => n183, A
                           => n182, ZN => N218);
   U783 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n751, B1 => 
                           REGISTERS_23_7_port, B2 => n734, ZN => n188);
   U784 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n785, B1 => 
                           REGISTERS_19_7_port, B2 => n768, ZN => n187);
   U785 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n819, B1 => 
                           REGISTERS_22_7_port, B2 => n802, ZN => n186);
   U786 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n844, B1 => 
                           REGISTERS_18_7_port, B2 => n830, ZN => n185);
   U787 : AND4_X1 port map( A1 => n188, A2 => n187, A3 => n186, A4 => n185, ZN 
                           => n205_port);
   U788 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n751, B1 => 
                           REGISTERS_31_7_port, B2 => n734, ZN => n192);
   U789 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n785, B1 => 
                           REGISTERS_27_7_port, B2 => n768, ZN => n191);
   U790 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n819, B1 => 
                           REGISTERS_30_7_port, B2 => n802, ZN => n190);
   U791 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n844, B1 => 
                           REGISTERS_26_7_port, B2 => n830, ZN => n189);
   U792 : AND4_X1 port map( A1 => n192, A2 => n191, A3 => n190, A4 => n189, ZN 
                           => n204_port);
   U793 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n751, B1 => 
                           REGISTERS_7_7_port, B2 => n734, ZN => n196_port);
   U794 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n785, B1 => 
                           REGISTERS_3_7_port, B2 => n768, ZN => n195_port);
   U795 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n819, B1 => 
                           REGISTERS_6_7_port, B2 => n802, ZN => n194_port);
   U796 : NAND4_X1 port map( A1 => n196_port, A2 => n195_port, A3 => n194_port,
                           A4 => n193_port, ZN => n202_port);
   U797 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n751, B1 => 
                           REGISTERS_15_7_port, B2 => n734, ZN => n200_port);
   U798 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n785, B1 => 
                           REGISTERS_11_7_port, B2 => n768, ZN => n199_port);
   U799 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n819, B1 => 
                           REGISTERS_14_7_port, B2 => n802, ZN => n198_port);
   U800 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n844, B1 => 
                           REGISTERS_10_7_port, B2 => n830, ZN => n197_port);
   U801 : NAND4_X1 port map( A1 => n200_port, A2 => n199_port, A3 => n198_port,
                           A4 => n197_port, ZN => n201_port);
   U802 : AOI22_X1 port map( A1 => n202_port, A2 => n853, B1 => n201_port, B2 
                           => n849, ZN => n203_port);
   U803 : OAI221_X1 port map( B1 => n861, B2 => n205_port, C1 => n855, C2 => 
                           n204_port, A => n203_port, ZN => N217);
   U804 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n751, B1 => 
                           REGISTERS_23_8_port, B2 => n734, ZN => n209_port);
   U805 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n785, B1 => 
                           REGISTERS_19_8_port, B2 => n768, ZN => n208_port);
   U806 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n819, B1 => 
                           REGISTERS_22_8_port, B2 => n802, ZN => n207_port);
   U807 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n843, B1 => 
                           REGISTERS_18_8_port, B2 => n830, ZN => n206_port);
   U808 : AND4_X1 port map( A1 => n209_port, A2 => n208_port, A3 => n207_port, 
                           A4 => n206_port, ZN => n226_port);
   U809 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n751, B1 => 
                           REGISTERS_31_8_port, B2 => n734, ZN => n213_port);
   U810 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n785, B1 => 
                           REGISTERS_27_8_port, B2 => n768, ZN => n212_port);
   U811 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n819, B1 => 
                           REGISTERS_30_8_port, B2 => n802, ZN => n211_port);
   U812 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n843, B1 => 
                           REGISTERS_26_8_port, B2 => n830, ZN => n210_port);
   U813 : AND4_X1 port map( A1 => n213_port, A2 => n212_port, A3 => n211_port, 
                           A4 => n210_port, ZN => n225_port);
   U814 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n751, B1 => 
                           REGISTERS_7_8_port, B2 => n734, ZN => n217_port);
   U815 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n785, B1 => 
                           REGISTERS_3_8_port, B2 => n768, ZN => n216_port);
   U816 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n819, B1 => 
                           REGISTERS_6_8_port, B2 => n802, ZN => n215_port);
   U817 : NAND4_X1 port map( A1 => n217_port, A2 => n216_port, A3 => n215_port,
                           A4 => n214_port, ZN => n223_port);
   U818 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n751, B1 => 
                           REGISTERS_15_8_port, B2 => n734, ZN => n221_port);
   U819 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n785, B1 => 
                           REGISTERS_11_8_port, B2 => n768, ZN => n220_port);
   U820 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n819, B1 => 
                           REGISTERS_14_8_port, B2 => n802, ZN => n219_port);
   U821 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n843, B1 => 
                           REGISTERS_10_8_port, B2 => n830, ZN => n218_port);
   U822 : NAND4_X1 port map( A1 => n221_port, A2 => n220_port, A3 => n219_port,
                           A4 => n218_port, ZN => n222_port);
   U823 : AOI22_X1 port map( A1 => n223_port, A2 => n853, B1 => n222_port, B2 
                           => n849, ZN => n224_port);
   U824 : OAI221_X1 port map( B1 => n861, B2 => n226_port, C1 => n856, C2 => 
                           n225_port, A => n224_port, ZN => N216);
   U825 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n750, B1 => 
                           REGISTERS_23_9_port, B2 => n733, ZN => n230_port);
   U826 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n784, B1 => 
                           REGISTERS_19_9_port, B2 => n767, ZN => n229_port);
   U827 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n818, B1 => 
                           REGISTERS_22_9_port, B2 => n801, ZN => n228_port);
   U828 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n843, B1 => 
                           REGISTERS_18_9_port, B2 => n829, ZN => n227_port);
   U829 : AND4_X1 port map( A1 => n230_port, A2 => n229_port, A3 => n228_port, 
                           A4 => n227_port, ZN => n247_port);
   U830 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n750, B1 => 
                           REGISTERS_31_9_port, B2 => n733, ZN => n234_port);
   U831 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n784, B1 => 
                           REGISTERS_27_9_port, B2 => n767, ZN => n233_port);
   U832 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n818, B1 => 
                           REGISTERS_30_9_port, B2 => n801, ZN => n232_port);
   U833 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n843, B1 => 
                           REGISTERS_26_9_port, B2 => n829, ZN => n231_port);
   U834 : AND4_X1 port map( A1 => n234_port, A2 => n233_port, A3 => n232_port, 
                           A4 => n231_port, ZN => n246_port);
   U835 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n750, B1 => 
                           REGISTERS_7_9_port, B2 => n733, ZN => n238_port);
   U836 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n784, B1 => 
                           REGISTERS_3_9_port, B2 => n767, ZN => n237_port);
   U837 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n818, B1 => 
                           REGISTERS_6_9_port, B2 => n801, ZN => n236_port);
   U838 : NAND4_X1 port map( A1 => n238_port, A2 => n237_port, A3 => n236_port,
                           A4 => n235_port, ZN => n244_port);
   U839 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n750, B1 => 
                           REGISTERS_15_9_port, B2 => n733, ZN => n242_port);
   U840 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n784, B1 => 
                           REGISTERS_11_9_port, B2 => n767, ZN => n241_port);
   U841 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n818, B1 => 
                           REGISTERS_14_9_port, B2 => n801, ZN => n240_port);
   U842 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n843, B1 => 
                           REGISTERS_10_9_port, B2 => n829, ZN => n239_port);
   U843 : NAND4_X1 port map( A1 => n242_port, A2 => n241_port, A3 => n240_port,
                           A4 => n239_port, ZN => n243_port);
   U844 : AOI22_X1 port map( A1 => n244_port, A2 => n853, B1 => n243_port, B2 
                           => n849, ZN => n245_port);
   U845 : OAI221_X1 port map( B1 => n861, B2 => n247_port, C1 => n856, C2 => 
                           n246_port, A => n245_port, ZN => N215);
   U846 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n750, B1 => 
                           REGISTERS_23_10_port, B2 => n733, ZN => n251_port);
   U847 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n784, B1 => 
                           REGISTERS_19_10_port, B2 => n767, ZN => n250_port);
   U848 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n818, B1 => 
                           REGISTERS_22_10_port, B2 => n801, ZN => n249_port);
   U849 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n843, B1 => 
                           REGISTERS_18_10_port, B2 => n829, ZN => n248_port);
   U850 : AND4_X1 port map( A1 => n251_port, A2 => n250_port, A3 => n249_port, 
                           A4 => n248_port, ZN => n268_port);
   U851 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n750, B1 => 
                           REGISTERS_31_10_port, B2 => n733, ZN => n255_port);
   U852 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n784, B1 => 
                           REGISTERS_27_10_port, B2 => n767, ZN => n254_port);
   U853 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n818, B1 => 
                           REGISTERS_30_10_port, B2 => n801, ZN => n253_port);
   U854 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n843, B1 => 
                           REGISTERS_26_10_port, B2 => n829, ZN => n252_port);
   U855 : AND4_X1 port map( A1 => n255_port, A2 => n254_port, A3 => n253_port, 
                           A4 => n252_port, ZN => n267_port);
   U856 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n750, B1 => 
                           REGISTERS_7_10_port, B2 => n733, ZN => n259_port);
   U857 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n784, B1 => 
                           REGISTERS_3_10_port, B2 => n767, ZN => n258);
   U858 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n818, B1 => 
                           REGISTERS_6_10_port, B2 => n801, ZN => n257);
   U859 : NAND4_X1 port map( A1 => n259_port, A2 => n258, A3 => n257, A4 => 
                           n256_port, ZN => n265_port);
   U860 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n750, B1 => 
                           REGISTERS_15_10_port, B2 => n733, ZN => n263_port);
   U861 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n784, B1 => 
                           REGISTERS_11_10_port, B2 => n767, ZN => n262_port);
   U862 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n818, B1 => 
                           REGISTERS_14_10_port, B2 => n801, ZN => n261_port);
   U863 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n843, B1 => 
                           REGISTERS_10_10_port, B2 => n829, ZN => n260_port);
   U864 : NAND4_X1 port map( A1 => n263_port, A2 => n262_port, A3 => n261_port,
                           A4 => n260_port, ZN => n264_port);
   U865 : AOI22_X1 port map( A1 => n265_port, A2 => n853, B1 => n264_port, B2 
                           => n849, ZN => n266_port);
   U866 : OAI221_X1 port map( B1 => n861, B2 => n268_port, C1 => n856, C2 => 
                           n267_port, A => n266_port, ZN => N214);
   U867 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n750, B1 => 
                           REGISTERS_23_11_port, B2 => n733, ZN => n272_port);
   U868 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n784, B1 => 
                           REGISTERS_19_11_port, B2 => n767, ZN => n271_port);
   U869 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n818, B1 => 
                           REGISTERS_22_11_port, B2 => n801, ZN => n270_port);
   U870 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n843, B1 => 
                           REGISTERS_18_11_port, B2 => n829, ZN => n269_port);
   U871 : AND4_X1 port map( A1 => n272_port, A2 => n271_port, A3 => n270_port, 
                           A4 => n269_port, ZN => n289_port);
   U872 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n750, B1 => 
                           REGISTERS_31_11_port, B2 => n733, ZN => n276_port);
   U873 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n784, B1 => 
                           REGISTERS_27_11_port, B2 => n767, ZN => n275_port);
   U874 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n818, B1 => 
                           REGISTERS_30_11_port, B2 => n801, ZN => n274_port);
   U875 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n843, B1 => 
                           REGISTERS_26_11_port, B2 => n829, ZN => n273_port);
   U876 : AND4_X1 port map( A1 => n276_port, A2 => n275_port, A3 => n274_port, 
                           A4 => n273_port, ZN => n288_port);
   U877 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n750, B1 => 
                           REGISTERS_7_11_port, B2 => n733, ZN => n280_port);
   U878 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n784, B1 => 
                           REGISTERS_3_11_port, B2 => n767, ZN => n279_port);
   U879 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n818, B1 => 
                           REGISTERS_6_11_port, B2 => n801, ZN => n278_port);
   U880 : NAND4_X1 port map( A1 => n280_port, A2 => n279_port, A3 => n278_port,
                           A4 => n277_port, ZN => n286_port);
   U881 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n750, B1 => 
                           REGISTERS_15_11_port, B2 => n733, ZN => n284_port);
   U882 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n784, B1 => 
                           REGISTERS_11_11_port, B2 => n767, ZN => n283_port);
   U883 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n818, B1 => 
                           REGISTERS_14_11_port, B2 => n801, ZN => n282_port);
   U884 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n843, B1 => 
                           REGISTERS_10_11_port, B2 => n829, ZN => n281_port);
   U885 : NAND4_X1 port map( A1 => n284_port, A2 => n283_port, A3 => n282_port,
                           A4 => n281_port, ZN => n285_port);
   U886 : AOI22_X1 port map( A1 => n286_port, A2 => n853, B1 => n285_port, B2 
                           => n849, ZN => n287_port);
   U887 : OAI221_X1 port map( B1 => n861, B2 => n289_port, C1 => n856, C2 => 
                           n288_port, A => n287_port, ZN => N213);
   U888 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n749, B1 => 
                           REGISTERS_23_12_port, B2 => n732, ZN => n293_port);
   U889 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n783, B1 => 
                           REGISTERS_19_12_port, B2 => n766, ZN => n292_port);
   U890 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n817, B1 => 
                           REGISTERS_22_12_port, B2 => n800, ZN => n291_port);
   U891 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n842, B1 => 
                           REGISTERS_18_12_port, B2 => n829, ZN => n290_port);
   U892 : AND4_X1 port map( A1 => n293_port, A2 => n292_port, A3 => n291_port, 
                           A4 => n290_port, ZN => n310_port);
   U893 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n749, B1 => 
                           REGISTERS_31_12_port, B2 => n732, ZN => n297_port);
   U894 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n783, B1 => 
                           REGISTERS_27_12_port, B2 => n766, ZN => n296_port);
   U895 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n817, B1 => 
                           REGISTERS_30_12_port, B2 => n800, ZN => n295_port);
   U896 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n842, B1 => 
                           REGISTERS_26_12_port, B2 => n829, ZN => n294_port);
   U897 : AND4_X1 port map( A1 => n297_port, A2 => n296_port, A3 => n295_port, 
                           A4 => n294_port, ZN => n309_port);
   U898 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n749, B1 => 
                           REGISTERS_7_12_port, B2 => n732, ZN => n301_port);
   U899 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n783, B1 => 
                           REGISTERS_3_12_port, B2 => n766, ZN => n300_port);
   U900 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n817, B1 => 
                           REGISTERS_6_12_port, B2 => n800, ZN => n299_port);
   U901 : NAND4_X1 port map( A1 => n301_port, A2 => n300_port, A3 => n299_port,
                           A4 => n298_port, ZN => n307_port);
   U902 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n749, B1 => 
                           REGISTERS_15_12_port, B2 => n732, ZN => n305_port);
   U903 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n783, B1 => 
                           REGISTERS_11_12_port, B2 => n766, ZN => n304_port);
   U904 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n817, B1 => 
                           REGISTERS_14_12_port, B2 => n800, ZN => n303_port);
   U905 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n842, B1 => 
                           REGISTERS_10_12_port, B2 => n829, ZN => n302_port);
   U906 : NAND4_X1 port map( A1 => n305_port, A2 => n304_port, A3 => n303_port,
                           A4 => n302_port, ZN => n306_port);
   U907 : AOI22_X1 port map( A1 => n307_port, A2 => n852, B1 => n306_port, B2 
                           => n848, ZN => n308_port);
   U908 : OAI221_X1 port map( B1 => n860, B2 => n310_port, C1 => n856, C2 => 
                           n309_port, A => n308_port, ZN => N212);
   U909 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n749, B1 => 
                           REGISTERS_23_13_port, B2 => n732, ZN => n314_port);
   U910 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n783, B1 => 
                           REGISTERS_19_13_port, B2 => n766, ZN => n313_port);
   U911 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n817, B1 => 
                           REGISTERS_22_13_port, B2 => n800, ZN => n312_port);
   U912 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n842, B1 => 
                           REGISTERS_18_13_port, B2 => n829, ZN => n311_port);
   U913 : AND4_X1 port map( A1 => n314_port, A2 => n313_port, A3 => n312_port, 
                           A4 => n311_port, ZN => n331_port);
   U914 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n749, B1 => 
                           REGISTERS_31_13_port, B2 => n732, ZN => n318_port);
   U915 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n783, B1 => 
                           REGISTERS_27_13_port, B2 => n766, ZN => n317_port);
   U916 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n817, B1 => 
                           REGISTERS_30_13_port, B2 => n800, ZN => n316_port);
   U917 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n842, B1 => 
                           REGISTERS_26_13_port, B2 => n829, ZN => n315_port);
   U918 : AND4_X1 port map( A1 => n318_port, A2 => n317_port, A3 => n316_port, 
                           A4 => n315_port, ZN => n330_port);
   U919 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n749, B1 => 
                           REGISTERS_7_13_port, B2 => n732, ZN => n322_port);
   U920 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n783, B1 => 
                           REGISTERS_3_13_port, B2 => n766, ZN => n321_port);
   U921 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n817, B1 => 
                           REGISTERS_6_13_port, B2 => n800, ZN => n320_port);
   U922 : NAND4_X1 port map( A1 => n322_port, A2 => n321_port, A3 => n320_port,
                           A4 => n319_port, ZN => n328_port);
   U923 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n749, B1 => 
                           REGISTERS_15_13_port, B2 => n732, ZN => n326_port);
   U924 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n783, B1 => 
                           REGISTERS_11_13_port, B2 => n766, ZN => n325_port);
   U925 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n817, B1 => 
                           REGISTERS_14_13_port, B2 => n800, ZN => n324_port);
   U926 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n842, B1 => 
                           REGISTERS_10_13_port, B2 => n829, ZN => n323_port);
   U927 : NAND4_X1 port map( A1 => n326_port, A2 => n325_port, A3 => n324_port,
                           A4 => n323_port, ZN => n327_port);
   U928 : AOI22_X1 port map( A1 => n328_port, A2 => n852, B1 => n327_port, B2 
                           => n848, ZN => n329_port);
   U929 : OAI221_X1 port map( B1 => n860, B2 => n331_port, C1 => n856, C2 => 
                           n330_port, A => n329_port, ZN => N211);
   U930 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n749, B1 => 
                           REGISTERS_23_14_port, B2 => n732, ZN => n335_port);
   U931 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n783, B1 => 
                           REGISTERS_19_14_port, B2 => n766, ZN => n334_port);
   U932 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n817, B1 => 
                           REGISTERS_22_14_port, B2 => n800, ZN => n333_port);
   U933 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n842, B1 => 
                           REGISTERS_18_14_port, B2 => n829, ZN => n332_port);
   U934 : AND4_X1 port map( A1 => n335_port, A2 => n334_port, A3 => n333_port, 
                           A4 => n332_port, ZN => n352_port);
   U935 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n749, B1 => 
                           REGISTERS_31_14_port, B2 => n732, ZN => n339_port);
   U936 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n783, B1 => 
                           REGISTERS_27_14_port, B2 => n766, ZN => n338_port);
   U937 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n817, B1 => 
                           REGISTERS_30_14_port, B2 => n800, ZN => n337_port);
   U938 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n842, B1 => 
                           REGISTERS_26_14_port, B2 => n829, ZN => n336_port);
   U939 : AND4_X1 port map( A1 => n339_port, A2 => n338_port, A3 => n337_port, 
                           A4 => n336_port, ZN => n351_port);
   U940 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n749, B1 => 
                           REGISTERS_7_14_port, B2 => n732, ZN => n343_port);
   U941 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n783, B1 => 
                           REGISTERS_3_14_port, B2 => n766, ZN => n342_port);
   U942 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n817, B1 => 
                           REGISTERS_6_14_port, B2 => n800, ZN => n341_port);
   U943 : NAND4_X1 port map( A1 => n343_port, A2 => n342_port, A3 => n341_port,
                           A4 => n340_port, ZN => n349_port);
   U944 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n749, B1 => 
                           REGISTERS_15_14_port, B2 => n732, ZN => n347_port);
   U945 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n783, B1 => 
                           REGISTERS_11_14_port, B2 => n766, ZN => n346_port);
   U946 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n817, B1 => 
                           REGISTERS_14_14_port, B2 => n800, ZN => n345_port);
   U947 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n842, B1 => 
                           REGISTERS_10_14_port, B2 => n829, ZN => n344_port);
   U948 : NAND4_X1 port map( A1 => n347_port, A2 => n346_port, A3 => n345_port,
                           A4 => n344_port, ZN => n348_port);
   U949 : AOI22_X1 port map( A1 => n349_port, A2 => n852, B1 => n348_port, B2 
                           => n848, ZN => n350_port);
   U950 : OAI221_X1 port map( B1 => n860, B2 => n352_port, C1 => n856, C2 => 
                           n351_port, A => n350_port, ZN => N210);
   U951 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n748, B1 => 
                           REGISTERS_23_15_port, B2 => n731, ZN => n356);
   U952 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n782, B1 => 
                           REGISTERS_19_15_port, B2 => n765, ZN => n355);
   U953 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n816, B1 => 
                           REGISTERS_22_15_port, B2 => n799, ZN => n354);
   U954 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n842, B1 => 
                           REGISTERS_18_15_port, B2 => n829, ZN => n353_port);
   U955 : AND4_X1 port map( A1 => n356, A2 => n355, A3 => n354, A4 => n353_port
                           , ZN => n373);
   U956 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n748, B1 => 
                           REGISTERS_31_15_port, B2 => n731, ZN => n360);
   U957 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n782, B1 => 
                           REGISTERS_27_15_port, B2 => n765, ZN => n359);
   U958 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n816, B1 => 
                           REGISTERS_30_15_port, B2 => n799, ZN => n358);
   U959 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n842, B1 => 
                           REGISTERS_26_15_port, B2 => n829, ZN => n357);
   U960 : AND4_X1 port map( A1 => n360, A2 => n359, A3 => n358, A4 => n357, ZN 
                           => n372);
   U961 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n748, B1 => 
                           REGISTERS_7_15_port, B2 => n731, ZN => n364);
   U962 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n782, B1 => 
                           REGISTERS_3_15_port, B2 => n765, ZN => n363);
   U963 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n816, B1 => 
                           REGISTERS_6_15_port, B2 => n799, ZN => n362);
   U964 : NAND4_X1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, ZN
                           => n370);
   U965 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n748, B1 => 
                           REGISTERS_15_15_port, B2 => n731, ZN => n368);
   U966 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n782, B1 => 
                           REGISTERS_11_15_port, B2 => n765, ZN => n367);
   U967 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n816, B1 => 
                           REGISTERS_14_15_port, B2 => n799, ZN => n366);
   U968 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n842, B1 => 
                           REGISTERS_10_15_port, B2 => n828, ZN => n365);
   U969 : NAND4_X1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, ZN
                           => n369);
   U970 : AOI22_X1 port map( A1 => n370, A2 => n852, B1 => n369, B2 => n848, ZN
                           => n371);
   U971 : OAI221_X1 port map( B1 => n860, B2 => n373, C1 => n856, C2 => n372, A
                           => n371, ZN => N209);
   U972 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n748, B1 => 
                           REGISTERS_23_16_port, B2 => n731, ZN => n377);
   U973 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n782, B1 => 
                           REGISTERS_19_16_port, B2 => n765, ZN => n376);
   U974 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n816, B1 => 
                           REGISTERS_22_16_port, B2 => n799, ZN => n375);
   U975 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n841, B1 => 
                           REGISTERS_18_16_port, B2 => n828, ZN => n374);
   U976 : AND4_X1 port map( A1 => n377, A2 => n376, A3 => n375, A4 => n374, ZN 
                           => n394);
   U977 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n748, B1 => 
                           REGISTERS_31_16_port, B2 => n731, ZN => n381);
   U978 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n782, B1 => 
                           REGISTERS_27_16_port, B2 => n765, ZN => n380);
   U979 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n816, B1 => 
                           REGISTERS_30_16_port, B2 => n799, ZN => n379);
   U980 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n841, B1 => 
                           REGISTERS_26_16_port, B2 => n828, ZN => n378);
   U981 : AND4_X1 port map( A1 => n381, A2 => n380, A3 => n379, A4 => n378, ZN 
                           => n393);
   U982 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n748, B1 => 
                           REGISTERS_7_16_port, B2 => n731, ZN => n385);
   U983 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n782, B1 => 
                           REGISTERS_3_16_port, B2 => n765, ZN => n384);
   U984 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n816, B1 => 
                           REGISTERS_6_16_port, B2 => n799, ZN => n383);
   U985 : NAND4_X1 port map( A1 => n385, A2 => n384, A3 => n383, A4 => n382, ZN
                           => n391);
   U986 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n748, B1 => 
                           REGISTERS_15_16_port, B2 => n731, ZN => n389);
   U987 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n782, B1 => 
                           REGISTERS_11_16_port, B2 => n765, ZN => n388);
   U988 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n816, B1 => 
                           REGISTERS_14_16_port, B2 => n799, ZN => n387);
   U989 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n841, B1 => 
                           REGISTERS_10_16_port, B2 => n828, ZN => n386);
   U990 : NAND4_X1 port map( A1 => n389, A2 => n388, A3 => n387, A4 => n386, ZN
                           => n390);
   U991 : AOI22_X1 port map( A1 => n391, A2 => n852, B1 => n390, B2 => n848, ZN
                           => n392);
   U992 : OAI221_X1 port map( B1 => n860, B2 => n394, C1 => n856, C2 => n393, A
                           => n392, ZN => N208);
   U993 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n748, B1 => 
                           REGISTERS_23_17_port, B2 => n731, ZN => n398);
   U994 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n782, B1 => 
                           REGISTERS_19_17_port, B2 => n765, ZN => n397);
   U995 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n816, B1 => 
                           REGISTERS_22_17_port, B2 => n799, ZN => n396);
   U996 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n841, B1 => 
                           REGISTERS_18_17_port, B2 => n828, ZN => n395);
   U997 : AND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN 
                           => n415);
   U998 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n748, B1 => 
                           REGISTERS_31_17_port, B2 => n731, ZN => n402);
   U999 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n782, B1 => 
                           REGISTERS_27_17_port, B2 => n765, ZN => n401);
   U1000 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n816, B1 => 
                           REGISTERS_30_17_port, B2 => n799, ZN => n400);
   U1001 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n841, B1 => 
                           REGISTERS_26_17_port, B2 => n828, ZN => n399);
   U1002 : AND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => n414);
   U1003 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n748, B1 => 
                           REGISTERS_7_17_port, B2 => n731, ZN => n406);
   U1004 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n782, B1 => 
                           REGISTERS_3_17_port, B2 => n765, ZN => n405);
   U1005 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n816, B1 => 
                           REGISTERS_6_17_port, B2 => n799, ZN => n404);
   U1006 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, 
                           ZN => n412);
   U1007 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n748, B1 => 
                           REGISTERS_15_17_port, B2 => n731, ZN => n410);
   U1008 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n782, B1 => 
                           REGISTERS_11_17_port, B2 => n765, ZN => n409);
   U1009 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n816, B1 => 
                           REGISTERS_14_17_port, B2 => n799, ZN => n408);
   U1010 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n841, B1 => 
                           REGISTERS_10_17_port, B2 => n828, ZN => n407);
   U1011 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, 
                           ZN => n411);
   U1012 : AOI22_X1 port map( A1 => n412, A2 => n852, B1 => n411, B2 => n848, 
                           ZN => n413);
   U1013 : OAI221_X1 port map( B1 => n860, B2 => n415, C1 => n856, C2 => n414, 
                           A => n413, ZN => N207);
   U1014 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n747, B1 => 
                           REGISTERS_23_18_port, B2 => n730, ZN => n419);
   U1015 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n781, B1 => 
                           REGISTERS_19_18_port, B2 => n764, ZN => n418);
   U1016 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n815, B1 => 
                           REGISTERS_22_18_port, B2 => n798, ZN => n417);
   U1017 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n841, B1 => 
                           REGISTERS_18_18_port, B2 => n828, ZN => n416);
   U1018 : AND4_X1 port map( A1 => n419, A2 => n418, A3 => n417, A4 => n416, ZN
                           => n436);
   U1019 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n747, B1 => 
                           REGISTERS_31_18_port, B2 => n730, ZN => n423);
   U1020 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n781, B1 => 
                           REGISTERS_27_18_port, B2 => n764, ZN => n422);
   U1021 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n815, B1 => 
                           REGISTERS_30_18_port, B2 => n798, ZN => n421);
   U1022 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n841, B1 => 
                           REGISTERS_26_18_port, B2 => n828, ZN => n420);
   U1023 : AND4_X1 port map( A1 => n423, A2 => n422, A3 => n421, A4 => n420, ZN
                           => n435);
   U1024 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n747, B1 => 
                           REGISTERS_7_18_port, B2 => n730, ZN => n427);
   U1025 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n781, B1 => 
                           REGISTERS_3_18_port, B2 => n764, ZN => n426);
   U1026 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n815, B1 => 
                           REGISTERS_6_18_port, B2 => n798, ZN => n425);
   U1027 : NAND4_X1 port map( A1 => n427, A2 => n426, A3 => n425, A4 => n424, 
                           ZN => n433);
   U1028 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n747, B1 => 
                           REGISTERS_15_18_port, B2 => n730, ZN => n431);
   U1029 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n781, B1 => 
                           REGISTERS_11_18_port, B2 => n764, ZN => n430);
   U1030 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n815, B1 => 
                           REGISTERS_14_18_port, B2 => n798, ZN => n429);
   U1031 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n841, B1 => 
                           REGISTERS_10_18_port, B2 => n828, ZN => n428);
   U1032 : NAND4_X1 port map( A1 => n431, A2 => n430, A3 => n429, A4 => n428, 
                           ZN => n432);
   U1033 : AOI22_X1 port map( A1 => n433, A2 => n852, B1 => n432, B2 => n848, 
                           ZN => n434);
   U1034 : OAI221_X1 port map( B1 => n860, B2 => n436, C1 => n856, C2 => n435, 
                           A => n434, ZN => N206);
   U1035 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n747, B1 => 
                           REGISTERS_23_19_port, B2 => n730, ZN => n440);
   U1036 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n781, B1 => 
                           REGISTERS_19_19_port, B2 => n764, ZN => n439);
   U1037 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n815, B1 => 
                           REGISTERS_22_19_port, B2 => n798, ZN => n438);
   U1038 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n841, B1 => 
                           REGISTERS_18_19_port, B2 => n828, ZN => n437);
   U1039 : AND4_X1 port map( A1 => n440, A2 => n439, A3 => n438, A4 => n437, ZN
                           => n457);
   U1040 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n747, B1 => 
                           REGISTERS_31_19_port, B2 => n730, ZN => n444);
   U1041 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n781, B1 => 
                           REGISTERS_27_19_port, B2 => n764, ZN => n443);
   U1042 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n815, B1 => 
                           REGISTERS_30_19_port, B2 => n798, ZN => n442);
   U1043 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n841, B1 => 
                           REGISTERS_26_19_port, B2 => n828, ZN => n441);
   U1044 : AND4_X1 port map( A1 => n444, A2 => n443, A3 => n442, A4 => n441, ZN
                           => n456);
   U1045 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n747, B1 => 
                           REGISTERS_7_19_port, B2 => n730, ZN => n448);
   U1046 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n781, B1 => 
                           REGISTERS_3_19_port, B2 => n764, ZN => n447);
   U1047 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n815, B1 => 
                           REGISTERS_6_19_port, B2 => n798, ZN => n446);
   U1048 : NAND4_X1 port map( A1 => n448, A2 => n447, A3 => n446, A4 => n445, 
                           ZN => n454);
   U1049 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n747, B1 => 
                           REGISTERS_15_19_port, B2 => n730, ZN => n452);
   U1050 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n781, B1 => 
                           REGISTERS_11_19_port, B2 => n764, ZN => n451);
   U1051 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n815, B1 => 
                           REGISTERS_14_19_port, B2 => n798, ZN => n450);
   U1052 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n841, B1 => 
                           REGISTERS_10_19_port, B2 => n828, ZN => n449);
   U1053 : NAND4_X1 port map( A1 => n452, A2 => n451, A3 => n450, A4 => n449, 
                           ZN => n453);
   U1054 : AOI22_X1 port map( A1 => n454, A2 => n852, B1 => n453, B2 => n848, 
                           ZN => n455);
   U1055 : OAI221_X1 port map( B1 => n860, B2 => n457, C1 => n856, C2 => n456, 
                           A => n455, ZN => N205);
   U1056 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n747, B1 => 
                           REGISTERS_23_20_port, B2 => n730, ZN => n461);
   U1057 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n781, B1 => 
                           REGISTERS_19_20_port, B2 => n764, ZN => n460);
   U1058 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n815, B1 => 
                           REGISTERS_22_20_port, B2 => n798, ZN => n459);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n840, B1 => 
                           REGISTERS_18_20_port, B2 => n828, ZN => n458);
   U1060 : AND4_X1 port map( A1 => n461, A2 => n460, A3 => n459, A4 => n458, ZN
                           => n478);
   U1061 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n747, B1 => 
                           REGISTERS_31_20_port, B2 => n730, ZN => n465);
   U1062 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n781, B1 => 
                           REGISTERS_27_20_port, B2 => n764, ZN => n464);
   U1063 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n815, B1 => 
                           REGISTERS_30_20_port, B2 => n798, ZN => n463);
   U1064 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n840, B1 => 
                           REGISTERS_26_20_port, B2 => n828, ZN => n462);
   U1065 : AND4_X1 port map( A1 => n465, A2 => n464, A3 => n463, A4 => n462, ZN
                           => n477);
   U1066 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n747, B1 => 
                           REGISTERS_7_20_port, B2 => n730, ZN => n469);
   U1067 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n781, B1 => 
                           REGISTERS_3_20_port, B2 => n764, ZN => n468);
   U1068 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n815, B1 => 
                           REGISTERS_6_20_port, B2 => n798, ZN => n467);
   U1069 : NAND4_X1 port map( A1 => n469, A2 => n468, A3 => n467, A4 => n466, 
                           ZN => n475);
   U1070 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n747, B1 => 
                           REGISTERS_15_20_port, B2 => n730, ZN => n473);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n781, B1 => 
                           REGISTERS_11_20_port, B2 => n764, ZN => n472);
   U1072 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n815, B1 => 
                           REGISTERS_14_20_port, B2 => n798, ZN => n471);
   U1073 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n840, B1 => 
                           REGISTERS_10_20_port, B2 => n828, ZN => n470);
   U1074 : NAND4_X1 port map( A1 => n473, A2 => n472, A3 => n471, A4 => n470, 
                           ZN => n474);
   U1075 : AOI22_X1 port map( A1 => n475, A2 => n852, B1 => n474, B2 => n848, 
                           ZN => n476);
   U1076 : OAI221_X1 port map( B1 => n860, B2 => n478, C1 => n857, C2 => n477, 
                           A => n476, ZN => N204);
   U1077 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n746, B1 => 
                           REGISTERS_23_21_port, B2 => n729, ZN => n482);
   U1078 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n780, B1 => 
                           REGISTERS_19_21_port, B2 => n763, ZN => n481);
   U1079 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n814, B1 => 
                           REGISTERS_22_21_port, B2 => n797, ZN => n480);
   U1080 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n840, B1 => 
                           REGISTERS_18_21_port, B2 => n828, ZN => n479);
   U1081 : AND4_X1 port map( A1 => n482, A2 => n481, A3 => n480, A4 => n479, ZN
                           => n499);
   U1082 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n746, B1 => 
                           REGISTERS_31_21_port, B2 => n729, ZN => n486);
   U1083 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n780, B1 => 
                           REGISTERS_27_21_port, B2 => n763, ZN => n485);
   U1084 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n814, B1 => 
                           REGISTERS_30_21_port, B2 => n797, ZN => n484);
   U1085 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n840, B1 => 
                           REGISTERS_26_21_port, B2 => n828, ZN => n483);
   U1086 : AND4_X1 port map( A1 => n486, A2 => n485, A3 => n484, A4 => n483, ZN
                           => n498);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n746, B1 => 
                           REGISTERS_7_21_port, B2 => n729, ZN => n490);
   U1088 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n780, B1 => 
                           REGISTERS_3_21_port, B2 => n763, ZN => n489);
   U1089 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n814, B1 => 
                           REGISTERS_6_21_port, B2 => n797, ZN => n488);
   U1090 : NAND4_X1 port map( A1 => n490, A2 => n489, A3 => n488, A4 => n487, 
                           ZN => n496);
   U1091 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n746, B1 => 
                           REGISTERS_15_21_port, B2 => n729, ZN => n494);
   U1092 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n780, B1 => 
                           REGISTERS_11_21_port, B2 => n763, ZN => n493);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n814, B1 => 
                           REGISTERS_14_21_port, B2 => n797, ZN => n492);
   U1094 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n840, B1 => 
                           REGISTERS_10_21_port, B2 => n828, ZN => n491);
   U1095 : NAND4_X1 port map( A1 => n494, A2 => n493, A3 => n492, A4 => n491, 
                           ZN => n495);
   U1096 : AOI22_X1 port map( A1 => n496, A2 => n852, B1 => n495, B2 => n848, 
                           ZN => n497);
   U1097 : OAI221_X1 port map( B1 => n860, B2 => n499, C1 => n857, C2 => n498, 
                           A => n497, ZN => N203);
   U1098 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n746, B1 => 
                           REGISTERS_23_22_port, B2 => n729, ZN => n503);
   U1099 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n780, B1 => 
                           REGISTERS_19_22_port, B2 => n763, ZN => n502);
   U1100 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n814, B1 => 
                           REGISTERS_22_22_port, B2 => n797, ZN => n501);
   U1101 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n840, B1 => 
                           REGISTERS_18_22_port, B2 => n828, ZN => n500);
   U1102 : AND4_X1 port map( A1 => n503, A2 => n502, A3 => n501, A4 => n500, ZN
                           => n520);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n746, B1 => 
                           REGISTERS_31_22_port, B2 => n729, ZN => n507);
   U1104 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n780, B1 => 
                           REGISTERS_27_22_port, B2 => n763, ZN => n506);
   U1105 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n814, B1 => 
                           REGISTERS_30_22_port, B2 => n797, ZN => n505);
   U1106 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n840, B1 => 
                           REGISTERS_26_22_port, B2 => n827, ZN => n504);
   U1107 : AND4_X1 port map( A1 => n507, A2 => n506, A3 => n505, A4 => n504, ZN
                           => n519);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n746, B1 => 
                           REGISTERS_7_22_port, B2 => n729, ZN => n511);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n780, B1 => 
                           REGISTERS_3_22_port, B2 => n763, ZN => n510);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n814, B1 => 
                           REGISTERS_6_22_port, B2 => n797, ZN => n509);
   U1111 : NAND4_X1 port map( A1 => n511, A2 => n510, A3 => n509, A4 => n508, 
                           ZN => n517);
   U1112 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n746, B1 => 
                           REGISTERS_15_22_port, B2 => n729, ZN => n515);
   U1113 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n780, B1 => 
                           REGISTERS_11_22_port, B2 => n763, ZN => n514);
   U1114 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n814, B1 => 
                           REGISTERS_14_22_port, B2 => n797, ZN => n513);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n840, B1 => 
                           REGISTERS_10_22_port, B2 => n827, ZN => n512);
   U1116 : NAND4_X1 port map( A1 => n515, A2 => n514, A3 => n513, A4 => n512, 
                           ZN => n516);
   U1117 : AOI22_X1 port map( A1 => n517, A2 => n852, B1 => n516, B2 => n848, 
                           ZN => n518);
   U1118 : OAI221_X1 port map( B1 => n860, B2 => n520, C1 => n857, C2 => n519, 
                           A => n518, ZN => N202);
   U1119 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n746, B1 => 
                           REGISTERS_23_23_port, B2 => n729, ZN => n524);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n780, B1 => 
                           REGISTERS_19_23_port, B2 => n763, ZN => n523);
   U1121 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n814, B1 => 
                           REGISTERS_22_23_port, B2 => n797, ZN => n522);
   U1122 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n840, B1 => 
                           REGISTERS_18_23_port, B2 => n827, ZN => n521);
   U1123 : AND4_X1 port map( A1 => n524, A2 => n523, A3 => n522, A4 => n521, ZN
                           => n541);
   U1124 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n746, B1 => 
                           REGISTERS_31_23_port, B2 => n729, ZN => n528);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n780, B1 => 
                           REGISTERS_27_23_port, B2 => n763, ZN => n527);
   U1126 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n814, B1 => 
                           REGISTERS_30_23_port, B2 => n797, ZN => n526);
   U1127 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n840, B1 => 
                           REGISTERS_26_23_port, B2 => n827, ZN => n525);
   U1128 : AND4_X1 port map( A1 => n528, A2 => n527, A3 => n526, A4 => n525, ZN
                           => n540);
   U1129 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n746, B1 => 
                           REGISTERS_7_23_port, B2 => n729, ZN => n532);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n780, B1 => 
                           REGISTERS_3_23_port, B2 => n763, ZN => n531);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n814, B1 => 
                           REGISTERS_6_23_port, B2 => n797, ZN => n530);
   U1132 : NAND4_X1 port map( A1 => n532, A2 => n531, A3 => n530, A4 => n529, 
                           ZN => n538);
   U1133 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n746, B1 => 
                           REGISTERS_15_23_port, B2 => n729, ZN => n536);
   U1134 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n780, B1 => 
                           REGISTERS_11_23_port, B2 => n763, ZN => n535);
   U1135 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n814, B1 => 
                           REGISTERS_14_23_port, B2 => n797, ZN => n534);
   U1136 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n840, B1 => 
                           REGISTERS_10_23_port, B2 => n827, ZN => n533);
   U1137 : NAND4_X1 port map( A1 => n536, A2 => n535, A3 => n534, A4 => n533, 
                           ZN => n537);
   U1138 : AOI22_X1 port map( A1 => n538, A2 => n852, B1 => n537, B2 => n848, 
                           ZN => n539);
   U1139 : OAI221_X1 port map( B1 => n860, B2 => n541, C1 => n857, C2 => n540, 
                           A => n539, ZN => N201);
   U1140 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n745, B1 => 
                           REGISTERS_23_24_port, B2 => n728, ZN => n545);
   U1141 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n779, B1 => 
                           REGISTERS_19_24_port, B2 => n762, ZN => n544);
   U1142 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n813, B1 => 
                           REGISTERS_22_24_port, B2 => n796, ZN => n543);
   U1143 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n839, B1 => 
                           REGISTERS_18_24_port, B2 => n827, ZN => n542);
   U1144 : AND4_X1 port map( A1 => n545, A2 => n544, A3 => n543, A4 => n542, ZN
                           => n562);
   U1145 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n745, B1 => 
                           REGISTERS_31_24_port, B2 => n728, ZN => n549);
   U1146 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n779, B1 => 
                           REGISTERS_27_24_port, B2 => n762, ZN => n548);
   U1147 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n813, B1 => 
                           REGISTERS_30_24_port, B2 => n796, ZN => n547);
   U1148 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n839, B1 => 
                           REGISTERS_26_24_port, B2 => n827, ZN => n546);
   U1149 : AND4_X1 port map( A1 => n549, A2 => n548, A3 => n547, A4 => n546, ZN
                           => n561);
   U1150 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n745, B1 => 
                           REGISTERS_7_24_port, B2 => n728, ZN => n553);
   U1151 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n779, B1 => 
                           REGISTERS_3_24_port, B2 => n762, ZN => n552);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n813, B1 => 
                           REGISTERS_6_24_port, B2 => n796, ZN => n551);
   U1153 : NAND4_X1 port map( A1 => n553, A2 => n552, A3 => n551, A4 => n550, 
                           ZN => n559);
   U1154 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n745, B1 => 
                           REGISTERS_15_24_port, B2 => n728, ZN => n557);
   U1155 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n779, B1 => 
                           REGISTERS_11_24_port, B2 => n762, ZN => n556);
   U1156 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n813, B1 => 
                           REGISTERS_14_24_port, B2 => n796, ZN => n555);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n839, B1 => 
                           REGISTERS_10_24_port, B2 => n827, ZN => n554);
   U1158 : NAND4_X1 port map( A1 => n557, A2 => n556, A3 => n555, A4 => n554, 
                           ZN => n558);
   U1159 : AOI22_X1 port map( A1 => n559, A2 => n851, B1 => n558, B2 => n847, 
                           ZN => n560);
   U1160 : OAI221_X1 port map( B1 => n859, B2 => n562, C1 => n857, C2 => n561, 
                           A => n560, ZN => N200);
   U1161 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n745, B1 => 
                           REGISTERS_23_25_port, B2 => n728, ZN => n566);
   U1162 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n779, B1 => 
                           REGISTERS_19_25_port, B2 => n762, ZN => n565);
   U1163 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n813, B1 => 
                           REGISTERS_22_25_port, B2 => n796, ZN => n564);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n839, B1 => 
                           REGISTERS_18_25_port, B2 => n827, ZN => n563);
   U1165 : AND4_X1 port map( A1 => n566, A2 => n565, A3 => n564, A4 => n563, ZN
                           => n583);
   U1166 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n745, B1 => 
                           REGISTERS_31_25_port, B2 => n728, ZN => n570);
   U1167 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n779, B1 => 
                           REGISTERS_27_25_port, B2 => n762, ZN => n569);
   U1168 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n813, B1 => 
                           REGISTERS_30_25_port, B2 => n796, ZN => n568);
   U1169 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n839, B1 => 
                           REGISTERS_26_25_port, B2 => n827, ZN => n567);
   U1170 : AND4_X1 port map( A1 => n570, A2 => n569, A3 => n568, A4 => n567, ZN
                           => n582);
   U1171 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n745, B1 => 
                           REGISTERS_7_25_port, B2 => n728, ZN => n574);
   U1172 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n779, B1 => 
                           REGISTERS_3_25_port, B2 => n762, ZN => n573);
   U1173 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n813, B1 => 
                           REGISTERS_6_25_port, B2 => n796, ZN => n572);
   U1174 : NAND4_X1 port map( A1 => n574, A2 => n573, A3 => n572, A4 => n571, 
                           ZN => n580);
   U1175 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n745, B1 => 
                           REGISTERS_15_25_port, B2 => n728, ZN => n578);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n779, B1 => 
                           REGISTERS_11_25_port, B2 => n762, ZN => n577);
   U1177 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n813, B1 => 
                           REGISTERS_14_25_port, B2 => n796, ZN => n576);
   U1178 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n839, B1 => 
                           REGISTERS_10_25_port, B2 => n827, ZN => n575);
   U1179 : NAND4_X1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, 
                           ZN => n579);
   U1180 : AOI22_X1 port map( A1 => n580, A2 => n851, B1 => n579, B2 => n847, 
                           ZN => n581);
   U1181 : OAI221_X1 port map( B1 => n859, B2 => n583, C1 => n857, C2 => n582, 
                           A => n581, ZN => N199);
   U1182 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n745, B1 => 
                           REGISTERS_23_26_port, B2 => n728, ZN => n587);
   U1183 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n779, B1 => 
                           REGISTERS_19_26_port, B2 => n762, ZN => n586);
   U1184 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n813, B1 => 
                           REGISTERS_22_26_port, B2 => n796, ZN => n585);
   U1185 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n839, B1 => 
                           REGISTERS_18_26_port, B2 => n827, ZN => n584);
   U1186 : AND4_X1 port map( A1 => n587, A2 => n586, A3 => n585, A4 => n584, ZN
                           => n604);
   U1187 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n745, B1 => 
                           REGISTERS_31_26_port, B2 => n728, ZN => n591);
   U1188 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n779, B1 => 
                           REGISTERS_27_26_port, B2 => n762, ZN => n590);
   U1189 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n813, B1 => 
                           REGISTERS_30_26_port, B2 => n796, ZN => n589);
   U1190 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n839, B1 => 
                           REGISTERS_26_26_port, B2 => n827, ZN => n588);
   U1191 : AND4_X1 port map( A1 => n591, A2 => n590, A3 => n589, A4 => n588, ZN
                           => n603);
   U1192 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n745, B1 => 
                           REGISTERS_7_26_port, B2 => n728, ZN => n595);
   U1193 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n779, B1 => 
                           REGISTERS_3_26_port, B2 => n762, ZN => n594);
   U1194 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n813, B1 => 
                           REGISTERS_6_26_port, B2 => n796, ZN => n593);
   U1195 : NAND4_X1 port map( A1 => n595, A2 => n594, A3 => n593, A4 => n592, 
                           ZN => n601);
   U1196 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n745, B1 => 
                           REGISTERS_15_26_port, B2 => n728, ZN => n599);
   U1197 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n779, B1 => 
                           REGISTERS_11_26_port, B2 => n762, ZN => n598);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n813, B1 => 
                           REGISTERS_14_26_port, B2 => n796, ZN => n597);
   U1199 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n839, B1 => 
                           REGISTERS_10_26_port, B2 => n827, ZN => n596);
   U1200 : NAND4_X1 port map( A1 => n599, A2 => n598, A3 => n597, A4 => n596, 
                           ZN => n600);
   U1201 : AOI22_X1 port map( A1 => n601, A2 => n851, B1 => n600, B2 => n847, 
                           ZN => n602);
   U1202 : OAI221_X1 port map( B1 => n859, B2 => n604, C1 => n857, C2 => n603, 
                           A => n602, ZN => N198);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n744, B1 => 
                           REGISTERS_23_27_port, B2 => n727, ZN => n608);
   U1204 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n778, B1 => 
                           REGISTERS_19_27_port, B2 => n761, ZN => n607);
   U1205 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n812, B1 => 
                           REGISTERS_22_27_port, B2 => n795, ZN => n606);
   U1206 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n839, B1 => 
                           REGISTERS_18_27_port, B2 => n827, ZN => n605);
   U1207 : AND4_X1 port map( A1 => n608, A2 => n607, A3 => n606, A4 => n605, ZN
                           => n625);
   U1208 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n744, B1 => 
                           REGISTERS_31_27_port, B2 => n727, ZN => n612);
   U1209 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n778, B1 => 
                           REGISTERS_27_27_port, B2 => n761, ZN => n611);
   U1210 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n812, B1 => 
                           REGISTERS_30_27_port, B2 => n795, ZN => n610);
   U1211 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n839, B1 => 
                           REGISTERS_26_27_port, B2 => n827, ZN => n609);
   U1212 : AND4_X1 port map( A1 => n612, A2 => n611, A3 => n610, A4 => n609, ZN
                           => n624);
   U1213 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n744, B1 => 
                           REGISTERS_7_27_port, B2 => n727, ZN => n616);
   U1214 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n778, B1 => 
                           REGISTERS_3_27_port, B2 => n761, ZN => n615);
   U1215 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n812, B1 => 
                           REGISTERS_6_27_port, B2 => n795, ZN => n614);
   U1216 : NAND4_X1 port map( A1 => n616, A2 => n615, A3 => n614, A4 => n613, 
                           ZN => n622);
   U1217 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n744, B1 => 
                           REGISTERS_15_27_port, B2 => n727, ZN => n620);
   U1218 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n778, B1 => 
                           REGISTERS_11_27_port, B2 => n761, ZN => n619);
   U1219 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n812, B1 => 
                           REGISTERS_14_27_port, B2 => n795, ZN => n618);
   U1220 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n839, B1 => 
                           REGISTERS_10_27_port, B2 => n827, ZN => n617);
   U1221 : NAND4_X1 port map( A1 => n620, A2 => n619, A3 => n618, A4 => n617, 
                           ZN => n621);
   U1222 : AOI22_X1 port map( A1 => n622, A2 => n851, B1 => n621, B2 => n847, 
                           ZN => n623);
   U1223 : OAI221_X1 port map( B1 => n859, B2 => n625, C1 => n857, C2 => n624, 
                           A => n623, ZN => N197);
   U1224 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n744, B1 => 
                           REGISTERS_23_28_port, B2 => n727, ZN => n629);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n778, B1 => 
                           REGISTERS_19_28_port, B2 => n761, ZN => n628);
   U1226 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n812, B1 => 
                           REGISTERS_22_28_port, B2 => n795, ZN => n627);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n838, B1 => 
                           REGISTERS_18_28_port, B2 => n827, ZN => n626);
   U1228 : AND4_X1 port map( A1 => n629, A2 => n628, A3 => n627, A4 => n626, ZN
                           => n646);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n744, B1 => 
                           REGISTERS_31_28_port, B2 => n727, ZN => n633);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n778, B1 => 
                           REGISTERS_27_28_port, B2 => n761, ZN => n632);
   U1231 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n812, B1 => 
                           REGISTERS_30_28_port, B2 => n795, ZN => n631);
   U1232 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n838, B1 => 
                           REGISTERS_26_28_port, B2 => n827, ZN => n630);
   U1233 : AND4_X1 port map( A1 => n633, A2 => n632, A3 => n631, A4 => n630, ZN
                           => n645);
   U1234 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n744, B1 => 
                           REGISTERS_7_28_port, B2 => n727, ZN => n637);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n778, B1 => 
                           REGISTERS_3_28_port, B2 => n761, ZN => n636);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n812, B1 => 
                           REGISTERS_6_28_port, B2 => n795, ZN => n635);
   U1237 : NAND4_X1 port map( A1 => n637, A2 => n636, A3 => n635, A4 => n634, 
                           ZN => n643);
   U1238 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n744, B1 => 
                           REGISTERS_15_28_port, B2 => n727, ZN => n641);
   U1239 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n778, B1 => 
                           REGISTERS_11_28_port, B2 => n761, ZN => n640);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n812, B1 => 
                           REGISTERS_14_28_port, B2 => n795, ZN => n639);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n838, B1 => 
                           REGISTERS_10_28_port, B2 => n827, ZN => n638);
   U1242 : NAND4_X1 port map( A1 => n641, A2 => n640, A3 => n639, A4 => n638, 
                           ZN => n642);
   U1243 : AOI22_X1 port map( A1 => n643, A2 => n851, B1 => n642, B2 => n847, 
                           ZN => n644);
   U1244 : OAI221_X1 port map( B1 => n859, B2 => n646, C1 => n857, C2 => n645, 
                           A => n644, ZN => N196);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n744, B1 => 
                           REGISTERS_23_29_port, B2 => n727, ZN => n650);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n778, B1 => 
                           REGISTERS_19_29_port, B2 => n761, ZN => n649);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n812, B1 => 
                           REGISTERS_22_29_port, B2 => n795, ZN => n648);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n838, B1 => 
                           REGISTERS_18_29_port, B2 => n826, ZN => n647);
   U1249 : AND4_X1 port map( A1 => n650, A2 => n649, A3 => n648, A4 => n647, ZN
                           => n667);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n744, B1 => 
                           REGISTERS_31_29_port, B2 => n727, ZN => n654);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n778, B1 => 
                           REGISTERS_27_29_port, B2 => n761, ZN => n653);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n812, B1 => 
                           REGISTERS_30_29_port, B2 => n795, ZN => n652);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n838, B1 => 
                           REGISTERS_26_29_port, B2 => n826, ZN => n651);
   U1254 : AND4_X1 port map( A1 => n654, A2 => n653, A3 => n652, A4 => n651, ZN
                           => n666);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n744, B1 => 
                           REGISTERS_7_29_port, B2 => n727, ZN => n658);
   U1256 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n778, B1 => 
                           REGISTERS_3_29_port, B2 => n761, ZN => n657);
   U1257 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n812, B1 => 
                           REGISTERS_6_29_port, B2 => n795, ZN => n656);
   U1258 : NAND4_X1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, 
                           ZN => n664);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n744, B1 => 
                           REGISTERS_15_29_port, B2 => n727, ZN => n662);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n778, B1 => 
                           REGISTERS_11_29_port, B2 => n761, ZN => n661);
   U1261 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n812, B1 => 
                           REGISTERS_14_29_port, B2 => n795, ZN => n660);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n838, B1 => 
                           REGISTERS_10_29_port, B2 => n826, ZN => n659);
   U1263 : NAND4_X1 port map( A1 => n662, A2 => n661, A3 => n660, A4 => n659, 
                           ZN => n663);
   U1264 : AOI22_X1 port map( A1 => n664, A2 => n851, B1 => n663, B2 => n847, 
                           ZN => n665);
   U1265 : OAI221_X1 port map( B1 => n859, B2 => n667, C1 => n857, C2 => n666, 
                           A => n665, ZN => N195);
   U1266 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n743, B1 => 
                           REGISTERS_23_30_port, B2 => n726, ZN => n671);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n777, B1 => 
                           REGISTERS_19_30_port, B2 => n760, ZN => n670);
   U1268 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n811, B1 => 
                           REGISTERS_22_30_port, B2 => n794, ZN => n669);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n838, B1 => 
                           REGISTERS_18_30_port, B2 => n826, ZN => n668);
   U1270 : AND4_X1 port map( A1 => n671, A2 => n670, A3 => n669, A4 => n668, ZN
                           => n688);
   U1271 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n743, B1 => 
                           REGISTERS_31_30_port, B2 => n726, ZN => n675);
   U1272 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n777, B1 => 
                           REGISTERS_27_30_port, B2 => n760, ZN => n674);
   U1273 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n811, B1 => 
                           REGISTERS_30_30_port, B2 => n794, ZN => n673);
   U1274 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n838, B1 => 
                           REGISTERS_26_30_port, B2 => n826, ZN => n672);
   U1275 : AND4_X1 port map( A1 => n675, A2 => n674, A3 => n673, A4 => n672, ZN
                           => n687);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n743, B1 => 
                           REGISTERS_7_30_port, B2 => n726, ZN => n679);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n777, B1 => 
                           REGISTERS_3_30_port, B2 => n760, ZN => n678);
   U1278 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n811, B1 => 
                           REGISTERS_6_30_port, B2 => n794, ZN => n677);
   U1279 : NAND4_X1 port map( A1 => n679, A2 => n678, A3 => n677, A4 => n676, 
                           ZN => n685);
   U1280 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n743, B1 => 
                           REGISTERS_15_30_port, B2 => n726, ZN => n683);
   U1281 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n777, B1 => 
                           REGISTERS_11_30_port, B2 => n760, ZN => n682);
   U1282 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n811, B1 => 
                           REGISTERS_14_30_port, B2 => n794, ZN => n681);
   U1283 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n838, B1 => 
                           REGISTERS_10_30_port, B2 => n826, ZN => n680);
   U1284 : NAND4_X1 port map( A1 => n683, A2 => n682, A3 => n681, A4 => n680, 
                           ZN => n684);
   U1285 : AOI22_X1 port map( A1 => n685, A2 => n851, B1 => n684, B2 => n847, 
                           ZN => n686);
   U1286 : OAI221_X1 port map( B1 => n859, B2 => n688, C1 => n857, C2 => n687, 
                           A => n686, ZN => N194);
   U1287 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n743, B1 => 
                           REGISTERS_23_31_port, B2 => n726, ZN => n692);
   U1288 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n777, B1 => 
                           REGISTERS_19_31_port, B2 => n760, ZN => n691);
   U1289 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n811, B1 => 
                           REGISTERS_22_31_port, B2 => n794, ZN => n690);
   U1290 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n838, B1 => 
                           REGISTERS_18_31_port, B2 => n826, ZN => n689);
   U1291 : AND4_X1 port map( A1 => n692, A2 => n691, A3 => n690, A4 => n689, ZN
                           => n715);
   U1292 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n743, B1 => 
                           REGISTERS_31_31_port, B2 => n726, ZN => n696);
   U1293 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n777, B1 => 
                           REGISTERS_27_31_port, B2 => n760, ZN => n695);
   U1294 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n811, B1 => 
                           REGISTERS_30_31_port, B2 => n794, ZN => n694);
   U1295 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n838, B1 => 
                           REGISTERS_26_31_port, B2 => n826, ZN => n693);
   U1296 : AND4_X1 port map( A1 => n696, A2 => n695, A3 => n694, A4 => n693, ZN
                           => n713);
   U1297 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n743, B1 => 
                           REGISTERS_7_31_port, B2 => n726, ZN => n700);
   U1298 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n777, B1 => 
                           REGISTERS_3_31_port, B2 => n760, ZN => n699);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n811, B1 => 
                           REGISTERS_6_31_port, B2 => n794, ZN => n698);
   U1300 : NAND4_X1 port map( A1 => n700, A2 => n699, A3 => n698, A4 => n697, 
                           ZN => n709);
   U1301 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n743, B1 => 
                           REGISTERS_15_31_port, B2 => n726, ZN => n706);
   U1302 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n777, B1 => 
                           REGISTERS_11_31_port, B2 => n760, ZN => n705);
   U1303 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n811, B1 => 
                           REGISTERS_14_31_port, B2 => n794, ZN => n704);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n838, B1 => 
                           REGISTERS_10_31_port, B2 => n826, ZN => n703);
   U1305 : NAND4_X1 port map( A1 => n706, A2 => n705, A3 => n704, A4 => n703, 
                           ZN => n707);
   U1306 : AOI22_X1 port map( A1 => n851, A2 => n709, B1 => n847, B2 => n707, 
                           ZN => n711);
   U1307 : OAI221_X1 port map( B1 => n715, B2 => n859, C1 => n713, C2 => n857, 
                           A => n711, ZN => N193);
   U1308 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n1547, ZN => n1542);
   U1309 : NOR2_X1 port map( A1 => n1546, A2 => ADD_RD2(1), ZN => n862);
   U1310 : NOR2_X1 port map( A1 => n1546, A2 => n1545, ZN => n863);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n1581, B1 => 
                           REGISTERS_23_0_port, B2 => n1564, ZN => n869);
   U1312 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n864);
   U1313 : NOR2_X1 port map( A1 => n1545, A2 => ADD_RD2(2), ZN => n865);
   U1314 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n1615, B1 => 
                           REGISTERS_19_0_port, B2 => n1598, ZN => n868);
   U1315 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n1649, B1 => 
                           REGISTERS_22_0_port, B2 => n1632, ZN => n867);
   U1316 : AND2_X1 port map( A1 => n864, A2 => n1544, ZN => n1530);
   U1317 : AND2_X1 port map( A1 => n865, A2 => n1544, ZN => n1529);
   U1318 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n1673, B1 => 
                           REGISTERS_18_0_port, B2 => n1659, ZN => n866);
   U1319 : AND4_X1 port map( A1 => n869, A2 => n868, A3 => n867, A4 => n866, ZN
                           => n886);
   U1320 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1540);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n1581, B1 => 
                           REGISTERS_31_0_port, B2 => n1564, ZN => n873);
   U1322 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n1615, B1 => 
                           REGISTERS_27_0_port, B2 => n1598, ZN => n872);
   U1323 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n1649, B1 => 
                           REGISTERS_30_0_port, B2 => n1632, ZN => n871);
   U1324 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n1673, B1 => 
                           REGISTERS_26_0_port, B2 => n1659, ZN => n870);
   U1325 : AND4_X1 port map( A1 => n873, A2 => n872, A3 => n871, A4 => n870, ZN
                           => n885);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n1581, B1 => 
                           REGISTERS_7_0_port, B2 => n1564, ZN => n877);
   U1327 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n1615, B1 => 
                           REGISTERS_3_0_port, B2 => n1598, ZN => n876);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n1649, B1 => 
                           REGISTERS_6_0_port, B2 => n1632, ZN => n875);
   U1329 : NAND4_X1 port map( A1 => n877, A2 => n876, A3 => n875, A4 => n874, 
                           ZN => n883);
   U1330 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1538);
   U1331 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n1581, B1 => 
                           REGISTERS_15_0_port, B2 => n1564, ZN => n881);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n1615, B1 => 
                           REGISTERS_11_0_port, B2 => n1598, ZN => n880);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n1649, B1 => 
                           REGISTERS_14_0_port, B2 => n1632, ZN => n879);
   U1334 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n1673, B1 => 
                           REGISTERS_10_0_port, B2 => n1659, ZN => n878);
   U1335 : NAND4_X1 port map( A1 => n881, A2 => n880, A3 => n879, A4 => n878, 
                           ZN => n882);
   U1336 : NOR2_X1 port map( A1 => n1547, A2 => ADD_RD2(4), ZN => n1536);
   U1337 : AOI22_X1 port map( A1 => n883, A2 => n1681, B1 => n882, B2 => n1677,
                           ZN => n884);
   U1338 : OAI221_X1 port map( B1 => n1689, B2 => n886, C1 => n1683, C2 => n885
                           , A => n884, ZN => N290);
   U1339 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n1581, B1 => 
                           REGISTERS_23_1_port, B2 => n1564, ZN => n890);
   U1340 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n1615, B1 => 
                           REGISTERS_19_1_port, B2 => n1598, ZN => n889);
   U1341 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n1649, B1 => 
                           REGISTERS_22_1_port, B2 => n1632, ZN => n888);
   U1342 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n1673, B1 => 
                           REGISTERS_18_1_port, B2 => n1659, ZN => n887);
   U1343 : AND4_X1 port map( A1 => n890, A2 => n889, A3 => n888, A4 => n887, ZN
                           => n907);
   U1344 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n1581, B1 => 
                           REGISTERS_31_1_port, B2 => n1564, ZN => n894);
   U1345 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n1615, B1 => 
                           REGISTERS_27_1_port, B2 => n1598, ZN => n893);
   U1346 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n1649, B1 => 
                           REGISTERS_30_1_port, B2 => n1632, ZN => n892);
   U1347 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n1673, B1 => 
                           REGISTERS_26_1_port, B2 => n1659, ZN => n891);
   U1348 : AND4_X1 port map( A1 => n894, A2 => n893, A3 => n892, A4 => n891, ZN
                           => n906);
   U1349 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n1581, B1 => 
                           REGISTERS_7_1_port, B2 => n1564, ZN => n898);
   U1350 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n1615, B1 => 
                           REGISTERS_3_1_port, B2 => n1598, ZN => n897);
   U1351 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n1649, B1 => 
                           REGISTERS_6_1_port, B2 => n1632, ZN => n896);
   U1352 : NAND4_X1 port map( A1 => n898, A2 => n897, A3 => n896, A4 => n895, 
                           ZN => n904);
   U1353 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n1581, B1 => 
                           REGISTERS_15_1_port, B2 => n1564, ZN => n902);
   U1354 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n1615, B1 => 
                           REGISTERS_11_1_port, B2 => n1598, ZN => n901);
   U1355 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n1649, B1 => 
                           REGISTERS_14_1_port, B2 => n1632, ZN => n900);
   U1356 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n1673, B1 => 
                           REGISTERS_10_1_port, B2 => n1659, ZN => n899);
   U1357 : NAND4_X1 port map( A1 => n902, A2 => n901, A3 => n900, A4 => n899, 
                           ZN => n903);
   U1358 : AOI22_X1 port map( A1 => n904, A2 => n1681, B1 => n903, B2 => n1677,
                           ZN => n905);
   U1359 : OAI221_X1 port map( B1 => n1689, B2 => n907, C1 => n1683, C2 => n906
                           , A => n905, ZN => N289);
   U1360 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n1581, B1 => 
                           REGISTERS_23_2_port, B2 => n1564, ZN => n911);
   U1361 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n1615, B1 => 
                           REGISTERS_19_2_port, B2 => n1598, ZN => n910);
   U1362 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n1649, B1 => 
                           REGISTERS_22_2_port, B2 => n1632, ZN => n909);
   U1363 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n1673, B1 => 
                           REGISTERS_18_2_port, B2 => n1659, ZN => n908);
   U1364 : AND4_X1 port map( A1 => n911, A2 => n910, A3 => n909, A4 => n908, ZN
                           => n928);
   U1365 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n1581, B1 => 
                           REGISTERS_31_2_port, B2 => n1564, ZN => n915);
   U1366 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n1615, B1 => 
                           REGISTERS_27_2_port, B2 => n1598, ZN => n914);
   U1367 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n1649, B1 => 
                           REGISTERS_30_2_port, B2 => n1632, ZN => n913);
   U1368 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n1673, B1 => 
                           REGISTERS_26_2_port, B2 => n1658, ZN => n912);
   U1369 : AND4_X1 port map( A1 => n915, A2 => n914, A3 => n913, A4 => n912, ZN
                           => n927);
   U1370 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n1581, B1 => 
                           REGISTERS_7_2_port, B2 => n1564, ZN => n919);
   U1371 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n1615, B1 => 
                           REGISTERS_3_2_port, B2 => n1598, ZN => n918);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n1649, B1 => 
                           REGISTERS_6_2_port, B2 => n1632, ZN => n917);
   U1373 : NAND4_X1 port map( A1 => n919, A2 => n918, A3 => n917, A4 => n916, 
                           ZN => n925);
   U1374 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n1581, B1 => 
                           REGISTERS_15_2_port, B2 => n1564, ZN => n923);
   U1375 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n1615, B1 => 
                           REGISTERS_11_2_port, B2 => n1598, ZN => n922);
   U1376 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n1649, B1 => 
                           REGISTERS_14_2_port, B2 => n1632, ZN => n921);
   U1377 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n1673, B1 => 
                           REGISTERS_10_2_port, B2 => n1658, ZN => n920);
   U1378 : NAND4_X1 port map( A1 => n923, A2 => n922, A3 => n921, A4 => n920, 
                           ZN => n924);
   U1379 : AOI22_X1 port map( A1 => n925, A2 => n1681, B1 => n924, B2 => n1677,
                           ZN => n926);
   U1380 : OAI221_X1 port map( B1 => n1689, B2 => n928, C1 => n1683, C2 => n927
                           , A => n926, ZN => N288);
   U1381 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n1580, B1 => 
                           REGISTERS_23_3_port, B2 => n1563, ZN => n932);
   U1382 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n1614, B1 => 
                           REGISTERS_19_3_port, B2 => n1597, ZN => n931);
   U1383 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n1648, B1 => 
                           REGISTERS_22_3_port, B2 => n1631, ZN => n930);
   U1384 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n1673, B1 => 
                           REGISTERS_18_3_port, B2 => n1658, ZN => n929);
   U1385 : AND4_X1 port map( A1 => n932, A2 => n931, A3 => n930, A4 => n929, ZN
                           => n949);
   U1386 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n1580, B1 => 
                           REGISTERS_31_3_port, B2 => n1563, ZN => n936);
   U1387 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n1614, B1 => 
                           REGISTERS_27_3_port, B2 => n1597, ZN => n935);
   U1388 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n1648, B1 => 
                           REGISTERS_30_3_port, B2 => n1631, ZN => n934);
   U1389 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n1673, B1 => 
                           REGISTERS_26_3_port, B2 => n1658, ZN => n933);
   U1390 : AND4_X1 port map( A1 => n936, A2 => n935, A3 => n934, A4 => n933, ZN
                           => n948);
   U1391 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n1580, B1 => 
                           REGISTERS_7_3_port, B2 => n1563, ZN => n940);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n1614, B1 => 
                           REGISTERS_3_3_port, B2 => n1597, ZN => n939);
   U1393 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n1648, B1 => 
                           REGISTERS_6_3_port, B2 => n1631, ZN => n938);
   U1394 : NAND4_X1 port map( A1 => n940, A2 => n939, A3 => n938, A4 => n937, 
                           ZN => n946);
   U1395 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n1580, B1 => 
                           REGISTERS_15_3_port, B2 => n1563, ZN => n944);
   U1396 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n1614, B1 => 
                           REGISTERS_11_3_port, B2 => n1597, ZN => n943);
   U1397 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n1648, B1 => 
                           REGISTERS_14_3_port, B2 => n1631, ZN => n942);
   U1398 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n1673, B1 => 
                           REGISTERS_10_3_port, B2 => n1658, ZN => n941);
   U1399 : NAND4_X1 port map( A1 => n944, A2 => n943, A3 => n942, A4 => n941, 
                           ZN => n945);
   U1400 : AOI22_X1 port map( A1 => n946, A2 => n1681, B1 => n945, B2 => n1677,
                           ZN => n947);
   U1401 : OAI221_X1 port map( B1 => n1689, B2 => n949, C1 => n1683, C2 => n948
                           , A => n947, ZN => N287);
   U1402 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n1580, B1 => 
                           REGISTERS_23_4_port, B2 => n1563, ZN => n953);
   U1403 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n1614, B1 => 
                           REGISTERS_19_4_port, B2 => n1597, ZN => n952);
   U1404 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n1648, B1 => 
                           REGISTERS_22_4_port, B2 => n1631, ZN => n951);
   U1405 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n1672, B1 => 
                           REGISTERS_18_4_port, B2 => n1658, ZN => n950);
   U1406 : AND4_X1 port map( A1 => n953, A2 => n952, A3 => n951, A4 => n950, ZN
                           => n970);
   U1407 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n1580, B1 => 
                           REGISTERS_31_4_port, B2 => n1563, ZN => n957);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n1614, B1 => 
                           REGISTERS_27_4_port, B2 => n1597, ZN => n956);
   U1409 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n1648, B1 => 
                           REGISTERS_30_4_port, B2 => n1631, ZN => n955);
   U1410 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n1672, B1 => 
                           REGISTERS_26_4_port, B2 => n1658, ZN => n954);
   U1411 : AND4_X1 port map( A1 => n957, A2 => n956, A3 => n955, A4 => n954, ZN
                           => n969);
   U1412 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n1580, B1 => 
                           REGISTERS_7_4_port, B2 => n1563, ZN => n961);
   U1413 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n1614, B1 => 
                           REGISTERS_3_4_port, B2 => n1597, ZN => n960);
   U1414 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n1648, B1 => 
                           REGISTERS_6_4_port, B2 => n1631, ZN => n959);
   U1415 : NAND4_X1 port map( A1 => n961, A2 => n960, A3 => n959, A4 => n958, 
                           ZN => n967);
   U1416 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n1580, B1 => 
                           REGISTERS_15_4_port, B2 => n1563, ZN => n965);
   U1417 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n1614, B1 => 
                           REGISTERS_11_4_port, B2 => n1597, ZN => n964);
   U1418 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n1648, B1 => 
                           REGISTERS_14_4_port, B2 => n1631, ZN => n963);
   U1419 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n1672, B1 => 
                           REGISTERS_10_4_port, B2 => n1658, ZN => n962);
   U1420 : NAND4_X1 port map( A1 => n965, A2 => n964, A3 => n963, A4 => n962, 
                           ZN => n966);
   U1421 : AOI22_X1 port map( A1 => n967, A2 => n1681, B1 => n966, B2 => n1677,
                           ZN => n968);
   U1422 : OAI221_X1 port map( B1 => n1689, B2 => n970, C1 => n1683, C2 => n969
                           , A => n968, ZN => N286);
   U1423 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n1580, B1 => 
                           REGISTERS_23_5_port, B2 => n1563, ZN => n974);
   U1424 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n1614, B1 => 
                           REGISTERS_19_5_port, B2 => n1597, ZN => n973);
   U1425 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n1648, B1 => 
                           REGISTERS_22_5_port, B2 => n1631, ZN => n972);
   U1426 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n1672, B1 => 
                           REGISTERS_18_5_port, B2 => n1658, ZN => n971);
   U1427 : AND4_X1 port map( A1 => n974, A2 => n973, A3 => n972, A4 => n971, ZN
                           => n991);
   U1428 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n1580, B1 => 
                           REGISTERS_31_5_port, B2 => n1563, ZN => n978);
   U1429 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n1614, B1 => 
                           REGISTERS_27_5_port, B2 => n1597, ZN => n977);
   U1430 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n1648, B1 => 
                           REGISTERS_30_5_port, B2 => n1631, ZN => n976);
   U1431 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n1672, B1 => 
                           REGISTERS_26_5_port, B2 => n1658, ZN => n975);
   U1432 : AND4_X1 port map( A1 => n978, A2 => n977, A3 => n976, A4 => n975, ZN
                           => n990);
   U1433 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n1580, B1 => 
                           REGISTERS_7_5_port, B2 => n1563, ZN => n982);
   U1434 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n1614, B1 => 
                           REGISTERS_3_5_port, B2 => n1597, ZN => n981);
   U1435 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n1648, B1 => 
                           REGISTERS_6_5_port, B2 => n1631, ZN => n980);
   U1436 : NAND4_X1 port map( A1 => n982, A2 => n981, A3 => n980, A4 => n979, 
                           ZN => n988);
   U1437 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n1580, B1 => 
                           REGISTERS_15_5_port, B2 => n1563, ZN => n986);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n1614, B1 => 
                           REGISTERS_11_5_port, B2 => n1597, ZN => n985);
   U1439 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n1648, B1 => 
                           REGISTERS_14_5_port, B2 => n1631, ZN => n984);
   U1440 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n1672, B1 => 
                           REGISTERS_10_5_port, B2 => n1658, ZN => n983);
   U1441 : NAND4_X1 port map( A1 => n986, A2 => n985, A3 => n984, A4 => n983, 
                           ZN => n987);
   U1442 : AOI22_X1 port map( A1 => n988, A2 => n1681, B1 => n987, B2 => n1677,
                           ZN => n989);
   U1443 : OAI221_X1 port map( B1 => n1689, B2 => n991, C1 => n1683, C2 => n990
                           , A => n989, ZN => N285);
   U1444 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n1579, B1 => 
                           REGISTERS_23_6_port, B2 => n1562, ZN => n995);
   U1445 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n1613, B1 => 
                           REGISTERS_19_6_port, B2 => n1596, ZN => n994);
   U1446 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n1647, B1 => 
                           REGISTERS_22_6_port, B2 => n1630, ZN => n993);
   U1447 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n1672, B1 => 
                           REGISTERS_18_6_port, B2 => n1658, ZN => n992);
   U1448 : AND4_X1 port map( A1 => n995, A2 => n994, A3 => n993, A4 => n992, ZN
                           => n1012);
   U1449 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n1579, B1 => 
                           REGISTERS_31_6_port, B2 => n1562, ZN => n999);
   U1450 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n1613, B1 => 
                           REGISTERS_27_6_port, B2 => n1596, ZN => n998);
   U1451 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n1647, B1 => 
                           REGISTERS_30_6_port, B2 => n1630, ZN => n997);
   U1452 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n1672, B1 => 
                           REGISTERS_26_6_port, B2 => n1658, ZN => n996);
   U1453 : AND4_X1 port map( A1 => n999, A2 => n998, A3 => n997, A4 => n996, ZN
                           => n1011);
   U1454 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n1579, B1 => 
                           REGISTERS_7_6_port, B2 => n1562, ZN => n1003);
   U1455 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n1613, B1 => 
                           REGISTERS_3_6_port, B2 => n1596, ZN => n1002);
   U1456 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n1647, B1 => 
                           REGISTERS_6_6_port, B2 => n1630, ZN => n1001);
   U1457 : NAND4_X1 port map( A1 => n1003, A2 => n1002, A3 => n1001, A4 => 
                           n1000, ZN => n1009);
   U1458 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n1579, B1 => 
                           REGISTERS_15_6_port, B2 => n1562, ZN => n1007);
   U1459 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n1613, B1 => 
                           REGISTERS_11_6_port, B2 => n1596, ZN => n1006);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n1647, B1 => 
                           REGISTERS_14_6_port, B2 => n1630, ZN => n1005);
   U1461 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n1672, B1 => 
                           REGISTERS_10_6_port, B2 => n1658, ZN => n1004);
   U1462 : NAND4_X1 port map( A1 => n1007, A2 => n1006, A3 => n1005, A4 => 
                           n1004, ZN => n1008);
   U1463 : AOI22_X1 port map( A1 => n1009, A2 => n1681, B1 => n1008, B2 => 
                           n1677, ZN => n1010);
   U1464 : OAI221_X1 port map( B1 => n1689, B2 => n1012, C1 => n1683, C2 => 
                           n1011, A => n1010, ZN => N284);
   U1465 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n1579, B1 => 
                           REGISTERS_23_7_port, B2 => n1562, ZN => n1016);
   U1466 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n1613, B1 => 
                           REGISTERS_19_7_port, B2 => n1596, ZN => n1015);
   U1467 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n1647, B1 => 
                           REGISTERS_22_7_port, B2 => n1630, ZN => n1014);
   U1468 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n1672, B1 => 
                           REGISTERS_18_7_port, B2 => n1658, ZN => n1013);
   U1469 : AND4_X1 port map( A1 => n1016, A2 => n1015, A3 => n1014, A4 => n1013
                           , ZN => n1033);
   U1470 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n1579, B1 => 
                           REGISTERS_31_7_port, B2 => n1562, ZN => n1020);
   U1471 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n1613, B1 => 
                           REGISTERS_27_7_port, B2 => n1596, ZN => n1019);
   U1472 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n1647, B1 => 
                           REGISTERS_30_7_port, B2 => n1630, ZN => n1018);
   U1473 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n1672, B1 => 
                           REGISTERS_26_7_port, B2 => n1658, ZN => n1017);
   U1474 : AND4_X1 port map( A1 => n1020, A2 => n1019, A3 => n1018, A4 => n1017
                           , ZN => n1032);
   U1475 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n1579, B1 => 
                           REGISTERS_7_7_port, B2 => n1562, ZN => n1024);
   U1476 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n1613, B1 => 
                           REGISTERS_3_7_port, B2 => n1596, ZN => n1023);
   U1477 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n1647, B1 => 
                           REGISTERS_6_7_port, B2 => n1630, ZN => n1022);
   U1478 : NAND4_X1 port map( A1 => n1024, A2 => n1023, A3 => n1022, A4 => 
                           n1021, ZN => n1030);
   U1479 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n1579, B1 => 
                           REGISTERS_15_7_port, B2 => n1562, ZN => n1028);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n1613, B1 => 
                           REGISTERS_11_7_port, B2 => n1596, ZN => n1027);
   U1481 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n1647, B1 => 
                           REGISTERS_14_7_port, B2 => n1630, ZN => n1026);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n1672, B1 => 
                           REGISTERS_10_7_port, B2 => n1658, ZN => n1025);
   U1483 : NAND4_X1 port map( A1 => n1028, A2 => n1027, A3 => n1026, A4 => 
                           n1025, ZN => n1029);
   U1484 : AOI22_X1 port map( A1 => n1030, A2 => n1681, B1 => n1029, B2 => 
                           n1677, ZN => n1031);
   U1485 : OAI221_X1 port map( B1 => n1689, B2 => n1033, C1 => n1683, C2 => 
                           n1032, A => n1031, ZN => N283);
   U1486 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n1579, B1 => 
                           REGISTERS_23_8_port, B2 => n1562, ZN => n1037);
   U1487 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n1613, B1 => 
                           REGISTERS_19_8_port, B2 => n1596, ZN => n1036);
   U1488 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n1647, B1 => 
                           REGISTERS_22_8_port, B2 => n1630, ZN => n1035);
   U1489 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n1671, B1 => 
                           REGISTERS_18_8_port, B2 => n1658, ZN => n1034);
   U1490 : AND4_X1 port map( A1 => n1037, A2 => n1036, A3 => n1035, A4 => n1034
                           , ZN => n1054);
   U1491 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n1579, B1 => 
                           REGISTERS_31_8_port, B2 => n1562, ZN => n1041);
   U1492 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n1613, B1 => 
                           REGISTERS_27_8_port, B2 => n1596, ZN => n1040);
   U1493 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n1647, B1 => 
                           REGISTERS_30_8_port, B2 => n1630, ZN => n1039);
   U1494 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n1671, B1 => 
                           REGISTERS_26_8_port, B2 => n1658, ZN => n1038);
   U1495 : AND4_X1 port map( A1 => n1041, A2 => n1040, A3 => n1039, A4 => n1038
                           , ZN => n1053);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n1579, B1 => 
                           REGISTERS_7_8_port, B2 => n1562, ZN => n1045);
   U1497 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n1613, B1 => 
                           REGISTERS_3_8_port, B2 => n1596, ZN => n1044);
   U1498 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n1647, B1 => 
                           REGISTERS_6_8_port, B2 => n1630, ZN => n1043);
   U1499 : NAND4_X1 port map( A1 => n1045, A2 => n1044, A3 => n1043, A4 => 
                           n1042, ZN => n1051);
   U1500 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n1579, B1 => 
                           REGISTERS_15_8_port, B2 => n1562, ZN => n1049);
   U1501 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n1613, B1 => 
                           REGISTERS_11_8_port, B2 => n1596, ZN => n1048);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n1647, B1 => 
                           REGISTERS_14_8_port, B2 => n1630, ZN => n1047);
   U1503 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n1671, B1 => 
                           REGISTERS_10_8_port, B2 => n1658, ZN => n1046);
   U1504 : NAND4_X1 port map( A1 => n1049, A2 => n1048, A3 => n1047, A4 => 
                           n1046, ZN => n1050);
   U1505 : AOI22_X1 port map( A1 => n1051, A2 => n1681, B1 => n1050, B2 => 
                           n1677, ZN => n1052);
   U1506 : OAI221_X1 port map( B1 => n1689, B2 => n1054, C1 => n1684, C2 => 
                           n1053, A => n1052, ZN => N282);
   U1507 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n1578, B1 => 
                           REGISTERS_23_9_port, B2 => n1561, ZN => n1058);
   U1508 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n1612, B1 => 
                           REGISTERS_19_9_port, B2 => n1595, ZN => n1057);
   U1509 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n1646, B1 => 
                           REGISTERS_22_9_port, B2 => n1629, ZN => n1056);
   U1510 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n1671, B1 => 
                           REGISTERS_18_9_port, B2 => n1657, ZN => n1055);
   U1511 : AND4_X1 port map( A1 => n1058, A2 => n1057, A3 => n1056, A4 => n1055
                           , ZN => n1075);
   U1512 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n1578, B1 => 
                           REGISTERS_31_9_port, B2 => n1561, ZN => n1062);
   U1513 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n1612, B1 => 
                           REGISTERS_27_9_port, B2 => n1595, ZN => n1061);
   U1514 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n1646, B1 => 
                           REGISTERS_30_9_port, B2 => n1629, ZN => n1060);
   U1515 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n1671, B1 => 
                           REGISTERS_26_9_port, B2 => n1657, ZN => n1059);
   U1516 : AND4_X1 port map( A1 => n1062, A2 => n1061, A3 => n1060, A4 => n1059
                           , ZN => n1074);
   U1517 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n1578, B1 => 
                           REGISTERS_7_9_port, B2 => n1561, ZN => n1066);
   U1518 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n1612, B1 => 
                           REGISTERS_3_9_port, B2 => n1595, ZN => n1065);
   U1519 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n1646, B1 => 
                           REGISTERS_6_9_port, B2 => n1629, ZN => n1064);
   U1520 : NAND4_X1 port map( A1 => n1066, A2 => n1065, A3 => n1064, A4 => 
                           n1063, ZN => n1072);
   U1521 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n1578, B1 => 
                           REGISTERS_15_9_port, B2 => n1561, ZN => n1070);
   U1522 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n1612, B1 => 
                           REGISTERS_11_9_port, B2 => n1595, ZN => n1069);
   U1523 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n1646, B1 => 
                           REGISTERS_14_9_port, B2 => n1629, ZN => n1068);
   U1524 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n1671, B1 => 
                           REGISTERS_10_9_port, B2 => n1657, ZN => n1067);
   U1525 : NAND4_X1 port map( A1 => n1070, A2 => n1069, A3 => n1068, A4 => 
                           n1067, ZN => n1071);
   U1526 : AOI22_X1 port map( A1 => n1072, A2 => n1681, B1 => n1071, B2 => 
                           n1677, ZN => n1073);
   U1527 : OAI221_X1 port map( B1 => n1689, B2 => n1075, C1 => n1684, C2 => 
                           n1074, A => n1073, ZN => N281);
   U1528 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n1578, B1 => 
                           REGISTERS_23_10_port, B2 => n1561, ZN => n1079);
   U1529 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n1612, B1 => 
                           REGISTERS_19_10_port, B2 => n1595, ZN => n1078);
   U1530 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n1646, B1 => 
                           REGISTERS_22_10_port, B2 => n1629, ZN => n1077);
   U1531 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n1671, B1 => 
                           REGISTERS_18_10_port, B2 => n1657, ZN => n1076);
   U1532 : AND4_X1 port map( A1 => n1079, A2 => n1078, A3 => n1077, A4 => n1076
                           , ZN => n1096);
   U1533 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n1578, B1 => 
                           REGISTERS_31_10_port, B2 => n1561, ZN => n1083);
   U1534 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n1612, B1 => 
                           REGISTERS_27_10_port, B2 => n1595, ZN => n1082);
   U1535 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n1646, B1 => 
                           REGISTERS_30_10_port, B2 => n1629, ZN => n1081);
   U1536 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n1671, B1 => 
                           REGISTERS_26_10_port, B2 => n1657, ZN => n1080);
   U1537 : AND4_X1 port map( A1 => n1083, A2 => n1082, A3 => n1081, A4 => n1080
                           , ZN => n1095);
   U1538 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n1578, B1 => 
                           REGISTERS_7_10_port, B2 => n1561, ZN => n1087);
   U1539 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n1612, B1 => 
                           REGISTERS_3_10_port, B2 => n1595, ZN => n1086);
   U1540 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n1646, B1 => 
                           REGISTERS_6_10_port, B2 => n1629, ZN => n1085);
   U1541 : NAND4_X1 port map( A1 => n1087, A2 => n1086, A3 => n1085, A4 => 
                           n1084, ZN => n1093);
   U1542 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n1578, B1 => 
                           REGISTERS_15_10_port, B2 => n1561, ZN => n1091);
   U1543 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n1612, B1 => 
                           REGISTERS_11_10_port, B2 => n1595, ZN => n1090);
   U1544 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n1646, B1 => 
                           REGISTERS_14_10_port, B2 => n1629, ZN => n1089);
   U1545 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n1671, B1 => 
                           REGISTERS_10_10_port, B2 => n1657, ZN => n1088);
   U1546 : NAND4_X1 port map( A1 => n1091, A2 => n1090, A3 => n1089, A4 => 
                           n1088, ZN => n1092);
   U1547 : AOI22_X1 port map( A1 => n1093, A2 => n1681, B1 => n1092, B2 => 
                           n1677, ZN => n1094);
   U1548 : OAI221_X1 port map( B1 => n1689, B2 => n1096, C1 => n1684, C2 => 
                           n1095, A => n1094, ZN => N280);
   U1549 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n1578, B1 => 
                           REGISTERS_23_11_port, B2 => n1561, ZN => n1100);
   U1550 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n1612, B1 => 
                           REGISTERS_19_11_port, B2 => n1595, ZN => n1099);
   U1551 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n1646, B1 => 
                           REGISTERS_22_11_port, B2 => n1629, ZN => n1098);
   U1552 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n1671, B1 => 
                           REGISTERS_18_11_port, B2 => n1657, ZN => n1097);
   U1553 : AND4_X1 port map( A1 => n1100, A2 => n1099, A3 => n1098, A4 => n1097
                           , ZN => n1117);
   U1554 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n1578, B1 => 
                           REGISTERS_31_11_port, B2 => n1561, ZN => n1104);
   U1555 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n1612, B1 => 
                           REGISTERS_27_11_port, B2 => n1595, ZN => n1103);
   U1556 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n1646, B1 => 
                           REGISTERS_30_11_port, B2 => n1629, ZN => n1102);
   U1557 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n1671, B1 => 
                           REGISTERS_26_11_port, B2 => n1657, ZN => n1101);
   U1558 : AND4_X1 port map( A1 => n1104, A2 => n1103, A3 => n1102, A4 => n1101
                           , ZN => n1116);
   U1559 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n1578, B1 => 
                           REGISTERS_7_11_port, B2 => n1561, ZN => n1108);
   U1560 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n1612, B1 => 
                           REGISTERS_3_11_port, B2 => n1595, ZN => n1107);
   U1561 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n1646, B1 => 
                           REGISTERS_6_11_port, B2 => n1629, ZN => n1106);
   U1562 : NAND4_X1 port map( A1 => n1108, A2 => n1107, A3 => n1106, A4 => 
                           n1105, ZN => n1114);
   U1563 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n1578, B1 => 
                           REGISTERS_15_11_port, B2 => n1561, ZN => n1112);
   U1564 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n1612, B1 => 
                           REGISTERS_11_11_port, B2 => n1595, ZN => n1111);
   U1565 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n1646, B1 => 
                           REGISTERS_14_11_port, B2 => n1629, ZN => n1110);
   U1566 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n1671, B1 => 
                           REGISTERS_10_11_port, B2 => n1657, ZN => n1109);
   U1567 : NAND4_X1 port map( A1 => n1112, A2 => n1111, A3 => n1110, A4 => 
                           n1109, ZN => n1113);
   U1568 : AOI22_X1 port map( A1 => n1114, A2 => n1681, B1 => n1113, B2 => 
                           n1677, ZN => n1115);
   U1569 : OAI221_X1 port map( B1 => n1689, B2 => n1117, C1 => n1684, C2 => 
                           n1116, A => n1115, ZN => N279);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n1577, B1 => 
                           REGISTERS_23_12_port, B2 => n1560, ZN => n1121);
   U1571 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n1611, B1 => 
                           REGISTERS_19_12_port, B2 => n1594, ZN => n1120);
   U1572 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n1645, B1 => 
                           REGISTERS_22_12_port, B2 => n1628, ZN => n1119);
   U1573 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n1670, B1 => 
                           REGISTERS_18_12_port, B2 => n1657, ZN => n1118);
   U1574 : AND4_X1 port map( A1 => n1121, A2 => n1120, A3 => n1119, A4 => n1118
                           , ZN => n1138);
   U1575 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n1577, B1 => 
                           REGISTERS_31_12_port, B2 => n1560, ZN => n1125);
   U1576 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n1611, B1 => 
                           REGISTERS_27_12_port, B2 => n1594, ZN => n1124);
   U1577 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n1645, B1 => 
                           REGISTERS_30_12_port, B2 => n1628, ZN => n1123);
   U1578 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n1670, B1 => 
                           REGISTERS_26_12_port, B2 => n1657, ZN => n1122);
   U1579 : AND4_X1 port map( A1 => n1125, A2 => n1124, A3 => n1123, A4 => n1122
                           , ZN => n1137);
   U1580 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n1577, B1 => 
                           REGISTERS_7_12_port, B2 => n1560, ZN => n1129);
   U1581 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n1611, B1 => 
                           REGISTERS_3_12_port, B2 => n1594, ZN => n1128);
   U1582 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n1645, B1 => 
                           REGISTERS_6_12_port, B2 => n1628, ZN => n1127);
   U1583 : NAND4_X1 port map( A1 => n1129, A2 => n1128, A3 => n1127, A4 => 
                           n1126, ZN => n1135);
   U1584 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n1577, B1 => 
                           REGISTERS_15_12_port, B2 => n1560, ZN => n1133);
   U1585 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n1611, B1 => 
                           REGISTERS_11_12_port, B2 => n1594, ZN => n1132);
   U1586 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n1645, B1 => 
                           REGISTERS_14_12_port, B2 => n1628, ZN => n1131);
   U1587 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n1670, B1 => 
                           REGISTERS_10_12_port, B2 => n1657, ZN => n1130);
   U1588 : NAND4_X1 port map( A1 => n1133, A2 => n1132, A3 => n1131, A4 => 
                           n1130, ZN => n1134);
   U1589 : AOI22_X1 port map( A1 => n1135, A2 => n1680, B1 => n1134, B2 => 
                           n1676, ZN => n1136);
   U1590 : OAI221_X1 port map( B1 => n1688, B2 => n1138, C1 => n1684, C2 => 
                           n1137, A => n1136, ZN => N278);
   U1591 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n1577, B1 => 
                           REGISTERS_23_13_port, B2 => n1560, ZN => n1142);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n1611, B1 => 
                           REGISTERS_19_13_port, B2 => n1594, ZN => n1141);
   U1593 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n1645, B1 => 
                           REGISTERS_22_13_port, B2 => n1628, ZN => n1140);
   U1594 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n1670, B1 => 
                           REGISTERS_18_13_port, B2 => n1657, ZN => n1139);
   U1595 : AND4_X1 port map( A1 => n1142, A2 => n1141, A3 => n1140, A4 => n1139
                           , ZN => n1159);
   U1596 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n1577, B1 => 
                           REGISTERS_31_13_port, B2 => n1560, ZN => n1146);
   U1597 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n1611, B1 => 
                           REGISTERS_27_13_port, B2 => n1594, ZN => n1145);
   U1598 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n1645, B1 => 
                           REGISTERS_30_13_port, B2 => n1628, ZN => n1144);
   U1599 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n1670, B1 => 
                           REGISTERS_26_13_port, B2 => n1657, ZN => n1143);
   U1600 : AND4_X1 port map( A1 => n1146, A2 => n1145, A3 => n1144, A4 => n1143
                           , ZN => n1158);
   U1601 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n1577, B1 => 
                           REGISTERS_7_13_port, B2 => n1560, ZN => n1150);
   U1602 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n1611, B1 => 
                           REGISTERS_3_13_port, B2 => n1594, ZN => n1149);
   U1603 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n1645, B1 => 
                           REGISTERS_6_13_port, B2 => n1628, ZN => n1148);
   U1604 : NAND4_X1 port map( A1 => n1150, A2 => n1149, A3 => n1148, A4 => 
                           n1147, ZN => n1156);
   U1605 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n1577, B1 => 
                           REGISTERS_15_13_port, B2 => n1560, ZN => n1154);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n1611, B1 => 
                           REGISTERS_11_13_port, B2 => n1594, ZN => n1153);
   U1607 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n1645, B1 => 
                           REGISTERS_14_13_port, B2 => n1628, ZN => n1152);
   U1608 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n1670, B1 => 
                           REGISTERS_10_13_port, B2 => n1657, ZN => n1151);
   U1609 : NAND4_X1 port map( A1 => n1154, A2 => n1153, A3 => n1152, A4 => 
                           n1151, ZN => n1155);
   U1610 : AOI22_X1 port map( A1 => n1156, A2 => n1680, B1 => n1155, B2 => 
                           n1676, ZN => n1157);
   U1611 : OAI221_X1 port map( B1 => n1688, B2 => n1159, C1 => n1684, C2 => 
                           n1158, A => n1157, ZN => N277);
   U1612 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n1577, B1 => 
                           REGISTERS_23_14_port, B2 => n1560, ZN => n1163);
   U1613 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n1611, B1 => 
                           REGISTERS_19_14_port, B2 => n1594, ZN => n1162);
   U1614 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n1645, B1 => 
                           REGISTERS_22_14_port, B2 => n1628, ZN => n1161);
   U1615 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n1670, B1 => 
                           REGISTERS_18_14_port, B2 => n1657, ZN => n1160);
   U1616 : AND4_X1 port map( A1 => n1163, A2 => n1162, A3 => n1161, A4 => n1160
                           , ZN => n1180);
   U1617 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n1577, B1 => 
                           REGISTERS_31_14_port, B2 => n1560, ZN => n1167);
   U1618 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n1611, B1 => 
                           REGISTERS_27_14_port, B2 => n1594, ZN => n1166);
   U1619 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n1645, B1 => 
                           REGISTERS_30_14_port, B2 => n1628, ZN => n1165);
   U1620 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n1670, B1 => 
                           REGISTERS_26_14_port, B2 => n1657, ZN => n1164);
   U1621 : AND4_X1 port map( A1 => n1167, A2 => n1166, A3 => n1165, A4 => n1164
                           , ZN => n1179);
   U1622 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n1577, B1 => 
                           REGISTERS_7_14_port, B2 => n1560, ZN => n1171);
   U1623 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n1611, B1 => 
                           REGISTERS_3_14_port, B2 => n1594, ZN => n1170);
   U1624 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n1645, B1 => 
                           REGISTERS_6_14_port, B2 => n1628, ZN => n1169);
   U1625 : NAND4_X1 port map( A1 => n1171, A2 => n1170, A3 => n1169, A4 => 
                           n1168, ZN => n1177);
   U1626 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n1577, B1 => 
                           REGISTERS_15_14_port, B2 => n1560, ZN => n1175);
   U1627 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n1611, B1 => 
                           REGISTERS_11_14_port, B2 => n1594, ZN => n1174);
   U1628 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n1645, B1 => 
                           REGISTERS_14_14_port, B2 => n1628, ZN => n1173);
   U1629 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n1670, B1 => 
                           REGISTERS_10_14_port, B2 => n1657, ZN => n1172);
   U1630 : NAND4_X1 port map( A1 => n1175, A2 => n1174, A3 => n1173, A4 => 
                           n1172, ZN => n1176);
   U1631 : AOI22_X1 port map( A1 => n1177, A2 => n1680, B1 => n1176, B2 => 
                           n1676, ZN => n1178);
   U1632 : OAI221_X1 port map( B1 => n1688, B2 => n1180, C1 => n1684, C2 => 
                           n1179, A => n1178, ZN => N276);
   U1633 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n1576, B1 => 
                           REGISTERS_23_15_port, B2 => n1559, ZN => n1184);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n1610, B1 => 
                           REGISTERS_19_15_port, B2 => n1593, ZN => n1183);
   U1635 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n1644, B1 => 
                           REGISTERS_22_15_port, B2 => n1627, ZN => n1182);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n1670, B1 => 
                           REGISTERS_18_15_port, B2 => n1657, ZN => n1181);
   U1637 : AND4_X1 port map( A1 => n1184, A2 => n1183, A3 => n1182, A4 => n1181
                           , ZN => n1201);
   U1638 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n1576, B1 => 
                           REGISTERS_31_15_port, B2 => n1559, ZN => n1188);
   U1639 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n1610, B1 => 
                           REGISTERS_27_15_port, B2 => n1593, ZN => n1187);
   U1640 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n1644, B1 => 
                           REGISTERS_30_15_port, B2 => n1627, ZN => n1186);
   U1641 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n1670, B1 => 
                           REGISTERS_26_15_port, B2 => n1657, ZN => n1185);
   U1642 : AND4_X1 port map( A1 => n1188, A2 => n1187, A3 => n1186, A4 => n1185
                           , ZN => n1200);
   U1643 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n1576, B1 => 
                           REGISTERS_7_15_port, B2 => n1559, ZN => n1192);
   U1644 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n1610, B1 => 
                           REGISTERS_3_15_port, B2 => n1593, ZN => n1191);
   U1645 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n1644, B1 => 
                           REGISTERS_6_15_port, B2 => n1627, ZN => n1190);
   U1646 : NAND4_X1 port map( A1 => n1192, A2 => n1191, A3 => n1190, A4 => 
                           n1189, ZN => n1198);
   U1647 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n1576, B1 => 
                           REGISTERS_15_15_port, B2 => n1559, ZN => n1196);
   U1648 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n1610, B1 => 
                           REGISTERS_11_15_port, B2 => n1593, ZN => n1195);
   U1649 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n1644, B1 => 
                           REGISTERS_14_15_port, B2 => n1627, ZN => n1194);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n1670, B1 => 
                           REGISTERS_10_15_port, B2 => n1656, ZN => n1193);
   U1651 : NAND4_X1 port map( A1 => n1196, A2 => n1195, A3 => n1194, A4 => 
                           n1193, ZN => n1197);
   U1652 : AOI22_X1 port map( A1 => n1198, A2 => n1680, B1 => n1197, B2 => 
                           n1676, ZN => n1199);
   U1653 : OAI221_X1 port map( B1 => n1688, B2 => n1201, C1 => n1684, C2 => 
                           n1200, A => n1199, ZN => N275);
   U1654 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n1576, B1 => 
                           REGISTERS_23_16_port, B2 => n1559, ZN => n1205);
   U1655 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n1610, B1 => 
                           REGISTERS_19_16_port, B2 => n1593, ZN => n1204);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n1644, B1 => 
                           REGISTERS_22_16_port, B2 => n1627, ZN => n1203);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n1669, B1 => 
                           REGISTERS_18_16_port, B2 => n1656, ZN => n1202);
   U1658 : AND4_X1 port map( A1 => n1205, A2 => n1204, A3 => n1203, A4 => n1202
                           , ZN => n1222);
   U1659 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n1576, B1 => 
                           REGISTERS_31_16_port, B2 => n1559, ZN => n1209);
   U1660 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n1610, B1 => 
                           REGISTERS_27_16_port, B2 => n1593, ZN => n1208);
   U1661 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n1644, B1 => 
                           REGISTERS_30_16_port, B2 => n1627, ZN => n1207);
   U1662 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n1669, B1 => 
                           REGISTERS_26_16_port, B2 => n1656, ZN => n1206);
   U1663 : AND4_X1 port map( A1 => n1209, A2 => n1208, A3 => n1207, A4 => n1206
                           , ZN => n1221);
   U1664 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n1576, B1 => 
                           REGISTERS_7_16_port, B2 => n1559, ZN => n1213);
   U1665 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n1610, B1 => 
                           REGISTERS_3_16_port, B2 => n1593, ZN => n1212);
   U1666 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n1644, B1 => 
                           REGISTERS_6_16_port, B2 => n1627, ZN => n1211);
   U1667 : NAND4_X1 port map( A1 => n1213, A2 => n1212, A3 => n1211, A4 => 
                           n1210, ZN => n1219);
   U1668 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n1576, B1 => 
                           REGISTERS_15_16_port, B2 => n1559, ZN => n1217);
   U1669 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n1610, B1 => 
                           REGISTERS_11_16_port, B2 => n1593, ZN => n1216);
   U1670 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n1644, B1 => 
                           REGISTERS_14_16_port, B2 => n1627, ZN => n1215);
   U1671 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n1669, B1 => 
                           REGISTERS_10_16_port, B2 => n1656, ZN => n1214);
   U1672 : NAND4_X1 port map( A1 => n1217, A2 => n1216, A3 => n1215, A4 => 
                           n1214, ZN => n1218);
   U1673 : AOI22_X1 port map( A1 => n1219, A2 => n1680, B1 => n1218, B2 => 
                           n1676, ZN => n1220);
   U1674 : OAI221_X1 port map( B1 => n1688, B2 => n1222, C1 => n1684, C2 => 
                           n1221, A => n1220, ZN => N274);
   U1675 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n1576, B1 => 
                           REGISTERS_23_17_port, B2 => n1559, ZN => n1226);
   U1676 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n1610, B1 => 
                           REGISTERS_19_17_port, B2 => n1593, ZN => n1225);
   U1677 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n1644, B1 => 
                           REGISTERS_22_17_port, B2 => n1627, ZN => n1224);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n1669, B1 => 
                           REGISTERS_18_17_port, B2 => n1656, ZN => n1223);
   U1679 : AND4_X1 port map( A1 => n1226, A2 => n1225, A3 => n1224, A4 => n1223
                           , ZN => n1243);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n1576, B1 => 
                           REGISTERS_31_17_port, B2 => n1559, ZN => n1230);
   U1681 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n1610, B1 => 
                           REGISTERS_27_17_port, B2 => n1593, ZN => n1229);
   U1682 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n1644, B1 => 
                           REGISTERS_30_17_port, B2 => n1627, ZN => n1228);
   U1683 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n1669, B1 => 
                           REGISTERS_26_17_port, B2 => n1656, ZN => n1227);
   U1684 : AND4_X1 port map( A1 => n1230, A2 => n1229, A3 => n1228, A4 => n1227
                           , ZN => n1242);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n1576, B1 => 
                           REGISTERS_7_17_port, B2 => n1559, ZN => n1234);
   U1686 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n1610, B1 => 
                           REGISTERS_3_17_port, B2 => n1593, ZN => n1233);
   U1687 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n1644, B1 => 
                           REGISTERS_6_17_port, B2 => n1627, ZN => n1232);
   U1688 : NAND4_X1 port map( A1 => n1234, A2 => n1233, A3 => n1232, A4 => 
                           n1231, ZN => n1240);
   U1689 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n1576, B1 => 
                           REGISTERS_15_17_port, B2 => n1559, ZN => n1238);
   U1690 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n1610, B1 => 
                           REGISTERS_11_17_port, B2 => n1593, ZN => n1237);
   U1691 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n1644, B1 => 
                           REGISTERS_14_17_port, B2 => n1627, ZN => n1236);
   U1692 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n1669, B1 => 
                           REGISTERS_10_17_port, B2 => n1656, ZN => n1235);
   U1693 : NAND4_X1 port map( A1 => n1238, A2 => n1237, A3 => n1236, A4 => 
                           n1235, ZN => n1239);
   U1694 : AOI22_X1 port map( A1 => n1240, A2 => n1680, B1 => n1239, B2 => 
                           n1676, ZN => n1241);
   U1695 : OAI221_X1 port map( B1 => n1688, B2 => n1243, C1 => n1684, C2 => 
                           n1242, A => n1241, ZN => N273);
   U1696 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n1575, B1 => 
                           REGISTERS_23_18_port, B2 => n1558, ZN => n1247);
   U1697 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n1609, B1 => 
                           REGISTERS_19_18_port, B2 => n1592, ZN => n1246);
   U1698 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n1643, B1 => 
                           REGISTERS_22_18_port, B2 => n1626, ZN => n1245);
   U1699 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n1669, B1 => 
                           REGISTERS_18_18_port, B2 => n1656, ZN => n1244);
   U1700 : AND4_X1 port map( A1 => n1247, A2 => n1246, A3 => n1245, A4 => n1244
                           , ZN => n1264);
   U1701 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n1575, B1 => 
                           REGISTERS_31_18_port, B2 => n1558, ZN => n1251);
   U1702 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n1609, B1 => 
                           REGISTERS_27_18_port, B2 => n1592, ZN => n1250);
   U1703 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n1643, B1 => 
                           REGISTERS_30_18_port, B2 => n1626, ZN => n1249);
   U1704 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n1669, B1 => 
                           REGISTERS_26_18_port, B2 => n1656, ZN => n1248);
   U1705 : AND4_X1 port map( A1 => n1251, A2 => n1250, A3 => n1249, A4 => n1248
                           , ZN => n1263);
   U1706 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n1575, B1 => 
                           REGISTERS_7_18_port, B2 => n1558, ZN => n1255);
   U1707 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n1609, B1 => 
                           REGISTERS_3_18_port, B2 => n1592, ZN => n1254);
   U1708 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n1643, B1 => 
                           REGISTERS_6_18_port, B2 => n1626, ZN => n1253);
   U1709 : NAND4_X1 port map( A1 => n1255, A2 => n1254, A3 => n1253, A4 => 
                           n1252, ZN => n1261);
   U1710 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n1575, B1 => 
                           REGISTERS_15_18_port, B2 => n1558, ZN => n1259);
   U1711 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n1609, B1 => 
                           REGISTERS_11_18_port, B2 => n1592, ZN => n1258);
   U1712 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n1643, B1 => 
                           REGISTERS_14_18_port, B2 => n1626, ZN => n1257);
   U1713 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n1669, B1 => 
                           REGISTERS_10_18_port, B2 => n1656, ZN => n1256);
   U1714 : NAND4_X1 port map( A1 => n1259, A2 => n1258, A3 => n1257, A4 => 
                           n1256, ZN => n1260);
   U1715 : AOI22_X1 port map( A1 => n1261, A2 => n1680, B1 => n1260, B2 => 
                           n1676, ZN => n1262);
   U1716 : OAI221_X1 port map( B1 => n1688, B2 => n1264, C1 => n1684, C2 => 
                           n1263, A => n1262, ZN => N272);
   U1717 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n1575, B1 => 
                           REGISTERS_23_19_port, B2 => n1558, ZN => n1268);
   U1718 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n1609, B1 => 
                           REGISTERS_19_19_port, B2 => n1592, ZN => n1267);
   U1719 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n1643, B1 => 
                           REGISTERS_22_19_port, B2 => n1626, ZN => n1266);
   U1720 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n1669, B1 => 
                           REGISTERS_18_19_port, B2 => n1656, ZN => n1265);
   U1721 : AND4_X1 port map( A1 => n1268, A2 => n1267, A3 => n1266, A4 => n1265
                           , ZN => n1285);
   U1722 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n1575, B1 => 
                           REGISTERS_31_19_port, B2 => n1558, ZN => n1272);
   U1723 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n1609, B1 => 
                           REGISTERS_27_19_port, B2 => n1592, ZN => n1271);
   U1724 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n1643, B1 => 
                           REGISTERS_30_19_port, B2 => n1626, ZN => n1270);
   U1725 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n1669, B1 => 
                           REGISTERS_26_19_port, B2 => n1656, ZN => n1269);
   U1726 : AND4_X1 port map( A1 => n1272, A2 => n1271, A3 => n1270, A4 => n1269
                           , ZN => n1284);
   U1727 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n1575, B1 => 
                           REGISTERS_7_19_port, B2 => n1558, ZN => n1276);
   U1728 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n1609, B1 => 
                           REGISTERS_3_19_port, B2 => n1592, ZN => n1275);
   U1729 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n1643, B1 => 
                           REGISTERS_6_19_port, B2 => n1626, ZN => n1274);
   U1730 : NAND4_X1 port map( A1 => n1276, A2 => n1275, A3 => n1274, A4 => 
                           n1273, ZN => n1282);
   U1731 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n1575, B1 => 
                           REGISTERS_15_19_port, B2 => n1558, ZN => n1280);
   U1732 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n1609, B1 => 
                           REGISTERS_11_19_port, B2 => n1592, ZN => n1279);
   U1733 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n1643, B1 => 
                           REGISTERS_14_19_port, B2 => n1626, ZN => n1278);
   U1734 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n1669, B1 => 
                           REGISTERS_10_19_port, B2 => n1656, ZN => n1277);
   U1735 : NAND4_X1 port map( A1 => n1280, A2 => n1279, A3 => n1278, A4 => 
                           n1277, ZN => n1281);
   U1736 : AOI22_X1 port map( A1 => n1282, A2 => n1680, B1 => n1281, B2 => 
                           n1676, ZN => n1283);
   U1737 : OAI221_X1 port map( B1 => n1688, B2 => n1285, C1 => n1684, C2 => 
                           n1284, A => n1283, ZN => N271);
   U1738 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n1575, B1 => 
                           REGISTERS_23_20_port, B2 => n1558, ZN => n1289);
   U1739 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n1609, B1 => 
                           REGISTERS_19_20_port, B2 => n1592, ZN => n1288);
   U1740 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n1643, B1 => 
                           REGISTERS_22_20_port, B2 => n1626, ZN => n1287);
   U1741 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n1668, B1 => 
                           REGISTERS_18_20_port, B2 => n1656, ZN => n1286);
   U1742 : AND4_X1 port map( A1 => n1289, A2 => n1288, A3 => n1287, A4 => n1286
                           , ZN => n1306);
   U1743 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n1575, B1 => 
                           REGISTERS_31_20_port, B2 => n1558, ZN => n1293);
   U1744 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n1609, B1 => 
                           REGISTERS_27_20_port, B2 => n1592, ZN => n1292);
   U1745 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n1643, B1 => 
                           REGISTERS_30_20_port, B2 => n1626, ZN => n1291);
   U1746 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n1668, B1 => 
                           REGISTERS_26_20_port, B2 => n1656, ZN => n1290);
   U1747 : AND4_X1 port map( A1 => n1293, A2 => n1292, A3 => n1291, A4 => n1290
                           , ZN => n1305);
   U1748 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n1575, B1 => 
                           REGISTERS_7_20_port, B2 => n1558, ZN => n1297);
   U1749 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n1609, B1 => 
                           REGISTERS_3_20_port, B2 => n1592, ZN => n1296);
   U1750 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n1643, B1 => 
                           REGISTERS_6_20_port, B2 => n1626, ZN => n1295);
   U1751 : NAND4_X1 port map( A1 => n1297, A2 => n1296, A3 => n1295, A4 => 
                           n1294, ZN => n1303);
   U1752 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n1575, B1 => 
                           REGISTERS_15_20_port, B2 => n1558, ZN => n1301);
   U1753 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n1609, B1 => 
                           REGISTERS_11_20_port, B2 => n1592, ZN => n1300);
   U1754 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n1643, B1 => 
                           REGISTERS_14_20_port, B2 => n1626, ZN => n1299);
   U1755 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n1668, B1 => 
                           REGISTERS_10_20_port, B2 => n1656, ZN => n1298);
   U1756 : NAND4_X1 port map( A1 => n1301, A2 => n1300, A3 => n1299, A4 => 
                           n1298, ZN => n1302);
   U1757 : AOI22_X1 port map( A1 => n1303, A2 => n1680, B1 => n1302, B2 => 
                           n1676, ZN => n1304);
   U1758 : OAI221_X1 port map( B1 => n1688, B2 => n1306, C1 => n1685, C2 => 
                           n1305, A => n1304, ZN => N270);
   U1759 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n1574, B1 => 
                           REGISTERS_23_21_port, B2 => n1557, ZN => n1310);
   U1760 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n1608, B1 => 
                           REGISTERS_19_21_port, B2 => n1591, ZN => n1309);
   U1761 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n1642, B1 => 
                           REGISTERS_22_21_port, B2 => n1625, ZN => n1308);
   U1762 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n1668, B1 => 
                           REGISTERS_18_21_port, B2 => n1656, ZN => n1307);
   U1763 : AND4_X1 port map( A1 => n1310, A2 => n1309, A3 => n1308, A4 => n1307
                           , ZN => n1327);
   U1764 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n1574, B1 => 
                           REGISTERS_31_21_port, B2 => n1557, ZN => n1314);
   U1765 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n1608, B1 => 
                           REGISTERS_27_21_port, B2 => n1591, ZN => n1313);
   U1766 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n1642, B1 => 
                           REGISTERS_30_21_port, B2 => n1625, ZN => n1312);
   U1767 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n1668, B1 => 
                           REGISTERS_26_21_port, B2 => n1656, ZN => n1311);
   U1768 : AND4_X1 port map( A1 => n1314, A2 => n1313, A3 => n1312, A4 => n1311
                           , ZN => n1326);
   U1769 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n1574, B1 => 
                           REGISTERS_7_21_port, B2 => n1557, ZN => n1318);
   U1770 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n1608, B1 => 
                           REGISTERS_3_21_port, B2 => n1591, ZN => n1317);
   U1771 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n1642, B1 => 
                           REGISTERS_6_21_port, B2 => n1625, ZN => n1316);
   U1772 : NAND4_X1 port map( A1 => n1318, A2 => n1317, A3 => n1316, A4 => 
                           n1315, ZN => n1324);
   U1773 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n1574, B1 => 
                           REGISTERS_15_21_port, B2 => n1557, ZN => n1322);
   U1774 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n1608, B1 => 
                           REGISTERS_11_21_port, B2 => n1591, ZN => n1321);
   U1775 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n1642, B1 => 
                           REGISTERS_14_21_port, B2 => n1625, ZN => n1320);
   U1776 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n1668, B1 => 
                           REGISTERS_10_21_port, B2 => n1656, ZN => n1319);
   U1777 : NAND4_X1 port map( A1 => n1322, A2 => n1321, A3 => n1320, A4 => 
                           n1319, ZN => n1323);
   U1778 : AOI22_X1 port map( A1 => n1324, A2 => n1680, B1 => n1323, B2 => 
                           n1676, ZN => n1325);
   U1779 : OAI221_X1 port map( B1 => n1688, B2 => n1327, C1 => n1685, C2 => 
                           n1326, A => n1325, ZN => N269);
   U1780 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n1574, B1 => 
                           REGISTERS_23_22_port, B2 => n1557, ZN => n1331);
   U1781 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n1608, B1 => 
                           REGISTERS_19_22_port, B2 => n1591, ZN => n1330);
   U1782 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n1642, B1 => 
                           REGISTERS_22_22_port, B2 => n1625, ZN => n1329);
   U1783 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n1668, B1 => 
                           REGISTERS_18_22_port, B2 => n1656, ZN => n1328);
   U1784 : AND4_X1 port map( A1 => n1331, A2 => n1330, A3 => n1329, A4 => n1328
                           , ZN => n1348);
   U1785 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n1574, B1 => 
                           REGISTERS_31_22_port, B2 => n1557, ZN => n1335);
   U1786 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n1608, B1 => 
                           REGISTERS_27_22_port, B2 => n1591, ZN => n1334);
   U1787 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n1642, B1 => 
                           REGISTERS_30_22_port, B2 => n1625, ZN => n1333);
   U1788 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n1668, B1 => 
                           REGISTERS_26_22_port, B2 => n1655, ZN => n1332);
   U1789 : AND4_X1 port map( A1 => n1335, A2 => n1334, A3 => n1333, A4 => n1332
                           , ZN => n1347);
   U1790 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n1574, B1 => 
                           REGISTERS_7_22_port, B2 => n1557, ZN => n1339);
   U1791 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n1608, B1 => 
                           REGISTERS_3_22_port, B2 => n1591, ZN => n1338);
   U1792 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n1642, B1 => 
                           REGISTERS_6_22_port, B2 => n1625, ZN => n1337);
   U1793 : NAND4_X1 port map( A1 => n1339, A2 => n1338, A3 => n1337, A4 => 
                           n1336, ZN => n1345);
   U1794 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n1574, B1 => 
                           REGISTERS_15_22_port, B2 => n1557, ZN => n1343);
   U1795 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n1608, B1 => 
                           REGISTERS_11_22_port, B2 => n1591, ZN => n1342);
   U1796 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n1642, B1 => 
                           REGISTERS_14_22_port, B2 => n1625, ZN => n1341);
   U1797 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n1668, B1 => 
                           REGISTERS_10_22_port, B2 => n1655, ZN => n1340);
   U1798 : NAND4_X1 port map( A1 => n1343, A2 => n1342, A3 => n1341, A4 => 
                           n1340, ZN => n1344);
   U1799 : AOI22_X1 port map( A1 => n1345, A2 => n1680, B1 => n1344, B2 => 
                           n1676, ZN => n1346);
   U1800 : OAI221_X1 port map( B1 => n1688, B2 => n1348, C1 => n1685, C2 => 
                           n1347, A => n1346, ZN => N268);
   U1801 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n1574, B1 => 
                           REGISTERS_23_23_port, B2 => n1557, ZN => n1352);
   U1802 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n1608, B1 => 
                           REGISTERS_19_23_port, B2 => n1591, ZN => n1351);
   U1803 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n1642, B1 => 
                           REGISTERS_22_23_port, B2 => n1625, ZN => n1350);
   U1804 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n1668, B1 => 
                           REGISTERS_18_23_port, B2 => n1655, ZN => n1349);
   U1805 : AND4_X1 port map( A1 => n1352, A2 => n1351, A3 => n1350, A4 => n1349
                           , ZN => n1369);
   U1806 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n1574, B1 => 
                           REGISTERS_31_23_port, B2 => n1557, ZN => n1356);
   U1807 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n1608, B1 => 
                           REGISTERS_27_23_port, B2 => n1591, ZN => n1355);
   U1808 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n1642, B1 => 
                           REGISTERS_30_23_port, B2 => n1625, ZN => n1354);
   U1809 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n1668, B1 => 
                           REGISTERS_26_23_port, B2 => n1655, ZN => n1353);
   U1810 : AND4_X1 port map( A1 => n1356, A2 => n1355, A3 => n1354, A4 => n1353
                           , ZN => n1368);
   U1811 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n1574, B1 => 
                           REGISTERS_7_23_port, B2 => n1557, ZN => n1360);
   U1812 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n1608, B1 => 
                           REGISTERS_3_23_port, B2 => n1591, ZN => n1359);
   U1813 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n1642, B1 => 
                           REGISTERS_6_23_port, B2 => n1625, ZN => n1358);
   U1814 : NAND4_X1 port map( A1 => n1360, A2 => n1359, A3 => n1358, A4 => 
                           n1357, ZN => n1366);
   U1815 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n1574, B1 => 
                           REGISTERS_15_23_port, B2 => n1557, ZN => n1364);
   U1816 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n1608, B1 => 
                           REGISTERS_11_23_port, B2 => n1591, ZN => n1363);
   U1817 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n1642, B1 => 
                           REGISTERS_14_23_port, B2 => n1625, ZN => n1362);
   U1818 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n1668, B1 => 
                           REGISTERS_10_23_port, B2 => n1655, ZN => n1361);
   U1819 : NAND4_X1 port map( A1 => n1364, A2 => n1363, A3 => n1362, A4 => 
                           n1361, ZN => n1365);
   U1820 : AOI22_X1 port map( A1 => n1366, A2 => n1680, B1 => n1365, B2 => 
                           n1676, ZN => n1367);
   U1821 : OAI221_X1 port map( B1 => n1688, B2 => n1369, C1 => n1685, C2 => 
                           n1368, A => n1367, ZN => N267);
   U1822 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n1573, B1 => 
                           REGISTERS_23_24_port, B2 => n1556, ZN => n1373);
   U1823 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n1607, B1 => 
                           REGISTERS_19_24_port, B2 => n1590, ZN => n1372);
   U1824 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n1641, B1 => 
                           REGISTERS_22_24_port, B2 => n1624, ZN => n1371);
   U1825 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n1667, B1 => 
                           REGISTERS_18_24_port, B2 => n1655, ZN => n1370);
   U1826 : AND4_X1 port map( A1 => n1373, A2 => n1372, A3 => n1371, A4 => n1370
                           , ZN => n1390);
   U1827 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n1573, B1 => 
                           REGISTERS_31_24_port, B2 => n1556, ZN => n1377);
   U1828 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n1607, B1 => 
                           REGISTERS_27_24_port, B2 => n1590, ZN => n1376);
   U1829 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n1641, B1 => 
                           REGISTERS_30_24_port, B2 => n1624, ZN => n1375);
   U1830 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n1667, B1 => 
                           REGISTERS_26_24_port, B2 => n1655, ZN => n1374);
   U1831 : AND4_X1 port map( A1 => n1377, A2 => n1376, A3 => n1375, A4 => n1374
                           , ZN => n1389);
   U1832 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n1573, B1 => 
                           REGISTERS_7_24_port, B2 => n1556, ZN => n1381);
   U1833 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n1607, B1 => 
                           REGISTERS_3_24_port, B2 => n1590, ZN => n1380);
   U1834 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n1641, B1 => 
                           REGISTERS_6_24_port, B2 => n1624, ZN => n1379);
   U1835 : NAND4_X1 port map( A1 => n1381, A2 => n1380, A3 => n1379, A4 => 
                           n1378, ZN => n1387);
   U1836 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n1573, B1 => 
                           REGISTERS_15_24_port, B2 => n1556, ZN => n1385);
   U1837 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n1607, B1 => 
                           REGISTERS_11_24_port, B2 => n1590, ZN => n1384);
   U1838 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n1641, B1 => 
                           REGISTERS_14_24_port, B2 => n1624, ZN => n1383);
   U1839 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n1667, B1 => 
                           REGISTERS_10_24_port, B2 => n1655, ZN => n1382);
   U1840 : NAND4_X1 port map( A1 => n1385, A2 => n1384, A3 => n1383, A4 => 
                           n1382, ZN => n1386);
   U1841 : AOI22_X1 port map( A1 => n1387, A2 => n1679, B1 => n1386, B2 => 
                           n1675, ZN => n1388);
   U1842 : OAI221_X1 port map( B1 => n1687, B2 => n1390, C1 => n1685, C2 => 
                           n1389, A => n1388, ZN => N266);
   U1843 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n1573, B1 => 
                           REGISTERS_23_25_port, B2 => n1556, ZN => n1394);
   U1844 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n1607, B1 => 
                           REGISTERS_19_25_port, B2 => n1590, ZN => n1393);
   U1845 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n1641, B1 => 
                           REGISTERS_22_25_port, B2 => n1624, ZN => n1392);
   U1846 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n1667, B1 => 
                           REGISTERS_18_25_port, B2 => n1655, ZN => n1391);
   U1847 : AND4_X1 port map( A1 => n1394, A2 => n1393, A3 => n1392, A4 => n1391
                           , ZN => n1411);
   U1848 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n1573, B1 => 
                           REGISTERS_31_25_port, B2 => n1556, ZN => n1398);
   U1849 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n1607, B1 => 
                           REGISTERS_27_25_port, B2 => n1590, ZN => n1397);
   U1850 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n1641, B1 => 
                           REGISTERS_30_25_port, B2 => n1624, ZN => n1396);
   U1851 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n1667, B1 => 
                           REGISTERS_26_25_port, B2 => n1655, ZN => n1395);
   U1852 : AND4_X1 port map( A1 => n1398, A2 => n1397, A3 => n1396, A4 => n1395
                           , ZN => n1410);
   U1853 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n1573, B1 => 
                           REGISTERS_7_25_port, B2 => n1556, ZN => n1402);
   U1854 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n1607, B1 => 
                           REGISTERS_3_25_port, B2 => n1590, ZN => n1401);
   U1855 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n1641, B1 => 
                           REGISTERS_6_25_port, B2 => n1624, ZN => n1400);
   U1856 : NAND4_X1 port map( A1 => n1402, A2 => n1401, A3 => n1400, A4 => 
                           n1399, ZN => n1408);
   U1857 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n1573, B1 => 
                           REGISTERS_15_25_port, B2 => n1556, ZN => n1406);
   U1858 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n1607, B1 => 
                           REGISTERS_11_25_port, B2 => n1590, ZN => n1405);
   U1859 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n1641, B1 => 
                           REGISTERS_14_25_port, B2 => n1624, ZN => n1404);
   U1860 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n1667, B1 => 
                           REGISTERS_10_25_port, B2 => n1655, ZN => n1403);
   U1861 : NAND4_X1 port map( A1 => n1406, A2 => n1405, A3 => n1404, A4 => 
                           n1403, ZN => n1407);
   U1862 : AOI22_X1 port map( A1 => n1408, A2 => n1679, B1 => n1407, B2 => 
                           n1675, ZN => n1409);
   U1863 : OAI221_X1 port map( B1 => n1687, B2 => n1411, C1 => n1685, C2 => 
                           n1410, A => n1409, ZN => N265);
   U1864 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n1573, B1 => 
                           REGISTERS_23_26_port, B2 => n1556, ZN => n1415);
   U1865 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n1607, B1 => 
                           REGISTERS_19_26_port, B2 => n1590, ZN => n1414);
   U1866 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n1641, B1 => 
                           REGISTERS_22_26_port, B2 => n1624, ZN => n1413);
   U1867 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n1667, B1 => 
                           REGISTERS_18_26_port, B2 => n1655, ZN => n1412);
   U1868 : AND4_X1 port map( A1 => n1415, A2 => n1414, A3 => n1413, A4 => n1412
                           , ZN => n1432);
   U1869 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n1573, B1 => 
                           REGISTERS_31_26_port, B2 => n1556, ZN => n1419);
   U1870 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n1607, B1 => 
                           REGISTERS_27_26_port, B2 => n1590, ZN => n1418);
   U1871 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n1641, B1 => 
                           REGISTERS_30_26_port, B2 => n1624, ZN => n1417);
   U1872 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n1667, B1 => 
                           REGISTERS_26_26_port, B2 => n1655, ZN => n1416);
   U1873 : AND4_X1 port map( A1 => n1419, A2 => n1418, A3 => n1417, A4 => n1416
                           , ZN => n1431);
   U1874 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n1573, B1 => 
                           REGISTERS_7_26_port, B2 => n1556, ZN => n1423);
   U1875 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n1607, B1 => 
                           REGISTERS_3_26_port, B2 => n1590, ZN => n1422);
   U1876 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n1641, B1 => 
                           REGISTERS_6_26_port, B2 => n1624, ZN => n1421);
   U1877 : NAND4_X1 port map( A1 => n1423, A2 => n1422, A3 => n1421, A4 => 
                           n1420, ZN => n1429);
   U1878 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n1573, B1 => 
                           REGISTERS_15_26_port, B2 => n1556, ZN => n1427);
   U1879 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n1607, B1 => 
                           REGISTERS_11_26_port, B2 => n1590, ZN => n1426);
   U1880 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n1641, B1 => 
                           REGISTERS_14_26_port, B2 => n1624, ZN => n1425);
   U1881 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n1667, B1 => 
                           REGISTERS_10_26_port, B2 => n1655, ZN => n1424);
   U1882 : NAND4_X1 port map( A1 => n1427, A2 => n1426, A3 => n1425, A4 => 
                           n1424, ZN => n1428);
   U1883 : AOI22_X1 port map( A1 => n1429, A2 => n1679, B1 => n1428, B2 => 
                           n1675, ZN => n1430);
   U1884 : OAI221_X1 port map( B1 => n1687, B2 => n1432, C1 => n1685, C2 => 
                           n1431, A => n1430, ZN => N264);
   U1885 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n1572, B1 => 
                           REGISTERS_23_27_port, B2 => n1555, ZN => n1436);
   U1886 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n1606, B1 => 
                           REGISTERS_19_27_port, B2 => n1589, ZN => n1435);
   U1887 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n1640, B1 => 
                           REGISTERS_22_27_port, B2 => n1623, ZN => n1434);
   U1888 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n1667, B1 => 
                           REGISTERS_18_27_port, B2 => n1655, ZN => n1433);
   U1889 : AND4_X1 port map( A1 => n1436, A2 => n1435, A3 => n1434, A4 => n1433
                           , ZN => n1453);
   U1890 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n1572, B1 => 
                           REGISTERS_31_27_port, B2 => n1555, ZN => n1440);
   U1891 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n1606, B1 => 
                           REGISTERS_27_27_port, B2 => n1589, ZN => n1439);
   U1892 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n1640, B1 => 
                           REGISTERS_30_27_port, B2 => n1623, ZN => n1438);
   U1893 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n1667, B1 => 
                           REGISTERS_26_27_port, B2 => n1655, ZN => n1437);
   U1894 : AND4_X1 port map( A1 => n1440, A2 => n1439, A3 => n1438, A4 => n1437
                           , ZN => n1452);
   U1895 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n1572, B1 => 
                           REGISTERS_7_27_port, B2 => n1555, ZN => n1444);
   U1896 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n1606, B1 => 
                           REGISTERS_3_27_port, B2 => n1589, ZN => n1443);
   U1897 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n1640, B1 => 
                           REGISTERS_6_27_port, B2 => n1623, ZN => n1442);
   U1898 : NAND4_X1 port map( A1 => n1444, A2 => n1443, A3 => n1442, A4 => 
                           n1441, ZN => n1450);
   U1899 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n1572, B1 => 
                           REGISTERS_15_27_port, B2 => n1555, ZN => n1448);
   U1900 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n1606, B1 => 
                           REGISTERS_11_27_port, B2 => n1589, ZN => n1447);
   U1901 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n1640, B1 => 
                           REGISTERS_14_27_port, B2 => n1623, ZN => n1446);
   U1902 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n1667, B1 => 
                           REGISTERS_10_27_port, B2 => n1655, ZN => n1445);
   U1903 : NAND4_X1 port map( A1 => n1448, A2 => n1447, A3 => n1446, A4 => 
                           n1445, ZN => n1449);
   U1904 : AOI22_X1 port map( A1 => n1450, A2 => n1679, B1 => n1449, B2 => 
                           n1675, ZN => n1451);
   U1905 : OAI221_X1 port map( B1 => n1687, B2 => n1453, C1 => n1685, C2 => 
                           n1452, A => n1451, ZN => N263);
   U1906 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n1572, B1 => 
                           REGISTERS_23_28_port, B2 => n1555, ZN => n1457);
   U1907 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n1606, B1 => 
                           REGISTERS_19_28_port, B2 => n1589, ZN => n1456);
   U1908 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n1640, B1 => 
                           REGISTERS_22_28_port, B2 => n1623, ZN => n1455);
   U1909 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n1666, B1 => 
                           REGISTERS_18_28_port, B2 => n1655, ZN => n1454);
   U1910 : AND4_X1 port map( A1 => n1457, A2 => n1456, A3 => n1455, A4 => n1454
                           , ZN => n1474);
   U1911 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n1572, B1 => 
                           REGISTERS_31_28_port, B2 => n1555, ZN => n1461);
   U1912 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n1606, B1 => 
                           REGISTERS_27_28_port, B2 => n1589, ZN => n1460);
   U1913 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n1640, B1 => 
                           REGISTERS_30_28_port, B2 => n1623, ZN => n1459);
   U1914 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n1666, B1 => 
                           REGISTERS_26_28_port, B2 => n1655, ZN => n1458);
   U1915 : AND4_X1 port map( A1 => n1461, A2 => n1460, A3 => n1459, A4 => n1458
                           , ZN => n1473);
   U1916 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n1572, B1 => 
                           REGISTERS_7_28_port, B2 => n1555, ZN => n1465);
   U1917 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n1606, B1 => 
                           REGISTERS_3_28_port, B2 => n1589, ZN => n1464);
   U1918 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n1640, B1 => 
                           REGISTERS_6_28_port, B2 => n1623, ZN => n1463);
   U1919 : NAND4_X1 port map( A1 => n1465, A2 => n1464, A3 => n1463, A4 => 
                           n1462, ZN => n1471);
   U1920 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n1572, B1 => 
                           REGISTERS_15_28_port, B2 => n1555, ZN => n1469);
   U1921 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n1606, B1 => 
                           REGISTERS_11_28_port, B2 => n1589, ZN => n1468);
   U1922 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n1640, B1 => 
                           REGISTERS_14_28_port, B2 => n1623, ZN => n1467);
   U1923 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n1666, B1 => 
                           REGISTERS_10_28_port, B2 => n1655, ZN => n1466);
   U1924 : NAND4_X1 port map( A1 => n1469, A2 => n1468, A3 => n1467, A4 => 
                           n1466, ZN => n1470);
   U1925 : AOI22_X1 port map( A1 => n1471, A2 => n1679, B1 => n1470, B2 => 
                           n1675, ZN => n1472);
   U1926 : OAI221_X1 port map( B1 => n1687, B2 => n1474, C1 => n1685, C2 => 
                           n1473, A => n1472, ZN => N262);
   U1927 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n1572, B1 => 
                           REGISTERS_23_29_port, B2 => n1555, ZN => n1478);
   U1928 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n1606, B1 => 
                           REGISTERS_19_29_port, B2 => n1589, ZN => n1477);
   U1929 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n1640, B1 => 
                           REGISTERS_22_29_port, B2 => n1623, ZN => n1476);
   U1930 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n1666, B1 => 
                           REGISTERS_18_29_port, B2 => n1654, ZN => n1475);
   U1931 : AND4_X1 port map( A1 => n1478, A2 => n1477, A3 => n1476, A4 => n1475
                           , ZN => n1495);
   U1932 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n1572, B1 => 
                           REGISTERS_31_29_port, B2 => n1555, ZN => n1482);
   U1933 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n1606, B1 => 
                           REGISTERS_27_29_port, B2 => n1589, ZN => n1481);
   U1934 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n1640, B1 => 
                           REGISTERS_30_29_port, B2 => n1623, ZN => n1480);
   U1935 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n1666, B1 => 
                           REGISTERS_26_29_port, B2 => n1654, ZN => n1479);
   U1936 : AND4_X1 port map( A1 => n1482, A2 => n1481, A3 => n1480, A4 => n1479
                           , ZN => n1494);
   U1937 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n1572, B1 => 
                           REGISTERS_7_29_port, B2 => n1555, ZN => n1486);
   U1938 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n1606, B1 => 
                           REGISTERS_3_29_port, B2 => n1589, ZN => n1485);
   U1939 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n1640, B1 => 
                           REGISTERS_6_29_port, B2 => n1623, ZN => n1484);
   U1940 : NAND4_X1 port map( A1 => n1486, A2 => n1485, A3 => n1484, A4 => 
                           n1483, ZN => n1492);
   U1941 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n1572, B1 => 
                           REGISTERS_15_29_port, B2 => n1555, ZN => n1490);
   U1942 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n1606, B1 => 
                           REGISTERS_11_29_port, B2 => n1589, ZN => n1489);
   U1943 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n1640, B1 => 
                           REGISTERS_14_29_port, B2 => n1623, ZN => n1488);
   U1944 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n1666, B1 => 
                           REGISTERS_10_29_port, B2 => n1654, ZN => n1487);
   U1945 : NAND4_X1 port map( A1 => n1490, A2 => n1489, A3 => n1488, A4 => 
                           n1487, ZN => n1491);
   U1946 : AOI22_X1 port map( A1 => n1492, A2 => n1679, B1 => n1491, B2 => 
                           n1675, ZN => n1493);
   U1947 : OAI221_X1 port map( B1 => n1687, B2 => n1495, C1 => n1685, C2 => 
                           n1494, A => n1493, ZN => N261);
   U1948 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n1571, B1 => 
                           REGISTERS_23_30_port, B2 => n1554, ZN => n1499);
   U1949 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n1605, B1 => 
                           REGISTERS_19_30_port, B2 => n1588, ZN => n1498);
   U1950 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n1639, B1 => 
                           REGISTERS_22_30_port, B2 => n1622, ZN => n1497);
   U1951 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n1666, B1 => 
                           REGISTERS_18_30_port, B2 => n1654, ZN => n1496);
   U1952 : AND4_X1 port map( A1 => n1499, A2 => n1498, A3 => n1497, A4 => n1496
                           , ZN => n1516);
   U1953 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n1571, B1 => 
                           REGISTERS_31_30_port, B2 => n1554, ZN => n1503);
   U1954 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n1605, B1 => 
                           REGISTERS_27_30_port, B2 => n1588, ZN => n1502);
   U1955 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n1639, B1 => 
                           REGISTERS_30_30_port, B2 => n1622, ZN => n1501);
   U1956 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n1666, B1 => 
                           REGISTERS_26_30_port, B2 => n1654, ZN => n1500);
   U1957 : AND4_X1 port map( A1 => n1503, A2 => n1502, A3 => n1501, A4 => n1500
                           , ZN => n1515);
   U1958 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n1571, B1 => 
                           REGISTERS_7_30_port, B2 => n1554, ZN => n1507);
   U1959 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n1605, B1 => 
                           REGISTERS_3_30_port, B2 => n1588, ZN => n1506);
   U1960 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n1639, B1 => 
                           REGISTERS_6_30_port, B2 => n1622, ZN => n1505);
   U1961 : NAND4_X1 port map( A1 => n1507, A2 => n1506, A3 => n1505, A4 => 
                           n1504, ZN => n1513);
   U1962 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n1571, B1 => 
                           REGISTERS_15_30_port, B2 => n1554, ZN => n1511);
   U1963 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n1605, B1 => 
                           REGISTERS_11_30_port, B2 => n1588, ZN => n1510);
   U1964 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n1639, B1 => 
                           REGISTERS_14_30_port, B2 => n1622, ZN => n1509);
   U1965 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n1666, B1 => 
                           REGISTERS_10_30_port, B2 => n1654, ZN => n1508);
   U1966 : NAND4_X1 port map( A1 => n1511, A2 => n1510, A3 => n1509, A4 => 
                           n1508, ZN => n1512);
   U1967 : AOI22_X1 port map( A1 => n1513, A2 => n1679, B1 => n1512, B2 => 
                           n1675, ZN => n1514);
   U1968 : OAI221_X1 port map( B1 => n1687, B2 => n1516, C1 => n1685, C2 => 
                           n1515, A => n1514, ZN => N260);
   U1969 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n1571, B1 => 
                           REGISTERS_23_31_port, B2 => n1554, ZN => n1520);
   U1970 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n1605, B1 => 
                           REGISTERS_19_31_port, B2 => n1588, ZN => n1519);
   U1971 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n1639, B1 => 
                           REGISTERS_22_31_port, B2 => n1622, ZN => n1518);
   U1972 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n1666, B1 => 
                           REGISTERS_18_31_port, B2 => n1654, ZN => n1517);
   U1973 : AND4_X1 port map( A1 => n1520, A2 => n1519, A3 => n1518, A4 => n1517
                           , ZN => n1543);
   U1974 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n1571, B1 => 
                           REGISTERS_31_31_port, B2 => n1554, ZN => n1524);
   U1975 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n1605, B1 => 
                           REGISTERS_27_31_port, B2 => n1588, ZN => n1523);
   U1976 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n1639, B1 => 
                           REGISTERS_30_31_port, B2 => n1622, ZN => n1522);
   U1977 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n1666, B1 => 
                           REGISTERS_26_31_port, B2 => n1654, ZN => n1521);
   U1978 : AND4_X1 port map( A1 => n1524, A2 => n1523, A3 => n1522, A4 => n1521
                           , ZN => n1541);
   U1979 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n1571, B1 => 
                           REGISTERS_7_31_port, B2 => n1554, ZN => n1528);
   U1980 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n1605, B1 => 
                           REGISTERS_3_31_port, B2 => n1588, ZN => n1527);
   U1981 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n1639, B1 => 
                           REGISTERS_6_31_port, B2 => n1622, ZN => n1526);
   U1982 : NAND4_X1 port map( A1 => n1528, A2 => n1527, A3 => n1526, A4 => 
                           n1525, ZN => n1537);
   U1983 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n1571, B1 => 
                           REGISTERS_15_31_port, B2 => n1554, ZN => n1534);
   U1984 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n1605, B1 => 
                           REGISTERS_11_31_port, B2 => n1588, ZN => n1533);
   U1985 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n1639, B1 => 
                           REGISTERS_14_31_port, B2 => n1622, ZN => n1532);
   U1986 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n1666, B1 => 
                           REGISTERS_10_31_port, B2 => n1654, ZN => n1531);
   U1987 : NAND4_X1 port map( A1 => n1534, A2 => n1533, A3 => n1532, A4 => 
                           n1531, ZN => n1535);
   U1988 : AOI22_X1 port map( A1 => n1679, A2 => n1537, B1 => n1675, B2 => 
                           n1535, ZN => n1539);
   U1989 : OAI221_X1 port map( B1 => n1543, B2 => n1687, C1 => n1541, C2 => 
                           n1685, A => n1539, ZN => N259);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CWBU is

   port( CLOCK : in std_logic;  ALU_OP : in std_logic_vector (0 to 4);  PSW : 
         in std_logic_vector (6 downto 0);  COND_SEL : out std_logic_vector (1 
         downto 0);  CWB_SEL : in std_logic_vector (1 downto 0);  CWB_MUW_SEL :
         out std_logic_vector (1 downto 0));

end CWBU;

architecture SYN_BEHAVIORAL of CWBU is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal ALUPIPE_4_port, ALUPIPE_2_port, ALUPIPE_1_port, ALUPIPE_0_port, n1, 
      n3, n4, n5, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n2, n6, n7, n8, n9, n10, n_1705, n_1706 : std_logic;

begin
   
   ALUPIPE_reg_2_inst : DFF_X1 port map( D => ALU_OP(2), CK => CLOCK, Q => 
                           ALUPIPE_2_port, QN => n_1705);
   U24 : NAND3_X1 port map( A1 => n10, A2 => n2, A3 => n11, ZN => 
                           CWB_MUW_SEL(1));
   U25 : NAND3_X1 port map( A1 => n5, A2 => n4, A3 => PSW(0), ZN => n23);
   ALUPIPE_reg_3_inst : DFF_X1 port map( D => ALU_OP(1), CK => CLOCK, Q => 
                           n_1706, QN => n3);
   ALUPIPE_reg_4_inst : DFF_X1 port map( D => ALU_OP(0), CK => CLOCK, Q => 
                           ALUPIPE_4_port, QN => n1);
   ALUPIPE_reg_1_inst : DFF_X1 port map( D => ALU_OP(3), CK => CLOCK, Q => 
                           ALUPIPE_1_port, QN => n4);
   ALUPIPE_reg_0_inst : DFF_X1 port map( D => ALU_OP(4), CK => CLOCK, Q => 
                           ALUPIPE_0_port, QN => n5);
   U3 : INV_X1 port map( A => n14, ZN => n2);
   U4 : INV_X1 port map( A => CWB_SEL(1), ZN => n10);
   U5 : AOI221_X1 port map( B1 => PSW(1), B2 => n17, C1 => PSW(3), C2 => n13, A
                           => n22, ZN => n21);
   U6 : OAI21_X1 port map( B1 => n19, B2 => n8, A => n23, ZN => n22);
   U7 : INV_X1 port map( A => PSW(2), ZN => n8);
   U8 : AOI221_X1 port map( B1 => n17, B2 => n9, C1 => n13, C2 => n7, A => n18,
                           ZN => n16);
   U9 : INV_X1 port map( A => PSW(1), ZN => n9);
   U10 : INV_X1 port map( A => PSW(3), ZN => n7);
   U11 : OAI21_X1 port map( B1 => PSW(2), B2 => n19, A => n20, ZN => n18);
   U12 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n13);
   U13 : NOR2_X1 port map( A1 => n4, A2 => ALUPIPE_0_port, ZN => n17);
   U14 : AND2_X1 port map( A1 => CWB_SEL(0), A2 => n12, ZN => CWB_MUW_SEL(0));
   U15 : OAI211_X1 port map( C1 => n13, C2 => n14, A => n1, B => n15, ZN => n12
                           );
   U16 : OAI22_X1 port map( A1 => n21, A2 => n2, B1 => n11, B2 => n6, ZN => 
                           COND_SEL(0));
   U17 : OAI22_X1 port map( A1 => n16, A2 => n2, B1 => PSW(5), B2 => n11, ZN =>
                           COND_SEL(1));
   U18 : NAND2_X1 port map( A1 => ALUPIPE_0_port, A2 => n4, ZN => n19);
   U19 : OR3_X1 port map( A1 => ALUPIPE_1_port, A2 => PSW(0), A3 => 
                           ALUPIPE_0_port, ZN => n20);
   U20 : INV_X1 port map( A => PSW(5), ZN => n6);
   U21 : XNOR2_X1 port map( A => n3, B => ALUPIPE_2_port, ZN => n15);
   U22 : NAND4_X1 port map( A1 => ALUPIPE_2_port, A2 => n13, A3 => n3, A4 => n1
                           , ZN => n11);
   U23 : NOR3_X1 port map( A1 => ALUPIPE_2_port, A2 => ALUPIPE_4_port, A3 => n3
                           , ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 is

   port( clock, rst : in std_logic;  address : in std_logic_vector (31 downto 
         0);  d_in, w_en : in std_logic;  d_out : out std_logic);

end BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0;

architecture SYN_Behavioral of BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal BHT_0_1_port, BHT_0_0_port, BHT_1_1_port, BHT_1_0_port, BHT_2_1_port,
      BHT_2_0_port, BHT_3_1_port, BHT_3_0_port, BHT_4_1_port, BHT_4_0_port, 
      BHT_5_1_port, BHT_5_0_port, BHT_6_1_port, BHT_6_0_port, BHT_7_1_port, 
      BHT_7_0_port, N55, n24, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
      n78, n79, n80, n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55_port
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n_1707, 
      n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714 : std_logic;

begin
   d_out <= N55;
   
   BHT_reg_7_1_inst : DFFR_X1 port map( D => n67, CK => n66, RN => n17, Q => 
                           BHT_7_1_port, QN => n_1707);
   BHT_reg_5_0_inst : DFFR_X1 port map( D => n71, CK => n66, RN => n17, Q => 
                           BHT_5_0_port, QN => n_1708);
   BHT_reg_3_1_inst : DFFR_X1 port map( D => n76, CK => n66, RN => n17, Q => 
                           BHT_3_1_port, QN => n_1709);
   BHT_reg_3_0_inst : DFFR_X1 port map( D => n75, CK => n66, RN => n17, Q => 
                           BHT_3_0_port, QN => n_1710);
   BHT_reg_2_1_inst : DFFR_X1 port map( D => n78, CK => n66, RN => n17, Q => 
                           BHT_2_1_port, QN => n_1711);
   BHT_reg_2_0_inst : DFFR_X1 port map( D => n77, CK => n66, RN => n17, Q => 
                           BHT_2_0_port, QN => n_1712);
   BHT_reg_4_0_inst : DFFR_X1 port map( D => n73, CK => n66, RN => n17, Q => 
                           BHT_4_0_port, QN => n_1713);
   BHT_reg_6_1_inst : DFFR_X1 port map( D => n70, CK => n66, RN => n17, Q => 
                           BHT_6_1_port, QN => n_1714);
   BHT_reg_7_0_inst : DFFR_X1 port map( D => n68, CK => n66, RN => n17, Q => 
                           BHT_7_0_port, QN => n24);
   BHT_reg_1_1_inst : DFFR_X1 port map( D => n80, CK => n66, RN => n17, Q => 
                           BHT_1_1_port, QN => n29);
   BHT_reg_1_0_inst : DFFR_X1 port map( D => n79, CK => n66, RN => n17, Q => 
                           BHT_1_0_port, QN => n19);
   BHT_reg_5_1_inst : DFFR_X1 port map( D => n72, CK => n66, RN => n17, Q => 
                           BHT_5_1_port, QN => n33);
   BHT_reg_4_1_inst : DFFR_X1 port map( D => n74, CK => n66, RN => n17, Q => 
                           BHT_4_1_port, QN => n35);
   BHT_reg_0_1_inst : DFFR_X1 port map( D => n82, CK => n66, RN => n17, Q => 
                           BHT_0_1_port, QN => n30);
   BHT_reg_0_0_inst : DFFR_X1 port map( D => n81, CK => n66, RN => n17, Q => 
                           BHT_0_0_port, QN => n20);
   BHT_reg_6_0_inst : DFFR_X1 port map( D => n69, CK => n66, RN => n17, Q => 
                           BHT_6_0_port, QN => n26);
   U3 : CLKBUF_X1 port map( A => w_en, Z => n15);
   U4 : AND2_X1 port map( A1 => n9, A2 => n2, ZN => n1);
   U5 : INV_X1 port map( A => rst, ZN => n17);
   U6 : INV_X1 port map( A => n15, ZN => n16);
   U7 : NAND2_X1 port map( A1 => N55, A2 => n56, ZN => n48);
   U8 : AND2_X1 port map( A1 => n51, A2 => n50, ZN => n2);
   U9 : AND2_X1 port map( A1 => n14, A2 => n2, ZN => n3);
   U10 : AND2_X1 port map( A1 => n2, A2 => n13, ZN => n4);
   U11 : AND2_X1 port map( A1 => n13, A2 => n12, ZN => n5);
   U12 : AND2_X1 port map( A1 => n14, A2 => n12, ZN => n6);
   U13 : AND2_X1 port map( A1 => n9, A2 => n12, ZN => n7);
   U14 : XNOR2_X1 port map( A => n54, B => n8, ZN => n65);
   U15 : XNOR2_X1 port map( A => d_in, B => n57, ZN => n8);
   U16 : AND2_X1 port map( A1 => n63, A2 => n62, ZN => n9);
   U17 : AND3_X1 port map( A1 => address(2), A2 => address(1), A3 => n2, ZN => 
                           n10);
   U18 : NAND2_X1 port map( A1 => n39, A2 => n38, ZN => n47);
   U19 : INV_X1 port map( A => n44, ZN => n38);
   U20 : AND2_X1 port map( A1 => address(1), A2 => address(0), ZN => n11);
   U21 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => n46);
   U22 : AND2_X1 port map( A1 => n51, A2 => address(0), ZN => n12);
   U23 : AND2_X1 port map( A1 => address(1), A2 => n63, ZN => n13);
   U24 : AND2_X1 port map( A1 => address(2), A2 => n62, ZN => n14);
   U25 : OAI221_X1 port map( B1 => n36, B2 => n20, C1 => n34, C2 => n19, A => 
                           n18, ZN => n37);
   U26 : OAI221_X1 port map( B1 => n36, B2 => n30, C1 => n34, C2 => n29, A => 
                           n28, ZN => n39);
   U27 : OAI221_X1 port map( B1 => n36, B2 => n35, C1 => n34, C2 => n33, A => 
                           n32, ZN => n42);
   U28 : INV_X1 port map( A => n43, ZN => n41);
   U29 : AOI21_X1 port map( B1 => n49, B2 => n48, A => n16, ZN => n51);
   U30 : INV_X1 port map( A => address(1), ZN => n62);
   U31 : INV_X1 port map( A => address(0), ZN => n50);
   U32 : NAND2_X1 port map( A1 => n62, A2 => n50, ZN => n36);
   U33 : NAND2_X1 port map( A1 => address(0), A2 => n62, ZN => n34);
   U34 : NAND2_X1 port map( A1 => address(1), A2 => n50, ZN => n27);
   U35 : INV_X1 port map( A => n27, ZN => n31);
   U36 : AOI22_X1 port map( A1 => BHT_2_0_port, A2 => n31, B1 => BHT_3_0_port, 
                           B2 => n11, ZN => n18);
   U37 : NAND3_X1 port map( A1 => BHT_7_0_port, A2 => address(1), A3 => 
                           address(0), ZN => n25);
   U38 : INV_X1 port map( A => n36, ZN => n22);
   U39 : INV_X1 port map( A => n34, ZN => n21);
   U40 : AOI22_X1 port map( A1 => BHT_4_0_port, A2 => n22, B1 => BHT_5_0_port, 
                           B2 => n21, ZN => n23);
   U41 : OAI211_X1 port map( C1 => n27, C2 => n26, A => n25, B => n23, ZN => 
                           n40);
   U42 : MUX2_X1 port map( A => n37, B => n40, S => address(2), Z => n54);
   U43 : AOI22_X1 port map( A1 => BHT_2_1_port, A2 => n31, B1 => BHT_3_1_port, 
                           B2 => n11, ZN => n28);
   U44 : AOI22_X1 port map( A1 => BHT_6_1_port, A2 => n31, B1 => BHT_7_1_port, 
                           B2 => n11, ZN => n32);
   U45 : MUX2_X1 port map( A => n39, B => n42, S => address(2), Z => N55);
   U46 : INV_X1 port map( A => N55, ZN => n57);
   U47 : INV_X1 port map( A => address(2), ZN => n63);
   U48 : NAND2_X1 port map( A1 => n37, A2 => n63, ZN => n44);
   U49 : NAND2_X1 port map( A1 => n40, A2 => address(2), ZN => n43);
   U50 : INV_X1 port map( A => d_in, ZN => n56);
   U51 : NAND3_X1 port map( A1 => n44, A2 => n56, A3 => n43, ZN => n45);
   U52 : NAND3_X1 port map( A1 => n47, A2 => n46, A3 => n45, ZN => n49);
   U53 : MUX2_X1 port map( A => BHT_4_1_port, B => n65, S => n3, Z => n74);
   U54 : INV_X1 port map( A => clock, ZN => n66);
   U55 : MUX2_X1 port map( A => BHT_5_1_port, B => n65, S => n6, Z => n72);
   U56 : MUX2_X1 port map( A => BHT_6_1_port, B => n65, S => n10, Z => n70);
   U57 : NAND3_X1 port map( A1 => n15, A2 => address(2), A3 => n11, ZN => 
                           n55_port);
   U58 : INV_X1 port map( A => n55_port, ZN => n61);
   U59 : OAI211_X1 port map( C1 => N55, C2 => n54, A => d_in, B => n61, ZN => 
                           n53);
   U60 : OAI21_X1 port map( B1 => n54, B2 => n55_port, A => BHT_7_1_port, ZN =>
                           n52);
   U61 : NAND2_X1 port map( A1 => n53, A2 => n52, ZN => n67);
   U62 : INV_X1 port map( A => n54, ZN => n64);
   U63 : MUX2_X1 port map( A => BHT_4_0_port, B => n64, S => n3, Z => n73);
   U64 : MUX2_X1 port map( A => BHT_5_0_port, B => n64, S => n6, Z => n71);
   U65 : MUX2_X1 port map( A => BHT_6_0_port, B => n64, S => n10, Z => n69);
   U66 : AOI21_X1 port map( B1 => n57, B2 => n56, A => n55_port, ZN => n58);
   U67 : OAI21_X1 port map( B1 => BHT_7_0_port, B2 => n58, A => n64, ZN => n60)
                           ;
   U68 : NAND3_X1 port map( A1 => d_in, A2 => BHT_7_0_port, A3 => N55, ZN => 
                           n59);
   U69 : OAI211_X1 port map( C1 => n24, C2 => n61, A => n60, B => n59, ZN => 
                           n68);
   U70 : MUX2_X1 port map( A => BHT_0_0_port, B => n64, S => n1, Z => n81);
   U71 : MUX2_X1 port map( A => BHT_1_0_port, B => n64, S => n7, Z => n79);
   U72 : MUX2_X1 port map( A => BHT_2_0_port, B => n64, S => n4, Z => n77);
   U73 : MUX2_X1 port map( A => BHT_3_0_port, B => n64, S => n5, Z => n75);
   U74 : MUX2_X1 port map( A => BHT_0_1_port, B => n65, S => n1, Z => n82);
   U75 : MUX2_X1 port map( A => BHT_1_1_port, B => n65, S => n7, Z => n80);
   U76 : MUX2_X1 port map( A => BHT_2_1_port, B => n65, S => n4, Z => n78);
   U77 : MUX2_X1 port map( A => BHT_3_1_port, B => n65, S => n5, Z => n76);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HDU_IR_SIZE32 is

   port( clk, rst : in std_logic;  IR : in std_logic_vector (31 downto 0);  
         STALL_CODE : out std_logic_vector (1 downto 0);  IF_STALL, ID_STALL, 
         EX_STALL, MEM_STALL, WB_STALL : out std_logic);

end HDU_IR_SIZE32;

architecture SYN_behavioural of HDU_IR_SIZE32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component HDU_IR_SIZE32_DW01_dec_1
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal STALL_CODE_1_port, IF_STALL_port, EX_STALL_port, cnt_mul_31_port, 
      cnt_mul_30_port, cnt_mul_29_port, cnt_mul_28_port, cnt_mul_27_port, 
      cnt_mul_26_port, cnt_mul_25_port, cnt_mul_24_port, cnt_mul_23_port, 
      cnt_mul_22_port, cnt_mul_21_port, cnt_mul_20_port, cnt_mul_19_port, 
      cnt_mul_18_port, cnt_mul_17_port, cnt_mul_16_port, cnt_mul_15_port, 
      cnt_mul_14_port, cnt_mul_13_port, cnt_mul_12_port, cnt_mul_11_port, 
      cnt_mul_10_port, cnt_mul_9_port, cnt_mul_8_port, cnt_mul_7_port, 
      cnt_mul_6_port, cnt_mul_5_port, cnt_mul_4_port, cnt_mul_3_port, 
      cnt_mul_2_port, cnt_mul_1_port, cnt_mul_0_port, N154, N155, N156, N157, 
      N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, 
      N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, 
      N182, N183, N184, n99, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n125, n126, n127, n128, 
      n149, n150, n151, n152, n153, n154_port, n155_port, n156_port, n157_port,
      n158_port, n159_port, n169_port, n170_port, n171_port, n172_port, 
      n173_port, n174_port, n175_port, n176_port, n177_port, n178_port, 
      n179_port, n180_port, n181_port, n182_port, n183_port, n184_port, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n202, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
      n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n100, n117, n118, n119, n120, n121, n122, n123, n124, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, STALL_CODE_0_port, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726 : std_logic;

begin
   STALL_CODE <= ( STALL_CODE_1_port, STALL_CODE_0_port );
   IF_STALL <= IF_STALL_port;
   ID_STALL <= IF_STALL_port;
   EX_STALL <= EX_STALL_port;
   MEM_STALL <= EX_STALL_port;
   WB_STALL <= EX_STALL_port;
   
   IR_EX_reg_28_inst : DFFR_X1 port map( D => n156_port, CK => clk, RN => n17, 
                           Q => n145, QN => n2);
   IR_EX_reg_27_inst : DFFR_X1 port map( D => n155_port, CK => clk, RN => n17, 
                           Q => n144, QN => n1);
   IR_EX_reg_20_inst : DFFR_X1 port map( D => n153, CK => clk, RN => n17, Q => 
                           n140, QN => n_1720);
   IR_EX_reg_19_inst : DFFR_X1 port map( D => n152, CK => clk, RN => n17, Q => 
                           n139, QN => n_1721);
   IR_EX_reg_18_inst : DFFR_X1 port map( D => n151, CK => clk, RN => n17, Q => 
                           n138, QN => n_1722);
   IR_EX_reg_17_inst : DFFR_X1 port map( D => n150, CK => clk, RN => n17, Q => 
                           n137, QN => n7);
   IR_EX_reg_16_inst : DFFR_X1 port map( D => n149, CK => clk, RN => n17, Q => 
                           n136, QN => n_1723);
   r100 : HDU_IR_SIZE32_DW01_dec_1 port map( A(31) => cnt_mul_31_port, A(30) =>
                           cnt_mul_30_port, A(29) => cnt_mul_29_port, A(28) => 
                           cnt_mul_28_port, A(27) => cnt_mul_27_port, A(26) => 
                           cnt_mul_26_port, A(25) => cnt_mul_25_port, A(24) => 
                           cnt_mul_24_port, A(23) => cnt_mul_23_port, A(22) => 
                           cnt_mul_22_port, A(21) => cnt_mul_21_port, A(20) => 
                           cnt_mul_20_port, A(19) => cnt_mul_19_port, A(18) => 
                           cnt_mul_18_port, A(17) => cnt_mul_17_port, A(16) => 
                           cnt_mul_16_port, A(15) => cnt_mul_15_port, A(14) => 
                           cnt_mul_14_port, A(13) => cnt_mul_13_port, A(12) => 
                           cnt_mul_12_port, A(11) => cnt_mul_11_port, A(10) => 
                           cnt_mul_10_port, A(9) => cnt_mul_9_port, A(8) => 
                           cnt_mul_8_port, A(7) => cnt_mul_7_port, A(6) => 
                           cnt_mul_6_port, A(5) => cnt_mul_5_port, A(4) => 
                           cnt_mul_4_port, A(3) => cnt_mul_3_port, A(2) => 
                           cnt_mul_2_port, A(1) => cnt_mul_1_port, A(0) => 
                           cnt_mul_0_port, SUM(31) => N184, SUM(30) => N183, 
                           SUM(29) => N182, SUM(28) => N181, SUM(27) => N180, 
                           SUM(26) => N179, SUM(25) => N178, SUM(24) => N177, 
                           SUM(23) => N176, SUM(22) => N175, SUM(21) => N174, 
                           SUM(20) => N173, SUM(19) => N172, SUM(18) => N171, 
                           SUM(17) => N170, SUM(16) => N169, SUM(15) => N168, 
                           SUM(14) => N167, SUM(13) => N166, SUM(12) => N165, 
                           SUM(11) => N164, SUM(10) => N163, SUM(9) => N162, 
                           SUM(8) => N161, SUM(7) => N160, SUM(6) => N159, 
                           SUM(5) => N158, SUM(4) => N157, SUM(3) => N156, 
                           SUM(2) => N155, SUM(1) => N154, SUM(0) => n_1724);
   STALL_MUL_reg : DFF_X1 port map( D => n3, CK => clk, Q => EX_STALL_port, QN 
                           => n199);
   cnt_mul_reg_7_inst : DFF_X1 port map( D => n192, CK => clk, Q => 
                           cnt_mul_7_port, QN => n106);
   cnt_mul_reg_6_inst : DFF_X1 port map( D => n193, CK => clk, Q => 
                           cnt_mul_6_port, QN => n105);
   cnt_mul_reg_5_inst : DFF_X1 port map( D => n194, CK => clk, Q => 
                           cnt_mul_5_port, QN => n104);
   cnt_mul_reg_4_inst : DFF_X1 port map( D => n195, CK => clk, Q => 
                           cnt_mul_4_port, QN => n103);
   cnt_mul_reg_3_inst : DFF_X1 port map( D => n196, CK => clk, Q => 
                           cnt_mul_3_port, QN => n102);
   cnt_mul_reg_2_inst : DFF_X1 port map( D => n197, CK => clk, Q => 
                           cnt_mul_2_port, QN => n101);
   cnt_mul_reg_30_inst : DFF_X1 port map( D => n169_port, CK => clk, Q => 
                           cnt_mul_30_port, QN => n31);
   cnt_mul_reg_29_inst : DFF_X1 port map( D => n170_port, CK => clk, Q => 
                           cnt_mul_29_port, QN => n128);
   cnt_mul_reg_28_inst : DFF_X1 port map( D => n171_port, CK => clk, Q => 
                           cnt_mul_28_port, QN => n127);
   cnt_mul_reg_31_inst : DFF_X1 port map( D => n198, CK => clk, Q => 
                           cnt_mul_31_port, QN => n99);
   cnt_mul_reg_13_inst : DFF_X1 port map( D => n186, CK => clk, Q => 
                           cnt_mul_13_port, QN => n112);
   cnt_mul_reg_12_inst : DFF_X1 port map( D => n187, CK => clk, Q => 
                           cnt_mul_12_port, QN => n111);
   cnt_mul_reg_11_inst : DFF_X1 port map( D => n188, CK => clk, Q => 
                           cnt_mul_11_port, QN => n110);
   cnt_mul_reg_10_inst : DFF_X1 port map( D => n189, CK => clk, Q => 
                           cnt_mul_10_port, QN => n109);
   cnt_mul_reg_9_inst : DFF_X1 port map( D => n190, CK => clk, Q => 
                           cnt_mul_9_port, QN => n108);
   cnt_mul_reg_8_inst : DFF_X1 port map( D => n191, CK => clk, Q => 
                           cnt_mul_8_port, QN => n107);
   cnt_mul_reg_27_inst : DFF_X1 port map( D => n172_port, CK => clk, Q => 
                           cnt_mul_27_port, QN => n126);
   cnt_mul_reg_26_inst : DFF_X1 port map( D => n173_port, CK => clk, Q => 
                           cnt_mul_26_port, QN => n125);
   cnt_mul_reg_25_inst : DFF_X1 port map( D => n174_port, CK => clk, Q => 
                           cnt_mul_25_port, QN => n33);
   cnt_mul_reg_24_inst : DFF_X1 port map( D => n175_port, CK => clk, Q => 
                           cnt_mul_24_port, QN => n34);
   cnt_mul_reg_23_inst : DFF_X1 port map( D => n176_port, CK => clk, Q => 
                           cnt_mul_23_port, QN => n35);
   cnt_mul_reg_22_inst : DFF_X1 port map( D => n177_port, CK => clk, Q => 
                           cnt_mul_22_port, QN => n36);
   cnt_mul_reg_21_inst : DFF_X1 port map( D => n178_port, CK => clk, Q => 
                           cnt_mul_21_port, QN => n37);
   cnt_mul_reg_20_inst : DFF_X1 port map( D => n179_port, CK => clk, Q => 
                           cnt_mul_20_port, QN => n38);
   cnt_mul_reg_19_inst : DFF_X1 port map( D => n180_port, CK => clk, Q => 
                           cnt_mul_19_port, QN => n39);
   cnt_mul_reg_18_inst : DFF_X1 port map( D => n181_port, CK => clk, Q => 
                           cnt_mul_18_port, QN => n40);
   cnt_mul_reg_17_inst : DFF_X1 port map( D => n182_port, CK => clk, Q => 
                           cnt_mul_17_port, QN => n116);
   cnt_mul_reg_16_inst : DFF_X1 port map( D => n183_port, CK => clk, Q => 
                           cnt_mul_16_port, QN => n115);
   cnt_mul_reg_15_inst : DFF_X1 port map( D => n184_port, CK => clk, Q => 
                           cnt_mul_15_port, QN => n114);
   cnt_mul_reg_14_inst : DFF_X1 port map( D => n185, CK => clk, Q => 
                           cnt_mul_14_port, QN => n113);
   cnt_mul_reg_1_inst : DFF_X1 port map( D => n200, CK => clk, Q => 
                           cnt_mul_1_port, QN => n32);
   cnt_mul_reg_0_inst : DFF_X1 port map( D => n202, CK => clk, Q => 
                           cnt_mul_0_port, QN => n30);
   IR_EX_reg_31_inst : DFFR_X1 port map( D => n159_port, CK => clk, RN => n17, 
                           Q => n146, QN => n_1725);
   IR_EX_reg_30_inst : DFFR_X1 port map( D => n158_port, CK => clk, RN => n17, 
                           Q => n142, QN => n133);
   IR_EX_reg_29_inst : DFFR_X1 port map( D => n157_port, CK => clk, RN => n17, 
                           Q => n143, QN => n132);
   IR_EX_reg_26_inst : DFFR_X1 port map( D => n154_port, CK => clk, RN => n17, 
                           Q => n141, QN => n_1726);
   U3 : BUF_X1 port map( A => n3, Z => n16);
   U4 : CLKBUF_X1 port map( A => n4, Z => n12);
   U5 : BUF_X1 port map( A => n4, Z => n11);
   U6 : AND2_X1 port map( A1 => n199, A2 => n45, ZN => n4);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n13);
   U9 : INV_X1 port map( A => n11, ZN => n8);
   U10 : CLKBUF_X1 port map( A => n16, Z => n15);
   U11 : INV_X1 port map( A => n11, ZN => n9);
   U12 : INV_X1 port map( A => n11, ZN => n10);
   U13 : INV_X1 port map( A => rst, ZN => n17);
   U14 : AND2_X1 port map( A1 => n76, A2 => n8, ZN => n3);
   U15 : NAND4_X1 port map( A1 => n134, A2 => n146, A3 => n133, A4 => n132, ZN 
                           => n135);
   U16 : AOI21_X1 port map( B1 => n131, B2 => n130, A => n129, ZN => n134);
   U17 : XNOR2_X1 port map( A => n136, B => IR(21), ZN => n96);
   U18 : NOR2_X1 port map( A1 => n5, A2 => n94, ZN => n95);
   U19 : OAI21_X1 port map( B1 => IR(30), B2 => n85, A => n84, ZN => n87);
   U20 : NAND2_X1 port map( A1 => IR(28), A2 => IR(26), ZN => n84);
   U21 : INV_X1 port map( A => n118, ZN => n85);
   U22 : XNOR2_X1 port map( A => IR(24), B => n139, ZN => n92);
   U23 : XNOR2_X1 port map( A => IR(23), B => n138, ZN => n91);
   U24 : XNOR2_X1 port map( A => IR(25), B => n140, ZN => n93);
   U25 : NOR4_X1 port map( A1 => n119, A2 => IR(29), A3 => IR(27), A4 => n118, 
                           ZN => n123);
   U26 : AND2_X1 port map( A1 => n121, A2 => n120, ZN => n122);
   U27 : NOR2_X1 port map( A1 => n6, A2 => n117, ZN => n124);
   U28 : NAND2_X1 port map( A1 => n100, A2 => n98, ZN => n117);
   U29 : XNOR2_X1 port map( A => IR(20), B => n140, ZN => n98);
   U30 : XNOR2_X1 port map( A => IR(16), B => n136, ZN => n100);
   U31 : XNOR2_X1 port map( A => n7, B => IR(22), ZN => n5);
   U32 : XNOR2_X1 port map( A => IR(17), B => n7, ZN => n6);
   U33 : XNOR2_X1 port map( A => n139, B => IR(19), ZN => n120);
   U34 : XNOR2_X1 port map( A => n138, B => IR(18), ZN => n121);
   U35 : INV_X1 port map( A => IR(29), ZN => n88);
   U36 : AOI21_X1 port map( B1 => n141, B2 => n2, A => n1, ZN => n129);
   U37 : XNOR2_X1 port map( A => n8, B => cnt_mul_0_port, ZN => n80);
   U38 : NAND3_X1 port map( A1 => IR(3), A2 => IR(26), A3 => IR(2), ZN => n19);
   U39 : INV_X1 port map( A => IR(1), ZN => n18);
   U40 : NOR3_X1 port map( A1 => n19, A2 => IR(0), A3 => n18, ZN => n24);
   U41 : NOR4_X1 port map( A1 => IR(7), A2 => IR(6), A3 => IR(5), A4 => IR(4), 
                           ZN => n23);
   U42 : NOR4_X1 port map( A1 => IR(27), A2 => IR(10), A3 => IR(9), A4 => IR(8)
                           , ZN => n22);
   U43 : INV_X1 port map( A => IR(30), ZN => n20);
   U44 : INV_X1 port map( A => IR(31), ZN => n90);
   U45 : NAND2_X1 port map( A1 => n20, A2 => n90, ZN => n119);
   U46 : NOR3_X1 port map( A1 => n119, A2 => IR(29), A3 => IR(28), ZN => n21);
   U47 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n45);
   U48 : NOR4_X1 port map( A1 => cnt_mul_5_port, A2 => cnt_mul_4_port, A3 => 
                           cnt_mul_3_port, A4 => cnt_mul_2_port, ZN => n28);
   U49 : NOR4_X1 port map( A1 => cnt_mul_9_port, A2 => cnt_mul_8_port, A3 => 
                           cnt_mul_7_port, A4 => cnt_mul_6_port, ZN => n27);
   U50 : NOR4_X1 port map( A1 => cnt_mul_13_port, A2 => cnt_mul_12_port, A3 => 
                           cnt_mul_11_port, A4 => cnt_mul_10_port, ZN => n26);
   U51 : NOR4_X1 port map( A1 => cnt_mul_17_port, A2 => cnt_mul_16_port, A3 => 
                           cnt_mul_15_port, A4 => cnt_mul_14_port, ZN => n25);
   U52 : NAND4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n44);
   U53 : NOR4_X1 port map( A1 => cnt_mul_29_port, A2 => cnt_mul_28_port, A3 => 
                           cnt_mul_27_port, A4 => cnt_mul_26_port, ZN => n29);
   U54 : NAND4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n43);
   U55 : NAND4_X1 port map( A1 => n36, A2 => n35, A3 => n34, A4 => n33, ZN => 
                           n42);
   U56 : NAND4_X1 port map( A1 => n40, A2 => n39, A3 => n38, A4 => n37, ZN => 
                           n41);
   U57 : NOR4_X1 port map( A1 => n44, A2 => n43, A3 => n42, A4 => n41, ZN => 
                           n46);
   U58 : OAI21_X1 port map( B1 => cnt_mul_31_port, B2 => n46, A => n45, ZN => 
                           n76);
   U59 : NAND2_X1 port map( A1 => N184, A2 => n13, ZN => n47);
   U60 : OAI21_X1 port map( B1 => n99, B2 => n8, A => n47, ZN => n198);
   U61 : NAND2_X1 port map( A1 => N183, A2 => n13, ZN => n48);
   U62 : OAI21_X1 port map( B1 => n31, B2 => n10, A => n48, ZN => n169_port);
   U63 : NAND2_X1 port map( A1 => N182, A2 => n13, ZN => n49);
   U64 : OAI21_X1 port map( B1 => n128, B2 => n10, A => n49, ZN => n170_port);
   U65 : NAND2_X1 port map( A1 => N181, A2 => n13, ZN => n50);
   U66 : OAI21_X1 port map( B1 => n127, B2 => n10, A => n50, ZN => n171_port);
   U67 : NAND2_X1 port map( A1 => N180, A2 => n13, ZN => n51);
   U68 : OAI21_X1 port map( B1 => n126, B2 => n9, A => n51, ZN => n172_port);
   U69 : NAND2_X1 port map( A1 => N179, A2 => n13, ZN => n52);
   U70 : OAI21_X1 port map( B1 => n125, B2 => n9, A => n52, ZN => n173_port);
   U71 : NAND2_X1 port map( A1 => N178, A2 => n13, ZN => n53);
   U72 : OAI21_X1 port map( B1 => n33, B2 => n9, A => n53, ZN => n174_port);
   U73 : NAND2_X1 port map( A1 => N177, A2 => n13, ZN => n54);
   U74 : OAI21_X1 port map( B1 => n34, B2 => n9, A => n54, ZN => n175_port);
   U75 : NAND2_X1 port map( A1 => N176, A2 => n13, ZN => n55);
   U76 : OAI21_X1 port map( B1 => n35, B2 => n9, A => n55, ZN => n176_port);
   U77 : NAND2_X1 port map( A1 => N175, A2 => n13, ZN => n56);
   U78 : OAI21_X1 port map( B1 => n36, B2 => n9, A => n56, ZN => n177_port);
   U79 : NAND2_X1 port map( A1 => N174, A2 => n13, ZN => n57);
   U80 : OAI21_X1 port map( B1 => n37, B2 => n9, A => n57, ZN => n178_port);
   U81 : NAND2_X1 port map( A1 => N173, A2 => n13, ZN => n58);
   U82 : OAI21_X1 port map( B1 => n38, B2 => n9, A => n58, ZN => n179_port);
   U83 : NAND2_X1 port map( A1 => N172, A2 => n14, ZN => n59);
   U84 : OAI21_X1 port map( B1 => n39, B2 => n9, A => n59, ZN => n180_port);
   U85 : NAND2_X1 port map( A1 => N171, A2 => n14, ZN => n60);
   U86 : OAI21_X1 port map( B1 => n40, B2 => n9, A => n60, ZN => n181_port);
   U87 : NAND2_X1 port map( A1 => N170, A2 => n14, ZN => n61);
   U88 : OAI21_X1 port map( B1 => n116, B2 => n9, A => n61, ZN => n182_port);
   U89 : NAND2_X1 port map( A1 => N169, A2 => n14, ZN => n62);
   U90 : OAI21_X1 port map( B1 => n115, B2 => n9, A => n62, ZN => n183_port);
   U91 : NAND2_X1 port map( A1 => N168, A2 => n14, ZN => n63);
   U92 : OAI21_X1 port map( B1 => n114, B2 => n9, A => n63, ZN => n184_port);
   U93 : NAND2_X1 port map( A1 => N167, A2 => n14, ZN => n64);
   U94 : OAI21_X1 port map( B1 => n113, B2 => n9, A => n64, ZN => n185);
   U95 : NAND2_X1 port map( A1 => N166, A2 => n14, ZN => n65);
   U96 : OAI21_X1 port map( B1 => n112, B2 => n8, A => n65, ZN => n186);
   U97 : NAND2_X1 port map( A1 => N165, A2 => n14, ZN => n66);
   U98 : OAI21_X1 port map( B1 => n111, B2 => n8, A => n66, ZN => n187);
   U99 : NAND2_X1 port map( A1 => N164, A2 => n14, ZN => n67);
   U100 : OAI21_X1 port map( B1 => n110, B2 => n8, A => n67, ZN => n188);
   U101 : NAND2_X1 port map( A1 => N163, A2 => n14, ZN => n68);
   U102 : OAI21_X1 port map( B1 => n109, B2 => n8, A => n68, ZN => n189);
   U103 : NAND2_X1 port map( A1 => N162, A2 => n14, ZN => n69);
   U104 : OAI21_X1 port map( B1 => n108, B2 => n8, A => n69, ZN => n190);
   U105 : NAND2_X1 port map( A1 => N161, A2 => n14, ZN => n70);
   U106 : OAI21_X1 port map( B1 => n107, B2 => n8, A => n70, ZN => n191);
   U107 : NAND2_X1 port map( A1 => N160, A2 => n15, ZN => n71);
   U108 : OAI21_X1 port map( B1 => n106, B2 => n8, A => n71, ZN => n192);
   U109 : NAND2_X1 port map( A1 => N159, A2 => n15, ZN => n72);
   U110 : OAI21_X1 port map( B1 => n105, B2 => n8, A => n72, ZN => n193);
   U111 : NAND2_X1 port map( A1 => N158, A2 => n15, ZN => n73);
   U112 : OAI21_X1 port map( B1 => n104, B2 => n8, A => n73, ZN => n194);
   U113 : NAND2_X1 port map( A1 => N157, A2 => n15, ZN => n74);
   U114 : OAI21_X1 port map( B1 => n103, B2 => n8, A => n74, ZN => n195);
   U115 : NAND2_X1 port map( A1 => N156, A2 => n15, ZN => n75);
   U116 : OAI21_X1 port map( B1 => n102, B2 => n8, A => n75, ZN => n196);
   U117 : MUX2_X1 port map( A => N154, B => cnt_mul_1_port, S => n12, Z => n79)
                           ;
   U118 : INV_X1 port map( A => n76, ZN => n77);
   U119 : NAND2_X1 port map( A1 => n77, A2 => n8, ZN => n81);
   U120 : INV_X1 port map( A => n81, ZN => n78);
   U121 : OR2_X1 port map( A1 => n79, A2 => n78, ZN => n200);
   U122 : NAND2_X1 port map( A1 => n81, A2 => n80, ZN => n202);
   U123 : NAND2_X1 port map( A1 => N155, A2 => n15, ZN => n82);
   U124 : OAI21_X1 port map( B1 => n101, B2 => n9, A => n82, ZN => n197);
   U125 : MUX2_X1 port map( A => n146, B => IR(31), S => n199, Z => n159_port);
   U126 : MUX2_X1 port map( A => n136, B => IR(16), S => n199, Z => n149);
   U127 : MUX2_X1 port map( A => n137, B => IR(17), S => n199, Z => n150);
   U128 : MUX2_X1 port map( A => n140, B => IR(20), S => n199, Z => n153);
   U129 : MUX2_X1 port map( A => n138, B => IR(18), S => n199, Z => n151);
   U130 : MUX2_X1 port map( A => n139, B => IR(19), S => n199, Z => n152);
   U131 : MUX2_X1 port map( A => n144, B => IR(27), S => n199, Z => n155_port);
   U132 : MUX2_X1 port map( A => n141, B => IR(26), S => n199, Z => n154_port);
   U133 : MUX2_X1 port map( A => n145, B => IR(28), S => n199, Z => n156_port);
   U134 : MUX2_X1 port map( A => n143, B => IR(29), S => n199, Z => n157_port);
   U135 : MUX2_X1 port map( A => n142, B => IR(30), S => n199, Z => n158_port);
   U136 : INV_X1 port map( A => IR(26), ZN => n83);
   U137 : INV_X1 port map( A => IR(28), ZN => n86);
   U138 : NAND2_X1 port map( A1 => n83, A2 => n86, ZN => n118);
   U139 : MUX2_X1 port map( A => n87, B => n86, S => IR(27), Z => n89);
   U140 : NAND3_X1 port map( A1 => n90, A2 => n89, A3 => n88, ZN => n97);
   U141 : NAND3_X1 port map( A1 => n93, A2 => n92, A3 => n91, ZN => n94);
   U142 : NAND3_X1 port map( A1 => n97, A2 => n96, A3 => n95, ZN => n131);
   U143 : NAND3_X1 port map( A1 => n124, A2 => n123, A3 => n122, ZN => n130);
   U144 : NAND2_X1 port map( A1 => n199, A2 => n135, ZN => IF_STALL_port);
   U145 : INV_X1 port map( A => n135, ZN => STALL_CODE_0_port);
   U146 : NOR2_X1 port map( A1 => n199, A2 => STALL_CODE_0_port, ZN => 
                           STALL_CODE_1_port);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWDU_IR_SIZE32 is

   port( CLOCK, RESET, EN : in std_logic;  IR : in std_logic_vector (31 downto 
         0);  FWD_A, FWD_B : out std_logic_vector (1 downto 0);  FWD_B2 : out 
         std_logic;  ZDU_SEL : out std_logic_vector (1 downto 0));

end FWDU_IR_SIZE32;

architecture SYN_BEHAVIORAL of FWDU_IR_SIZE32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal FWD_B2_port, n106, n107, n108, n109, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n175, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n174, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733 : std_logic;

begin
   FWD_B2 <= FWD_B2_port;
   
   IR_EX_reg_31_inst : DFFR_X1 port map( D => n175, CK => CLOCK, RN => n15, Q 
                           => n185, QN => n1);
   IR_EX_reg_30_inst : DFFR_X1 port map( D => n173, CK => CLOCK, RN => n15, Q 
                           => n187, QN => n3);
   IR_EX_reg_28_inst : DFFR_X1 port map( D => n171, CK => CLOCK, RN => n15, Q 
                           => n135, QN => n4);
   IR_EX_reg_27_inst : DFFR_X1 port map( D => n170, CK => CLOCK, RN => n15, Q 
                           => n134, QN => n2);
   FWD_B2_tmp2_reg : DFF_X1 port map( D => n143, CK => CLOCK, Q => n132, QN => 
                           n_1727);
   FWD_B2_reg : DFF_X1 port map( D => n142, CK => CLOCK, Q => FWD_B2_port, QN 
                           => n_1728);
   FWD_A_reg_1_inst : DFF_X1 port map( D => n141, CK => CLOCK, Q => FWD_A(1), 
                           QN => n109);
   FWD_A_reg_0_inst : DFF_X1 port map( D => n140, CK => CLOCK, Q => FWD_A(0), 
                           QN => n108);
   FWD_B_reg_1_inst : DFF_X1 port map( D => n139, CK => CLOCK, Q => FWD_B(1), 
                           QN => n107);
   FWD_B_reg_0_inst : DFF_X1 port map( D => n138, CK => CLOCK, Q => FWD_B(0), 
                           QN => n106);
   ZDU_SEL_reg_1_inst : DFF_X1 port map( D => n137, CK => CLOCK, Q => 
                           ZDU_SEL(1), QN => n61);
   ZDU_SEL_reg_0_inst : DFF_X1 port map( D => n136, CK => CLOCK, Q => 
                           ZDU_SEL(0), QN => n47);
   IR_EX_reg_12_inst : DFFR_X1 port map( D => n160, CK => CLOCK, RN => n17, Q 
                           => n177, QN => n_1729);
   IR_EX_reg_18_inst : DFFR_X1 port map( D => n166, CK => CLOCK, RN => n17, Q 
                           => n180, QN => n28);
   IR_MEM_reg_31_inst : DFFR_X1 port map( D => n158, CK => CLOCK, RN => n17, Q 
                           => n198, QN => n80);
   IR_MEM_reg_30_inst : DFFR_X1 port map( D => n157, CK => CLOCK, RN => n17, Q 
                           => n201, QN => n_1730);
   IR_MEM_reg_29_inst : DFFR_X1 port map( D => n156, CK => CLOCK, RN => n17, Q 
                           => n202, QN => n81);
   IR_MEM_reg_28_inst : DFFR_X1 port map( D => n155, CK => CLOCK, RN => n17, Q 
                           => n199, QN => n38);
   IR_MEM_reg_27_inst : DFFR_X1 port map( D => n154, CK => CLOCK, RN => n17, Q 
                           => n200, QN => n_1731);
   IR_MEM_reg_20_inst : DFFR_X1 port map( D => n153, CK => CLOCK, RN => n17, Q 
                           => n197, QN => n40);
   IR_MEM_reg_19_inst : DFFR_X1 port map( D => n152, CK => CLOCK, RN => n17, Q 
                           => n195, QN => n44);
   IR_MEM_reg_18_inst : DFFR_X1 port map( D => n151, CK => CLOCK, RN => n17, Q 
                           => n193, QN => n59);
   IR_MEM_reg_17_inst : DFFR_X1 port map( D => n150, CK => CLOCK, RN => n17, Q 
                           => n191, QN => n50);
   IR_MEM_reg_16_inst : DFFR_X1 port map( D => n149, CK => CLOCK, RN => n17, Q 
                           => n189, QN => n52);
   IR_MEM_reg_15_inst : DFFR_X1 port map( D => n148, CK => CLOCK, RN => n17, Q 
                           => n196, QN => n39);
   IR_MEM_reg_14_inst : DFFR_X1 port map( D => n147, CK => CLOCK, RN => n17, Q 
                           => n194, QN => n43);
   IR_MEM_reg_13_inst : DFFR_X1 port map( D => n146, CK => CLOCK, RN => n17, Q 
                           => n192, QN => n58);
   IR_MEM_reg_12_inst : DFFR_X1 port map( D => n145, CK => CLOCK, RN => n17, Q 
                           => n190, QN => n49);
   IR_MEM_reg_11_inst : DFFR_X1 port map( D => n144, CK => CLOCK, RN => n17, Q 
                           => n188, QN => n51);
   IR_EX_reg_26_inst : DFFR_X1 port map( D => n169, CK => CLOCK, RN => n17, Q 
                           => n133, QN => n_1732);
   IR_EX_reg_14_inst : DFFR_X1 port map( D => n162, CK => CLOCK, RN => n17, Q 
                           => n181, QN => n23);
   IR_EX_reg_13_inst : DFFR_X1 port map( D => n161, CK => CLOCK, RN => n17, Q 
                           => n179, QN => n27);
   IR_EX_reg_11_inst : DFFR_X1 port map( D => n159, CK => CLOCK, RN => n17, Q 
                           => n174, QN => n25);
   IR_EX_reg_17_inst : DFFR_X1 port map( D => n165, CK => CLOCK, RN => n17, Q 
                           => n178, QN => n_1733);
   IR_EX_reg_19_inst : DFFR_X1 port map( D => n167, CK => CLOCK, RN => n17, Q 
                           => n182, QN => n24);
   IR_EX_reg_20_inst : DFFR_X1 port map( D => n168, CK => CLOCK, RN => n17, Q 
                           => n184, QN => n22);
   IR_EX_reg_16_inst : DFFR_X1 port map( D => n164, CK => CLOCK, RN => n17, Q 
                           => n176, QN => n26);
   IR_EX_reg_15_inst : DFFR_X1 port map( D => n163, CK => CLOCK, RN => n17, Q 
                           => n183, QN => n21);
   IR_EX_reg_29_inst : DFFR_X1 port map( D => n172, CK => CLOCK, RN => n17, Q 
                           => n186, QN => n89);
   U2 : INV_X2 port map( A => RESET, ZN => n17);
   U3 : BUF_X1 port map( A => EN, Z => n14);
   U4 : BUF_X1 port map( A => n17, Z => n16);
   U5 : AND2_X1 port map( A1 => n13, A2 => n16, ZN => n5);
   U6 : BUF_X1 port map( A => n14, Z => n13);
   U7 : BUF_X1 port map( A => n14, Z => n12);
   U8 : BUF_X1 port map( A => n14, Z => n11);
   U9 : BUF_X1 port map( A => n16, Z => n15);
   U10 : INV_X1 port map( A => n48, ZN => n57);
   U11 : OR2_X1 port map( A1 => n93, A2 => n94, ZN => n117);
   U12 : OAI22_X1 port map( A1 => n63, A2 => n62, B1 => n5, B2 => n61, ZN => 
                           n137);
   U13 : NAND2_X1 port map( A1 => n123, A2 => n60, ZN => n62);
   U14 : NAND4_X1 port map( A1 => n87, A2 => n57, A3 => n85, A4 => n10, ZN => 
                           n63);
   U15 : AND3_X1 port map( A1 => n3, A2 => n1, A3 => n20, ZN => n6);
   U16 : XNOR2_X1 port map( A => IR(20), B => n69, ZN => n71);
   U17 : MUX2_X1 port map( A => n178, B => n177, S => n6, Z => n7);
   U18 : XNOR2_X1 port map( A => IR(19), B => n68, ZN => n72);
   U19 : XNOR2_X1 port map( A => IR(23), B => n67, ZN => n29);
   U20 : AND4_X1 port map( A1 => n9, A2 => n81, A3 => n80, A4 => n38, ZN => n8)
                           ;
   U21 : NOR2_X1 port map( A1 => n200, A2 => n201, ZN => n9);
   U22 : XNOR2_X1 port map( A => IR(21), B => n66, ZN => n31);
   U23 : AND4_X1 port map( A1 => n56, A2 => n55, A3 => n54, A4 => n53, ZN => 
                           n10);
   U24 : MUX2_X1 port map( A => n179, B => IR(13), S => n11, Z => n161);
   U25 : MUX2_X1 port map( A => n180, B => IR(18), S => n13, Z => n166);
   U26 : MUX2_X1 port map( A => n134, B => IR(27), S => n13, Z => n170);
   U27 : MUX2_X1 port map( A => n135, B => IR(28), S => n13, Z => n171);
   U28 : MUX2_X1 port map( A => n186, B => IR(29), S => n13, Z => n172);
   U29 : MUX2_X1 port map( A => n187, B => IR(30), S => n13, Z => n173);
   U30 : MUX2_X1 port map( A => n185, B => IR(31), S => n13, Z => n175);
   U31 : MUX2_X1 port map( A => n177, B => IR(12), S => n13, Z => n160);
   U32 : MUX2_X1 port map( A => n178, B => IR(17), S => n12, Z => n165);
   U33 : MUX2_X1 port map( A => n174, B => IR(11), S => n12, Z => n159);
   U34 : MUX2_X1 port map( A => n176, B => IR(16), S => n12, Z => n164);
   U35 : MUX2_X1 port map( A => n183, B => IR(15), S => n12, Z => n163);
   U36 : MUX2_X1 port map( A => n184, B => IR(20), S => n12, Z => n168);
   U37 : MUX2_X1 port map( A => n181, B => IR(14), S => n12, Z => n162);
   U38 : MUX2_X1 port map( A => n182, B => IR(19), S => n12, Z => n167);
   U39 : MUX2_X1 port map( A => n188, B => n174, S => n12, Z => n144);
   U40 : MUX2_X1 port map( A => n190, B => n177, S => n12, Z => n145);
   U41 : MUX2_X1 port map( A => n192, B => n179, S => n12, Z => n146);
   U42 : MUX2_X1 port map( A => n189, B => n176, S => n12, Z => n149);
   U43 : MUX2_X1 port map( A => n191, B => n178, S => n11, Z => n150);
   U44 : MUX2_X1 port map( A => n193, B => n180, S => n11, Z => n151);
   U45 : MUX2_X1 port map( A => n200, B => n134, S => n11, Z => n154);
   U46 : MUX2_X1 port map( A => n201, B => n187, S => n11, Z => n157);
   U47 : MUX2_X1 port map( A => n202, B => n186, S => n11, Z => n156);
   U48 : MUX2_X1 port map( A => n198, B => n185, S => n11, Z => n158);
   U49 : MUX2_X1 port map( A => n199, B => n135, S => n11, Z => n155);
   U50 : MUX2_X1 port map( A => n196, B => n183, S => n11, Z => n148);
   U51 : MUX2_X1 port map( A => n197, B => n184, S => n11, Z => n153);
   U52 : MUX2_X1 port map( A => n194, B => n181, S => n11, Z => n147);
   U53 : MUX2_X1 port map( A => n195, B => n182, S => n11, Z => n152);
   U54 : INV_X1 port map( A => IR(30), ZN => n64);
   U55 : INV_X1 port map( A => IR(31), ZN => n19);
   U56 : INV_X1 port map( A => IR(29), ZN => n18);
   U57 : INV_X1 port map( A => IR(27), ZN => n65);
   U58 : NAND4_X1 port map( A1 => n64, A2 => n19, A3 => n18, A4 => n65, ZN => 
                           n90);
   U59 : INV_X1 port map( A => n90, ZN => n120);
   U60 : NAND3_X1 port map( A1 => IR(28), A2 => n5, A3 => n120, ZN => n48);
   U61 : NOR3_X1 port map( A1 => n186, A2 => n135, A3 => n134, ZN => n20);
   U62 : MUX2_X1 port map( A => n22, B => n21, S => n6, Z => n69);
   U63 : XOR2_X1 port map( A => n69, B => IR(25), Z => n34);
   U64 : MUX2_X1 port map( A => n24, B => n23, S => n6, Z => n68);
   U65 : XOR2_X1 port map( A => n68, B => IR(24), Z => n33);
   U66 : MUX2_X1 port map( A => n26, B => n25, S => n6, Z => n66);
   U67 : XOR2_X1 port map( A => IR(22), B => n7, Z => n30);
   U68 : MUX2_X1 port map( A => n28, B => n27, S => n6, Z => n67);
   U69 : NOR3_X1 port map( A1 => n31, A2 => n30, A3 => n29, ZN => n32);
   U70 : NAND3_X1 port map( A1 => n34, A2 => n33, A3 => n32, ZN => n60);
   U71 : INV_X1 port map( A => n60, ZN => n126);
   U72 : NOR3_X1 port map( A1 => n180, A2 => n176, A3 => n178, ZN => n36);
   U73 : NOR3_X1 port map( A1 => n179, A2 => n174, A3 => n177, ZN => n35);
   U74 : MUX2_X1 port map( A => n36, B => n35, S => n6, Z => n37);
   U75 : NAND3_X1 port map( A1 => n68, A2 => n37, A3 => n69, ZN => n85);
   U76 : MUX2_X1 port map( A => n40, B => n39, S => n8, Z => n99);
   U77 : NOR3_X1 port map( A1 => n193, A2 => n191, A3 => n189, ZN => n42);
   U78 : NOR3_X1 port map( A1 => n192, A2 => n190, A3 => n188, ZN => n41);
   U79 : MUX2_X1 port map( A => n42, B => n41, S => n8, Z => n45);
   U80 : MUX2_X1 port map( A => n44, B => n43, S => n8, Z => n96);
   U81 : NAND3_X1 port map( A1 => n99, A2 => n45, A3 => n96, ZN => n87);
   U82 : NAND4_X1 port map( A1 => n57, A2 => n126, A3 => n85, A4 => n87, ZN => 
                           n46);
   U83 : OAI21_X1 port map( B1 => n5, B2 => n47, A => n46, ZN => n136);
   U84 : MUX2_X1 port map( A => n50, B => n49, S => n8, Z => n95);
   U85 : XOR2_X1 port map( A => n95, B => IR(22), Z => n56);
   U86 : MUX2_X1 port map( A => n52, B => n51, S => n8, Z => n97);
   U87 : XOR2_X1 port map( A => n97, B => IR(21), Z => n55);
   U88 : XOR2_X1 port map( A => n99, B => IR(25), Z => n54);
   U89 : XOR2_X1 port map( A => n96, B => IR(24), Z => n53);
   U90 : MUX2_X1 port map( A => n59, B => n58, S => n8, Z => n101);
   U91 : XOR2_X1 port map( A => n101, B => IR(23), Z => n123);
   U92 : INV_X1 port map( A => IR(28), ZN => n119);
   U93 : OAI211_X1 port map( C1 => IR(26), C2 => n65, A => n119, B => n64, ZN 
                           => n78);
   U94 : NAND2_X1 port map( A1 => IR(29), A2 => IR(31), ZN => n77);
   U95 : NOR4_X1 port map( A1 => n131, A2 => IR(18), A3 => IR(19), A4 => IR(20)
                           , ZN => n76);
   U96 : XOR2_X1 port map( A => n66, B => IR(16), Z => n75);
   U97 : XOR2_X1 port map( A => n67, B => IR(18), Z => n74);
   U98 : XOR2_X1 port map( A => IR(17), B => n7, Z => n70);
   U99 : NOR3_X1 port map( A1 => n72, A2 => n71, A3 => n70, ZN => n73);
   U100 : NAND3_X1 port map( A1 => n75, A2 => n74, A3 => n73, ZN => n94);
   U101 : NOR4_X1 port map( A1 => n78, A2 => n77, A3 => n76, A4 => n94, ZN => 
                           n79);
   U102 : MUX2_X1 port map( A => n132, B => n79, S => n5, Z => n143);
   U103 : MUX2_X1 port map( A => FWD_B2_port, B => n132, S => n5, Z => n142);
   U104 : MUX2_X1 port map( A => n133, B => IR(26), S => n12, Z => n169);
   U105 : MUX2_X1 port map( A => n200, B => n9, S => n199, Z => n82);
   U106 : NAND3_X1 port map( A1 => n82, A2 => n81, A3 => n80, ZN => n128);
   U107 : INV_X1 port map( A => n128, ZN => n115);
   U108 : NOR2_X1 port map( A1 => n187, A2 => n134, ZN => n83);
   U109 : MUX2_X1 port map( A => n134, B => n83, S => n135, Z => n84);
   U110 : NAND3_X1 port map( A1 => n84, A2 => n89, A3 => n1, ZN => n125);
   U111 : INV_X1 port map( A => n125, ZN => n86);
   U112 : OAI221_X1 port map( B1 => n115, B2 => n87, C1 => n86, C2 => n85, A =>
                           n5, ZN => n92);
   U113 : MUX2_X1 port map( A => n2, B => n4, S => n133, Z => n88);
   U114 : NAND4_X1 port map( A1 => n185, A2 => n89, A3 => n88, A4 => n3, ZN => 
                           n93);
   U115 : NOR3_X1 port map( A1 => IR(28), A2 => n90, A3 => n94, ZN => n91);
   U116 : OAI211_X1 port map( C1 => IR(26), C2 => n93, A => n125, B => n91, ZN 
                           => n113);
   U117 : OAI22_X1 port map( A1 => n92, A2 => n113, B1 => n106, B2 => n5, ZN =>
                           n138);
   U118 : INV_X1 port map( A => n92, ZN => n129);
   U119 : XOR2_X1 port map( A => n95, B => IR(17), Z => n112);
   U120 : XOR2_X1 port map( A => n96, B => IR(19), Z => n111);
   U121 : INV_X1 port map( A => n97, ZN => n98);
   U122 : XOR2_X1 port map( A => IR(16), B => n98, Z => n105);
   U123 : INV_X1 port map( A => n99, ZN => n100);
   U124 : XOR2_X1 port map( A => IR(20), B => n100, Z => n104);
   U125 : INV_X1 port map( A => n101, ZN => n102);
   U126 : XOR2_X1 port map( A => IR(18), B => n102, Z => n103);
   U127 : NOR3_X1 port map( A1 => n105, A2 => n104, A3 => n103, ZN => n110);
   U128 : NAND3_X1 port map( A1 => n112, A2 => n111, A3 => n110, ZN => n116);
   U129 : INV_X1 port map( A => n113, ZN => n114);
   U130 : AOI211_X1 port map( C1 => n117, C2 => n116, A => n115, B => n114, ZN 
                           => n118);
   U131 : NAND4_X1 port map( A1 => n120, A2 => n129, A3 => n119, A4 => n118, ZN
                           => n121);
   U132 : OAI21_X1 port map( B1 => n107, B2 => n5, A => n121, ZN => n139);
   U133 : NAND3_X1 port map( A1 => n126, A2 => n129, A3 => n125, ZN => n122);
   U134 : OAI21_X1 port map( B1 => n108, B2 => n5, A => n122, ZN => n140);
   U135 : INV_X1 port map( A => n123, ZN => n124);
   U136 : AOI21_X1 port map( B1 => n126, B2 => n125, A => n124, ZN => n127);
   U137 : NAND4_X1 port map( A1 => n129, A2 => n128, A3 => n127, A4 => n10, ZN 
                           => n130);
   U138 : OAI21_X1 port map( B1 => n109, B2 => n5, A => n130, ZN => n141);
   U139 : OR2_X1 port map( A1 => IR(17), A2 => IR(16), ZN => n131);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( CLOCK : in std_logic;  AluOpcode : in std_logic_vector (0 to 4);  A, B
         : in std_logic_vector (31 downto 0);  Cin : in std_logic;  ALU_out : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic;  COND : out
         std_logic_vector (5 downto 0));

end ALU_NBIT32;

architecture SYN_BEHAVIORAL of ALU_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX4to1_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUL
      port( CLOCK : in std_logic;  A, B : in std_logic_vector (15 downto 0);  Y
            : out std_logic_vector (31 downto 0));
   end component;
   
   component CMP_NBIT32
      port( SUM : in std_logic_vector (31 downto 0);  Cout : in std_logic;  
            A_L_B, A_LE_B, A_G_B, A_GE_B, A_E_B, A_NE_B : out std_logic);
   end component;
   
   component LOGIC_NBIT32_N_SELECTOR4
      port( S : in std_logic_vector (3 downto 0);  A, B : in std_logic_vector 
            (31 downto 0);  O : out std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER
      port( data_in : in std_logic_vector (31 downto 0);  R : in 
            std_logic_vector (4 downto 0);  conf : in std_logic_vector (1 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component AND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal Cout_port, cin_internal, en_adder, A_adder_31_port, A_adder_30_port, 
      A_adder_29_port, A_adder_28_port, A_adder_27_port, A_adder_26_port, 
      A_adder_25_port, A_adder_24_port, A_adder_23_port, A_adder_22_port, 
      A_adder_21_port, A_adder_20_port, A_adder_19_port, A_adder_18_port, 
      A_adder_17_port, A_adder_16_port, A_adder_15_port, A_adder_14_port, 
      A_adder_13_port, A_adder_12_port, A_adder_11_port, A_adder_10_port, 
      A_adder_9_port, A_adder_8_port, A_adder_7_port, A_adder_6_port, 
      A_adder_5_port, A_adder_4_port, A_adder_3_port, A_adder_2_port, 
      A_adder_1_port, A_adder_0_port, B_adder_31_port, B_adder_30_port, 
      B_adder_29_port, B_adder_28_port, B_adder_27_port, B_adder_26_port, 
      B_adder_25_port, B_adder_24_port, B_adder_23_port, B_adder_22_port, 
      B_adder_21_port, B_adder_20_port, B_adder_19_port, B_adder_18_port, 
      B_adder_17_port, B_adder_16_port, B_adder_15_port, B_adder_14_port, 
      B_adder_13_port, B_adder_12_port, B_adder_11_port, B_adder_10_port, 
      B_adder_9_port, B_adder_8_port, B_adder_7_port, B_adder_6_port, 
      B_adder_5_port, B_adder_4_port, B_adder_3_port, B_adder_2_port, 
      B_adder_1_port, B_adder_0_port, A_logic_31_port, A_logic_30_port, 
      A_logic_29_port, A_logic_28_port, A_logic_27_port, A_logic_26_port, 
      A_logic_25_port, A_logic_24_port, A_logic_23_port, A_logic_22_port, 
      A_logic_21_port, A_logic_20_port, A_logic_19_port, A_logic_18_port, 
      A_logic_17_port, A_logic_16_port, A_logic_15_port, A_logic_14_port, 
      A_logic_13_port, A_logic_12_port, A_logic_11_port, A_logic_10_port, 
      A_logic_9_port, A_logic_8_port, A_logic_7_port, A_logic_6_port, 
      A_logic_5_port, A_logic_4_port, A_logic_3_port, A_logic_2_port, 
      A_logic_1_port, A_logic_0_port, B_logic_31_port, B_logic_30_port, 
      B_logic_29_port, B_logic_28_port, B_logic_27_port, B_logic_26_port, 
      B_logic_25_port, B_logic_24_port, B_logic_23_port, B_logic_22_port, 
      B_logic_21_port, B_logic_20_port, B_logic_19_port, B_logic_18_port, 
      B_logic_17_port, B_logic_16_port, B_logic_15_port, B_logic_14_port, 
      B_logic_13_port, B_logic_12_port, B_logic_11_port, B_logic_10_port, 
      B_logic_9_port, B_logic_8_port, B_logic_7_port, B_logic_6_port, 
      B_logic_5_port, B_logic_4_port, B_logic_3_port, B_logic_2_port, 
      B_logic_1_port, B_logic_0_port, A_shifter_31_port, A_shifter_30_port, 
      A_shifter_29_port, A_shifter_28_port, A_shifter_27_port, 
      A_shifter_26_port, A_shifter_25_port, A_shifter_24_port, 
      A_shifter_23_port, A_shifter_22_port, A_shifter_21_port, 
      A_shifter_20_port, A_shifter_19_port, A_shifter_18_port, 
      A_shifter_17_port, A_shifter_16_port, A_shifter_15_port, 
      A_shifter_14_port, A_shifter_13_port, A_shifter_12_port, 
      A_shifter_11_port, A_shifter_10_port, A_shifter_9_port, A_shifter_8_port,
      A_shifter_7_port, A_shifter_6_port, A_shifter_5_port, A_shifter_4_port, 
      A_shifter_3_port, A_shifter_2_port, A_shifter_1_port, A_shifter_0_port, 
      B_shifter_4_port, B_shifter_3_port, B_shifter_2_port, B_shifter_1_port, 
      B_shifter_0_port, in_cmp_31_port, in_cmp_30_port, in_cmp_29_port, 
      in_cmp_28_port, in_cmp_27_port, in_cmp_26_port, in_cmp_25_port, 
      in_cmp_24_port, in_cmp_23_port, in_cmp_22_port, in_cmp_21_port, 
      in_cmp_20_port, in_cmp_19_port, in_cmp_18_port, in_cmp_17_port, 
      in_cmp_16_port, in_cmp_15_port, in_cmp_14_port, in_cmp_13_port, 
      in_cmp_12_port, in_cmp_11_port, in_cmp_10_port, in_cmp_9_port, 
      in_cmp_8_port, in_cmp_7_port, in_cmp_6_port, in_cmp_5_port, in_cmp_4_port
      , in_cmp_3_port, in_cmp_2_port, in_cmp_1_port, in_cmp_0_port, 
      out_adder_31_port, out_adder_30_port, out_adder_29_port, 
      out_adder_28_port, out_adder_27_port, out_adder_26_port, 
      out_adder_25_port, out_adder_24_port, out_adder_23_port, 
      out_adder_22_port, out_adder_21_port, out_adder_20_port, 
      out_adder_19_port, out_adder_18_port, out_adder_17_port, 
      out_adder_16_port, out_adder_15_port, out_adder_14_port, 
      out_adder_13_port, out_adder_12_port, out_adder_11_port, 
      out_adder_10_port, out_adder_9_port, out_adder_8_port, out_adder_7_port, 
      out_adder_6_port, out_adder_5_port, out_adder_4_port, out_adder_3_port, 
      out_adder_2_port, out_adder_1_port, out_adder_0_port, A_mul_15_port, 
      A_mul_14_port, A_mul_13_port, A_mul_12_port, A_mul_11_port, A_mul_10_port
      , A_mul_9_port, A_mul_8_port, A_mul_7_port, A_mul_6_port, A_mul_5_port, 
      A_mul_4_port, A_mul_3_port, A_mul_2_port, A_mul_1_port, A_mul_0_port, 
      B_mul_15_port, B_mul_14_port, B_mul_13_port, B_mul_12_port, B_mul_11_port
      , B_mul_10_port, B_mul_9_port, B_mul_8_port, B_mul_7_port, B_mul_6_port, 
      B_mul_5_port, B_mul_4_port, B_mul_3_port, B_mul_2_port, B_mul_1_port, 
      B_mul_0_port, conf_1_port, conf_0_port, out_shifter_31_port, 
      out_shifter_30_port, out_shifter_29_port, out_shifter_28_port, 
      out_shifter_27_port, out_shifter_26_port, out_shifter_25_port, 
      out_shifter_24_port, out_shifter_23_port, out_shifter_22_port, 
      out_shifter_21_port, out_shifter_20_port, out_shifter_19_port, 
      out_shifter_18_port, out_shifter_17_port, out_shifter_16_port, 
      out_shifter_15_port, out_shifter_14_port, out_shifter_13_port, 
      out_shifter_12_port, out_shifter_11_port, out_shifter_10_port, 
      out_shifter_9_port, out_shifter_8_port, out_shifter_7_port, 
      out_shifter_6_port, out_shifter_5_port, out_shifter_4_port, 
      out_shifter_3_port, out_shifter_2_port, out_shifter_1_port, 
      out_shifter_0_port, logic_sel_3_port, logic_sel_2_port, logic_sel_1_port,
      logic_sel_0_port, out_logic_31_port, out_logic_30_port, out_logic_29_port
      , out_logic_28_port, out_logic_27_port, out_logic_26_port, 
      out_logic_25_port, out_logic_24_port, out_logic_23_port, 
      out_logic_22_port, out_logic_21_port, out_logic_20_port, 
      out_logic_19_port, out_logic_18_port, out_logic_17_port, 
      out_logic_16_port, out_logic_15_port, out_logic_14_port, 
      out_logic_13_port, out_logic_12_port, out_logic_11_port, 
      out_logic_10_port, out_logic_9_port, out_logic_8_port, out_logic_7_port, 
      out_logic_6_port, out_logic_5_port, out_logic_4_port, out_logic_3_port, 
      out_logic_2_port, out_logic_1_port, out_logic_0_port, out_mul_31_port, 
      out_mul_30_port, out_mul_29_port, out_mul_28_port, out_mul_27_port, 
      out_mul_26_port, out_mul_25_port, out_mul_24_port, out_mul_23_port, 
      out_mul_22_port, out_mul_21_port, out_mul_20_port, out_mul_19_port, 
      out_mul_18_port, out_mul_17_port, out_mul_16_port, out_mul_15_port, 
      out_mul_14_port, out_mul_13_port, out_mul_12_port, out_mul_11_port, 
      out_mul_10_port, out_mul_9_port, out_mul_8_port, out_mul_7_port, 
      out_mul_6_port, out_mul_5_port, out_mul_4_port, out_mul_3_port, 
      out_mul_2_port, out_mul_1_port, out_mul_0_port, mux_out_1_port, 
      mux_out_0_port, N88, N89, N90, N91, N92, N93, n21, n1, n2, n3, n4, n5, n6
      , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n22,
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70 : std_logic;

begin
   Cout <= Cout_port;
   
   conf_reg_1_inst : DLH_X1 port map( G => N91, D => N93, Q => conf_1_port);
   conf_reg_0_inst : DLH_X1 port map( G => N91, D => N92, Q => conf_0_port);
   logic_sel_reg_3_inst : DLH_X1 port map( G => n28, D => N90, Q => 
                           logic_sel_3_port);
   logic_sel_reg_2_inst : DLH_X1 port map( G => n29, D => N89, Q => 
                           logic_sel_2_port);
   logic_sel_reg_1_inst : DLH_X1 port map( G => n29, D => N89, Q => 
                           logic_sel_1_port);
   logic_sel_reg_0_inst : DLH_X1 port map( G => n28, D => N88, Q => 
                           logic_sel_0_port);
   ADDER_A_i_0 : AND2_0 port map( A => A(0), B => en_adder, Y => A_adder_0_port
                           );
   ADDER_B_i_0 : AND2_228 port map( A => B(0), B => n66, Y => B_adder_0_port);
   ADDER_A_i_1 : AND2_227 port map( A => A(1), B => n17, Y => A_adder_1_port);
   ADDER_B_i_1 : AND2_226 port map( A => B(1), B => en_adder, Y => 
                           B_adder_1_port);
   ADDER_A_i_2 : AND2_225 port map( A => A(2), B => n13, Y => A_adder_2_port);
   ADDER_B_i_2 : AND2_224 port map( A => B(2), B => n67, Y => B_adder_2_port);
   ADDER_A_i_3 : AND2_223 port map( A => A(3), B => n18, Y => A_adder_3_port);
   ADDER_B_i_3 : AND2_222 port map( A => B(3), B => n67, Y => B_adder_3_port);
   ADDER_A_i_4 : AND2_221 port map( A => A(4), B => n13, Y => A_adder_4_port);
   ADDER_B_i_4 : AND2_220 port map( A => B(4), B => n67, Y => B_adder_4_port);
   ADDER_A_i_5 : AND2_219 port map( A => A(5), B => n17, Y => A_adder_5_port);
   ADDER_B_i_5 : AND2_218 port map( A => B(5), B => en_adder, Y => 
                           B_adder_5_port);
   ADDER_A_i_6 : AND2_217 port map( A => A(6), B => n13, Y => A_adder_6_port);
   ADDER_B_i_6 : AND2_216 port map( A => B(6), B => n67, Y => B_adder_6_port);
   ADDER_A_i_7 : AND2_215 port map( A => A(7), B => n18, Y => A_adder_7_port);
   ADDER_B_i_7 : AND2_214 port map( A => B(7), B => n67, Y => B_adder_7_port);
   ADDER_A_i_8 : AND2_213 port map( A => A(8), B => n13, Y => A_adder_8_port);
   ADDER_B_i_8 : AND2_212 port map( A => B(8), B => n13, Y => B_adder_8_port);
   ADDER_A_i_9 : AND2_211 port map( A => A(9), B => n14, Y => A_adder_9_port);
   ADDER_B_i_9 : AND2_210 port map( A => B(9), B => n13, Y => B_adder_9_port);
   ADDER_A_i_10 : AND2_209 port map( A => A(10), B => n4, Y => A_adder_10_port)
                           ;
   ADDER_B_i_10 : AND2_208 port map( A => B(10), B => n13, Y => B_adder_10_port
                           );
   ADDER_A_i_11 : AND2_207 port map( A => A(11), B => n16, Y => A_adder_11_port
                           );
   ADDER_B_i_11 : AND2_206 port map( A => B(11), B => n13, Y => B_adder_11_port
                           );
   ADDER_A_i_12 : AND2_205 port map( A => A(12), B => n14, Y => A_adder_12_port
                           );
   ADDER_B_i_12 : AND2_204 port map( A => B(12), B => n17, Y => B_adder_12_port
                           );
   ADDER_A_i_13 : AND2_203 port map( A => A(13), B => n14, Y => A_adder_13_port
                           );
   ADDER_B_i_13 : AND2_202 port map( A => B(13), B => n67, Y => B_adder_13_port
                           );
   ADDER_A_i_14 : AND2_201 port map( A => A(14), B => n14, Y => A_adder_14_port
                           );
   ADDER_B_i_14 : AND2_200 port map( A => B(14), B => n18, Y => B_adder_14_port
                           );
   ADDER_A_i_15 : AND2_199 port map( A => A(15), B => n16, Y => A_adder_15_port
                           );
   ADDER_B_i_15 : AND2_198 port map( A => B(15), B => n13, Y => B_adder_15_port
                           );
   ADDER_A_i_16 : AND2_197 port map( A => A(16), B => n16, Y => A_adder_16_port
                           );
   ADDER_B_i_16 : AND2_196 port map( A => B(16), B => n66, Y => B_adder_16_port
                           );
   ADDER_A_i_17 : AND2_195 port map( A => A(17), B => n16, Y => A_adder_17_port
                           );
   ADDER_B_i_17 : AND2_194 port map( A => B(17), B => n15, Y => B_adder_17_port
                           );
   ADDER_A_i_18 : AND2_193 port map( A => A(18), B => n4, Y => A_adder_18_port)
                           ;
   ADDER_B_i_18 : AND2_192 port map( A => B(18), B => n15, Y => B_adder_18_port
                           );
   ADDER_A_i_19 : AND2_191 port map( A => A(19), B => n14, Y => A_adder_19_port
                           );
   ADDER_B_i_19 : AND2_190 port map( A => B(19), B => n15, Y => B_adder_19_port
                           );
   ADDER_A_i_20 : AND2_189 port map( A => A(20), B => n15, Y => A_adder_20_port
                           );
   ADDER_B_i_20 : AND2_188 port map( A => B(20), B => n15, Y => B_adder_20_port
                           );
   ADDER_A_i_21 : AND2_187 port map( A => A(21), B => n4, Y => A_adder_21_port)
                           ;
   ADDER_B_i_21 : AND2_186 port map( A => B(21), B => n15, Y => B_adder_21_port
                           );
   ADDER_A_i_22 : AND2_185 port map( A => A(22), B => n15, Y => A_adder_22_port
                           );
   ADDER_B_i_22 : AND2_184 port map( A => B(22), B => n4, Y => B_adder_22_port)
                           ;
   ADDER_A_i_23 : AND2_183 port map( A => A(23), B => n15, Y => A_adder_23_port
                           );
   ADDER_B_i_23 : AND2_182 port map( A => B(23), B => n14, Y => B_adder_23_port
                           );
   ADDER_A_i_24 : AND2_181 port map( A => A(24), B => n14, Y => A_adder_24_port
                           );
   ADDER_B_i_24 : AND2_180 port map( A => B(24), B => n15, Y => B_adder_24_port
                           );
   ADDER_A_i_25 : AND2_179 port map( A => A(25), B => n15, Y => A_adder_25_port
                           );
   ADDER_B_i_25 : AND2_178 port map( A => B(25), B => n15, Y => B_adder_25_port
                           );
   ADDER_A_i_26 : AND2_177 port map( A => A(26), B => n15, Y => A_adder_26_port
                           );
   ADDER_B_i_26 : AND2_176 port map( A => B(26), B => n16, Y => B_adder_26_port
                           );
   ADDER_A_i_27 : AND2_175 port map( A => A(27), B => n14, Y => A_adder_27_port
                           );
   ADDER_B_i_27 : AND2_174 port map( A => B(27), B => n14, Y => B_adder_27_port
                           );
   ADDER_A_i_28 : AND2_173 port map( A => A(28), B => n14, Y => A_adder_28_port
                           );
   ADDER_B_i_28 : AND2_172 port map( A => B(28), B => n14, Y => B_adder_28_port
                           );
   ADDER_A_i_29 : AND2_171 port map( A => A(29), B => n14, Y => A_adder_29_port
                           );
   ADDER_B_i_29 : AND2_170 port map( A => B(29), B => n4, Y => B_adder_29_port)
                           ;
   ADDER_A_i_30 : AND2_169 port map( A => A(30), B => n4, Y => A_adder_30_port)
                           ;
   ADDER_B_i_30 : AND2_168 port map( A => B(30), B => n15, Y => B_adder_30_port
                           );
   ADDER_A_i_31 : AND2_167 port map( A => A(31), B => n15, Y => A_adder_31_port
                           );
   ADDER_B_i_31 : AND2_166 port map( A => B(31), B => n16, Y => B_adder_31_port
                           );
   LOGIC_A_i_0 : AND2_165 port map( A => A(0), B => n28, Y => A_logic_0_port);
   LOGIC_B_i_0 : AND2_164 port map( A => B(0), B => n28, Y => B_logic_0_port);
   LOGIC_A_i_1 : AND2_163 port map( A => A(1), B => n28, Y => A_logic_1_port);
   LOGIC_B_i_1 : AND2_162 port map( A => B(1), B => n28, Y => B_logic_1_port);
   LOGIC_A_i_2 : AND2_161 port map( A => A(2), B => n28, Y => A_logic_2_port);
   LOGIC_B_i_2 : AND2_160 port map( A => B(2), B => n28, Y => B_logic_2_port);
   LOGIC_A_i_3 : AND2_159 port map( A => A(3), B => n28, Y => A_logic_3_port);
   LOGIC_B_i_3 : AND2_158 port map( A => B(3), B => n28, Y => B_logic_3_port);
   LOGIC_A_i_4 : AND2_157 port map( A => A(4), B => n28, Y => A_logic_4_port);
   LOGIC_B_i_4 : AND2_156 port map( A => B(4), B => n28, Y => B_logic_4_port);
   LOGIC_A_i_5 : AND2_155 port map( A => A(5), B => n28, Y => A_logic_5_port);
   LOGIC_B_i_5 : AND2_154 port map( A => B(5), B => n29, Y => B_logic_5_port);
   LOGIC_A_i_6 : AND2_153 port map( A => A(6), B => n29, Y => A_logic_6_port);
   LOGIC_B_i_6 : AND2_152 port map( A => B(6), B => n29, Y => B_logic_6_port);
   LOGIC_A_i_7 : AND2_151 port map( A => A(7), B => n29, Y => A_logic_7_port);
   LOGIC_B_i_7 : AND2_150 port map( A => B(7), B => n29, Y => B_logic_7_port);
   LOGIC_A_i_8 : AND2_149 port map( A => A(8), B => n29, Y => A_logic_8_port);
   LOGIC_B_i_8 : AND2_148 port map( A => B(8), B => n29, Y => B_logic_8_port);
   LOGIC_A_i_9 : AND2_147 port map( A => A(9), B => n29, Y => A_logic_9_port);
   LOGIC_B_i_9 : AND2_146 port map( A => B(9), B => n29, Y => B_logic_9_port);
   LOGIC_A_i_10 : AND2_145 port map( A => A(10), B => n29, Y => A_logic_10_port
                           );
   LOGIC_B_i_10 : AND2_144 port map( A => B(10), B => n29, Y => B_logic_10_port
                           );
   LOGIC_A_i_11 : AND2_143 port map( A => A(11), B => n29, Y => A_logic_11_port
                           );
   LOGIC_B_i_11 : AND2_142 port map( A => B(11), B => n28, Y => B_logic_11_port
                           );
   LOGIC_A_i_12 : AND2_141 port map( A => A(12), B => n29, Y => A_logic_12_port
                           );
   LOGIC_B_i_12 : AND2_140 port map( A => B(12), B => n28, Y => B_logic_12_port
                           );
   LOGIC_A_i_13 : AND2_139 port map( A => A(13), B => n29, Y => A_logic_13_port
                           );
   LOGIC_B_i_13 : AND2_138 port map( A => B(13), B => n28, Y => B_logic_13_port
                           );
   LOGIC_A_i_14 : AND2_137 port map( A => A(14), B => n29, Y => A_logic_14_port
                           );
   LOGIC_B_i_14 : AND2_136 port map( A => B(14), B => n28, Y => B_logic_14_port
                           );
   LOGIC_A_i_15 : AND2_135 port map( A => A(15), B => n29, Y => A_logic_15_port
                           );
   LOGIC_B_i_15 : AND2_134 port map( A => B(15), B => n28, Y => B_logic_15_port
                           );
   LOGIC_A_i_16 : AND2_133 port map( A => A(16), B => n29, Y => A_logic_16_port
                           );
   LOGIC_B_i_16 : AND2_132 port map( A => B(16), B => n29, Y => B_logic_16_port
                           );
   LOGIC_A_i_17 : AND2_131 port map( A => A(17), B => n29, Y => A_logic_17_port
                           );
   LOGIC_B_i_17 : AND2_130 port map( A => B(17), B => n28, Y => B_logic_17_port
                           );
   LOGIC_A_i_18 : AND2_129 port map( A => A(18), B => n28, Y => A_logic_18_port
                           );
   LOGIC_B_i_18 : AND2_128 port map( A => B(18), B => n28, Y => B_logic_18_port
                           );
   LOGIC_A_i_19 : AND2_127 port map( A => A(19), B => n29, Y => A_logic_19_port
                           );
   LOGIC_B_i_19 : AND2_126 port map( A => B(19), B => n28, Y => B_logic_19_port
                           );
   LOGIC_A_i_20 : AND2_125 port map( A => A(20), B => n29, Y => A_logic_20_port
                           );
   LOGIC_B_i_20 : AND2_124 port map( A => B(20), B => n29, Y => B_logic_20_port
                           );
   LOGIC_A_i_21 : AND2_123 port map( A => A(21), B => n29, Y => A_logic_21_port
                           );
   LOGIC_B_i_21 : AND2_122 port map( A => B(21), B => n28, Y => B_logic_21_port
                           );
   LOGIC_A_i_22 : AND2_121 port map( A => A(22), B => n29, Y => A_logic_22_port
                           );
   LOGIC_B_i_22 : AND2_120 port map( A => B(22), B => n28, Y => B_logic_22_port
                           );
   LOGIC_A_i_23 : AND2_119 port map( A => A(23), B => n28, Y => A_logic_23_port
                           );
   LOGIC_B_i_23 : AND2_118 port map( A => B(23), B => n29, Y => B_logic_23_port
                           );
   LOGIC_A_i_24 : AND2_117 port map( A => A(24), B => n28, Y => A_logic_24_port
                           );
   LOGIC_B_i_24 : AND2_116 port map( A => B(24), B => n29, Y => B_logic_24_port
                           );
   LOGIC_A_i_25 : AND2_115 port map( A => A(25), B => n29, Y => A_logic_25_port
                           );
   LOGIC_B_i_25 : AND2_114 port map( A => B(25), B => n28, Y => B_logic_25_port
                           );
   LOGIC_A_i_26 : AND2_113 port map( A => A(26), B => n28, Y => A_logic_26_port
                           );
   LOGIC_B_i_26 : AND2_112 port map( A => B(26), B => n29, Y => B_logic_26_port
                           );
   LOGIC_A_i_27 : AND2_111 port map( A => A(27), B => n28, Y => A_logic_27_port
                           );
   LOGIC_B_i_27 : AND2_110 port map( A => B(27), B => n29, Y => B_logic_27_port
                           );
   LOGIC_A_i_28 : AND2_109 port map( A => A(28), B => n28, Y => A_logic_28_port
                           );
   LOGIC_B_i_28 : AND2_108 port map( A => B(28), B => n29, Y => B_logic_28_port
                           );
   LOGIC_A_i_29 : AND2_107 port map( A => A(29), B => n28, Y => A_logic_29_port
                           );
   LOGIC_B_i_29 : AND2_106 port map( A => B(29), B => n28, Y => B_logic_29_port
                           );
   LOGIC_A_i_30 : AND2_105 port map( A => A(30), B => n29, Y => A_logic_30_port
                           );
   LOGIC_B_i_30 : AND2_104 port map( A => B(30), B => n28, Y => B_logic_30_port
                           );
   LOGIC_A_i_31 : AND2_103 port map( A => A(31), B => n29, Y => A_logic_31_port
                           );
   LOGIC_B_i_31 : AND2_102 port map( A => B(31), B => n28, Y => B_logic_31_port
                           );
   SHIFTER_A_i_0 : AND2_101 port map( A => A(0), B => n22, Y => 
                           A_shifter_0_port);
   SHIFTER_A_i_1 : AND2_100 port map( A => A(1), B => n22, Y => 
                           A_shifter_1_port);
   SHIFTER_A_i_2 : AND2_99 port map( A => A(2), B => n22, Y => A_shifter_2_port
                           );
   SHIFTER_A_i_3 : AND2_98 port map( A => A(3), B => n22, Y => A_shifter_3_port
                           );
   SHIFTER_A_i_4 : AND2_97 port map( A => A(4), B => n22, Y => A_shifter_4_port
                           );
   SHIFTER_A_i_5 : AND2_96 port map( A => A(5), B => n22, Y => A_shifter_5_port
                           );
   SHIFTER_A_i_6 : AND2_95 port map( A => A(6), B => n22, Y => A_shifter_6_port
                           );
   SHIFTER_A_i_7 : AND2_94 port map( A => A(7), B => n22, Y => A_shifter_7_port
                           );
   SHIFTER_A_i_8 : AND2_93 port map( A => A(8), B => n22, Y => A_shifter_8_port
                           );
   SHIFTER_A_i_9 : AND2_92 port map( A => A(9), B => n22, Y => A_shifter_9_port
                           );
   SHIFTER_A_i_10 : AND2_91 port map( A => A(10), B => n22, Y => 
                           A_shifter_10_port);
   SHIFTER_A_i_11 : AND2_90 port map( A => A(11), B => n22, Y => 
                           A_shifter_11_port);
   SHIFTER_A_i_12 : AND2_89 port map( A => A(12), B => n23, Y => 
                           A_shifter_12_port);
   SHIFTER_A_i_13 : AND2_88 port map( A => A(13), B => n23, Y => 
                           A_shifter_13_port);
   SHIFTER_A_i_14 : AND2_87 port map( A => A(14), B => n23, Y => 
                           A_shifter_14_port);
   SHIFTER_A_i_15 : AND2_86 port map( A => A(15), B => n23, Y => 
                           A_shifter_15_port);
   SHIFTER_A_i_16 : AND2_85 port map( A => A(16), B => n23, Y => 
                           A_shifter_16_port);
   SHIFTER_A_i_17 : AND2_84 port map( A => A(17), B => n23, Y => 
                           A_shifter_17_port);
   SHIFTER_A_i_18 : AND2_83 port map( A => A(18), B => n23, Y => 
                           A_shifter_18_port);
   SHIFTER_A_i_19 : AND2_82 port map( A => A(19), B => n23, Y => 
                           A_shifter_19_port);
   SHIFTER_A_i_20 : AND2_81 port map( A => A(20), B => n23, Y => 
                           A_shifter_20_port);
   SHIFTER_A_i_21 : AND2_80 port map( A => A(21), B => n23, Y => 
                           A_shifter_21_port);
   SHIFTER_A_i_22 : AND2_79 port map( A => A(22), B => n23, Y => 
                           A_shifter_22_port);
   SHIFTER_A_i_23 : AND2_78 port map( A => A(23), B => n23, Y => 
                           A_shifter_23_port);
   SHIFTER_A_i_24 : AND2_77 port map( A => A(24), B => n24, Y => 
                           A_shifter_24_port);
   SHIFTER_A_i_25 : AND2_76 port map( A => A(25), B => n24, Y => 
                           A_shifter_25_port);
   SHIFTER_A_i_26 : AND2_75 port map( A => A(26), B => n24, Y => 
                           A_shifter_26_port);
   SHIFTER_A_i_27 : AND2_74 port map( A => A(27), B => n24, Y => 
                           A_shifter_27_port);
   SHIFTER_A_i_28 : AND2_73 port map( A => A(28), B => n24, Y => 
                           A_shifter_28_port);
   SHIFTER_A_i_29 : AND2_72 port map( A => A(29), B => n24, Y => 
                           A_shifter_29_port);
   SHIFTER_A_i_30 : AND2_71 port map( A => A(30), B => n24, Y => 
                           A_shifter_30_port);
   SHIFTER_A_i_31 : AND2_70 port map( A => A(31), B => n24, Y => 
                           A_shifter_31_port);
   SHIFTER_B_i_0 : AND2_69 port map( A => B(0), B => n24, Y => B_shifter_0_port
                           );
   SHIFTER_B_i_1 : AND2_68 port map( A => B(1), B => n24, Y => B_shifter_1_port
                           );
   SHIFTER_B_i_2 : AND2_67 port map( A => B(2), B => n24, Y => B_shifter_2_port
                           );
   SHIFTER_B_i_3 : AND2_66 port map( A => B(3), B => n24, Y => B_shifter_3_port
                           );
   SHIFTER_B_i_4 : AND2_65 port map( A => B(4), B => n24, Y => B_shifter_4_port
                           );
   SUM_i_0 : AND2_64 port map( A => out_adder_0_port, B => n1, Y => 
                           in_cmp_0_port);
   SUM_i_1 : AND2_63 port map( A => out_adder_1_port, B => n20, Y => 
                           in_cmp_1_port);
   SUM_i_2 : AND2_62 port map( A => out_adder_2_port, B => n20, Y => 
                           in_cmp_2_port);
   SUM_i_3 : AND2_61 port map( A => out_adder_3_port, B => n20, Y => 
                           in_cmp_3_port);
   SUM_i_4 : AND2_60 port map( A => out_adder_4_port, B => n20, Y => 
                           in_cmp_4_port);
   SUM_i_5 : AND2_59 port map( A => out_adder_5_port, B => n20, Y => 
                           in_cmp_5_port);
   SUM_i_6 : AND2_58 port map( A => out_adder_6_port, B => n20, Y => 
                           in_cmp_6_port);
   SUM_i_7 : AND2_57 port map( A => out_adder_7_port, B => n20, Y => 
                           in_cmp_7_port);
   SUM_i_8 : AND2_56 port map( A => out_adder_8_port, B => n20, Y => 
                           in_cmp_8_port);
   SUM_i_9 : AND2_55 port map( A => out_adder_9_port, B => n20, Y => 
                           in_cmp_9_port);
   SUM_i_10 : AND2_54 port map( A => out_adder_10_port, B => n20, Y => 
                           in_cmp_10_port);
   SUM_i_11 : AND2_53 port map( A => out_adder_11_port, B => n20, Y => 
                           in_cmp_11_port);
   SUM_i_12 : AND2_52 port map( A => out_adder_12_port, B => n20, Y => 
                           in_cmp_12_port);
   SUM_i_13 : AND2_51 port map( A => out_adder_13_port, B => n20, Y => 
                           in_cmp_13_port);
   SUM_i_14 : AND2_50 port map( A => out_adder_14_port, B => n20, Y => 
                           in_cmp_14_port);
   SUM_i_15 : AND2_49 port map( A => out_adder_15_port, B => n20, Y => 
                           in_cmp_15_port);
   SUM_i_16 : AND2_48 port map( A => out_adder_16_port, B => n20, Y => 
                           in_cmp_16_port);
   SUM_i_17 : AND2_47 port map( A => out_adder_17_port, B => n19, Y => 
                           in_cmp_17_port);
   SUM_i_18 : AND2_46 port map( A => out_adder_18_port, B => n19, Y => 
                           in_cmp_18_port);
   SUM_i_19 : AND2_45 port map( A => out_adder_19_port, B => n19, Y => 
                           in_cmp_19_port);
   SUM_i_20 : AND2_44 port map( A => out_adder_20_port, B => n19, Y => 
                           in_cmp_20_port);
   SUM_i_21 : AND2_43 port map( A => out_adder_21_port, B => n19, Y => 
                           in_cmp_21_port);
   SUM_i_22 : AND2_42 port map( A => out_adder_22_port, B => n19, Y => 
                           in_cmp_22_port);
   SUM_i_23 : AND2_41 port map( A => out_adder_23_port, B => n19, Y => 
                           in_cmp_23_port);
   SUM_i_24 : AND2_40 port map( A => out_adder_24_port, B => n19, Y => 
                           in_cmp_24_port);
   SUM_i_25 : AND2_39 port map( A => out_adder_25_port, B => n19, Y => 
                           in_cmp_25_port);
   SUM_i_26 : AND2_38 port map( A => out_adder_26_port, B => n19, Y => 
                           in_cmp_26_port);
   SUM_i_27 : AND2_37 port map( A => out_adder_27_port, B => n19, Y => 
                           in_cmp_27_port);
   SUM_i_28 : AND2_36 port map( A => out_adder_28_port, B => n19, Y => 
                           in_cmp_28_port);
   SUM_i_29 : AND2_35 port map( A => out_adder_29_port, B => n19, Y => 
                           in_cmp_29_port);
   SUM_i_30 : AND2_34 port map( A => out_adder_30_port, B => n19, Y => 
                           in_cmp_30_port);
   SUM_i_31 : AND2_33 port map( A => out_adder_31_port, B => n19, Y => 
                           in_cmp_31_port);
   MUL_A_i_0 : AND2_32 port map( A => A(0), B => n25, Y => A_mul_0_port);
   MUL_B_i_0 : AND2_31 port map( A => B(0), B => n25, Y => B_mul_0_port);
   MUL_A_i_1 : AND2_30 port map( A => A(1), B => n25, Y => A_mul_1_port);
   MUL_B_i_1 : AND2_29 port map( A => B(1), B => n25, Y => B_mul_1_port);
   MUL_A_i_2 : AND2_28 port map( A => A(2), B => n25, Y => A_mul_2_port);
   MUL_B_i_2 : AND2_27 port map( A => B(2), B => n25, Y => B_mul_2_port);
   MUL_A_i_3 : AND2_26 port map( A => A(3), B => n25, Y => A_mul_3_port);
   MUL_B_i_3 : AND2_25 port map( A => B(3), B => n25, Y => B_mul_3_port);
   MUL_A_i_4 : AND2_24 port map( A => A(4), B => n25, Y => A_mul_4_port);
   MUL_B_i_4 : AND2_23 port map( A => B(4), B => n25, Y => B_mul_4_port);
   MUL_A_i_5 : AND2_22 port map( A => A(5), B => n25, Y => A_mul_5_port);
   MUL_B_i_5 : AND2_21 port map( A => B(5), B => n25, Y => B_mul_5_port);
   MUL_A_i_6 : AND2_20 port map( A => A(6), B => n26, Y => A_mul_6_port);
   MUL_B_i_6 : AND2_19 port map( A => B(6), B => n26, Y => B_mul_6_port);
   MUL_A_i_7 : AND2_18 port map( A => A(7), B => n26, Y => A_mul_7_port);
   MUL_B_i_7 : AND2_17 port map( A => B(7), B => n26, Y => B_mul_7_port);
   MUL_A_i_8 : AND2_16 port map( A => A(8), B => n26, Y => A_mul_8_port);
   MUL_B_i_8 : AND2_15 port map( A => B(8), B => n26, Y => B_mul_8_port);
   MUL_A_i_9 : AND2_14 port map( A => A(9), B => n26, Y => A_mul_9_port);
   MUL_B_i_9 : AND2_13 port map( A => B(9), B => n26, Y => B_mul_9_port);
   MUL_A_i_10 : AND2_12 port map( A => A(10), B => n26, Y => A_mul_10_port);
   MUL_B_i_10 : AND2_11 port map( A => B(10), B => n26, Y => B_mul_10_port);
   MUL_A_i_11 : AND2_10 port map( A => A(11), B => n26, Y => A_mul_11_port);
   MUL_B_i_11 : AND2_9 port map( A => B(11), B => n26, Y => B_mul_11_port);
   MUL_A_i_12 : AND2_8 port map( A => A(12), B => n27, Y => A_mul_12_port);
   MUL_B_i_12 : AND2_7 port map( A => B(12), B => n27, Y => B_mul_12_port);
   MUL_A_i_13 : AND2_6 port map( A => A(13), B => n27, Y => A_mul_13_port);
   MUL_B_i_13 : AND2_5 port map( A => B(13), B => n27, Y => B_mul_13_port);
   MUL_A_i_14 : AND2_4 port map( A => A(14), B => n27, Y => A_mul_14_port);
   MUL_B_i_14 : AND2_3 port map( A => B(14), B => n27, Y => B_mul_14_port);
   MUL_A_i_15 : AND2_2 port map( A => A(15), B => n27, Y => A_mul_15_port);
   MUL_B_i_15 : AND2_1 port map( A => B(15), B => n27, Y => B_mul_15_port);
   ADD : ADDER_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A_adder_31_port, 
                           A(30) => A_adder_30_port, A(29) => A_adder_29_port, 
                           A(28) => A_adder_28_port, A(27) => A_adder_27_port, 
                           A(26) => A_adder_26_port, A(25) => A_adder_25_port, 
                           A(24) => A_adder_24_port, A(23) => A_adder_23_port, 
                           A(22) => A_adder_22_port, A(21) => A_adder_21_port, 
                           A(20) => A_adder_20_port, A(19) => A_adder_19_port, 
                           A(18) => A_adder_18_port, A(17) => A_adder_17_port, 
                           A(16) => A_adder_16_port, A(15) => A_adder_15_port, 
                           A(14) => A_adder_14_port, A(13) => A_adder_13_port, 
                           A(12) => A_adder_12_port, A(11) => A_adder_11_port, 
                           A(10) => A_adder_10_port, A(9) => A_adder_9_port, 
                           A(8) => A_adder_8_port, A(7) => A_adder_7_port, A(6)
                           => A_adder_6_port, A(5) => A_adder_5_port, A(4) => 
                           A_adder_4_port, A(3) => A_adder_3_port, A(2) => 
                           A_adder_2_port, A(1) => A_adder_1_port, A(0) => 
                           A_adder_0_port, B(31) => B_adder_31_port, B(30) => 
                           B_adder_30_port, B(29) => B_adder_29_port, B(28) => 
                           B_adder_28_port, B(27) => B_adder_27_port, B(26) => 
                           B_adder_26_port, B(25) => B_adder_25_port, B(24) => 
                           B_adder_24_port, B(23) => B_adder_23_port, B(22) => 
                           B_adder_22_port, B(21) => B_adder_21_port, B(20) => 
                           B_adder_20_port, B(19) => B_adder_19_port, B(18) => 
                           B_adder_18_port, B(17) => B_adder_17_port, B(16) => 
                           B_adder_16_port, B(15) => B_adder_15_port, B(14) => 
                           B_adder_14_port, B(13) => B_adder_13_port, B(12) => 
                           B_adder_12_port, B(11) => B_adder_11_port, B(10) => 
                           B_adder_10_port, B(9) => B_adder_9_port, B(8) => 
                           B_adder_8_port, B(7) => B_adder_7_port, B(6) => 
                           B_adder_6_port, B(5) => B_adder_5_port, B(4) => 
                           B_adder_4_port, B(3) => B_adder_3_port, B(2) => 
                           B_adder_2_port, B(1) => B_adder_1_port, B(0) => 
                           B_adder_0_port, ADD_SUB => n68, Cin => cin_internal,
                           S(31) => out_adder_31_port, S(30) => 
                           out_adder_30_port, S(29) => out_adder_29_port, S(28)
                           => out_adder_28_port, S(27) => out_adder_27_port, 
                           S(26) => out_adder_26_port, S(25) => 
                           out_adder_25_port, S(24) => out_adder_24_port, S(23)
                           => out_adder_23_port, S(22) => out_adder_22_port, 
                           S(21) => out_adder_21_port, S(20) => 
                           out_adder_20_port, S(19) => out_adder_19_port, S(18)
                           => out_adder_18_port, S(17) => out_adder_17_port, 
                           S(16) => out_adder_16_port, S(15) => 
                           out_adder_15_port, S(14) => out_adder_14_port, S(13)
                           => out_adder_13_port, S(12) => out_adder_12_port, 
                           S(11) => out_adder_11_port, S(10) => 
                           out_adder_10_port, S(9) => out_adder_9_port, S(8) =>
                           out_adder_8_port, S(7) => out_adder_7_port, S(6) => 
                           out_adder_6_port, S(5) => out_adder_5_port, S(4) => 
                           out_adder_4_port, S(3) => out_adder_3_port, S(2) => 
                           out_adder_2_port, S(1) => out_adder_1_port, S(0) => 
                           out_adder_0_port, Cout => Cout_port);
   SHIFT : SHIFTER port map( data_in(31) => A_shifter_31_port, data_in(30) => 
                           A_shifter_30_port, data_in(29) => A_shifter_29_port,
                           data_in(28) => A_shifter_28_port, data_in(27) => 
                           A_shifter_27_port, data_in(26) => A_shifter_26_port,
                           data_in(25) => A_shifter_25_port, data_in(24) => 
                           A_shifter_24_port, data_in(23) => A_shifter_23_port,
                           data_in(22) => A_shifter_22_port, data_in(21) => 
                           A_shifter_21_port, data_in(20) => A_shifter_20_port,
                           data_in(19) => A_shifter_19_port, data_in(18) => 
                           A_shifter_18_port, data_in(17) => A_shifter_17_port,
                           data_in(16) => A_shifter_16_port, data_in(15) => 
                           A_shifter_15_port, data_in(14) => A_shifter_14_port,
                           data_in(13) => A_shifter_13_port, data_in(12) => 
                           A_shifter_12_port, data_in(11) => A_shifter_11_port,
                           data_in(10) => A_shifter_10_port, data_in(9) => 
                           A_shifter_9_port, data_in(8) => A_shifter_8_port, 
                           data_in(7) => A_shifter_7_port, data_in(6) => 
                           A_shifter_6_port, data_in(5) => A_shifter_5_port, 
                           data_in(4) => A_shifter_4_port, data_in(3) => 
                           A_shifter_3_port, data_in(2) => A_shifter_2_port, 
                           data_in(1) => A_shifter_1_port, data_in(0) => 
                           A_shifter_0_port, R(4) => B_shifter_4_port, R(3) => 
                           B_shifter_3_port, R(2) => B_shifter_2_port, R(1) => 
                           B_shifter_1_port, R(0) => B_shifter_0_port, conf(1) 
                           => conf_1_port, conf(0) => conf_0_port, data_out(31)
                           => out_shifter_31_port, data_out(30) => 
                           out_shifter_30_port, data_out(29) => 
                           out_shifter_29_port, data_out(28) => 
                           out_shifter_28_port, data_out(27) => 
                           out_shifter_27_port, data_out(26) => 
                           out_shifter_26_port, data_out(25) => 
                           out_shifter_25_port, data_out(24) => 
                           out_shifter_24_port, data_out(23) => 
                           out_shifter_23_port, data_out(22) => 
                           out_shifter_22_port, data_out(21) => 
                           out_shifter_21_port, data_out(20) => 
                           out_shifter_20_port, data_out(19) => 
                           out_shifter_19_port, data_out(18) => 
                           out_shifter_18_port, data_out(17) => 
                           out_shifter_17_port, data_out(16) => 
                           out_shifter_16_port, data_out(15) => 
                           out_shifter_15_port, data_out(14) => 
                           out_shifter_14_port, data_out(13) => 
                           out_shifter_13_port, data_out(12) => 
                           out_shifter_12_port, data_out(11) => 
                           out_shifter_11_port, data_out(10) => 
                           out_shifter_10_port, data_out(9) => 
                           out_shifter_9_port, data_out(8) => 
                           out_shifter_8_port, data_out(7) => 
                           out_shifter_7_port, data_out(6) => 
                           out_shifter_6_port, data_out(5) => 
                           out_shifter_5_port, data_out(4) => 
                           out_shifter_4_port, data_out(3) => 
                           out_shifter_3_port, data_out(2) => 
                           out_shifter_2_port, data_out(1) => 
                           out_shifter_1_port, data_out(0) => 
                           out_shifter_0_port);
   LOGICALS : LOGIC_NBIT32_N_SELECTOR4 port map( S(3) => logic_sel_3_port, S(2)
                           => logic_sel_2_port, S(1) => logic_sel_1_port, S(0) 
                           => logic_sel_0_port, A(31) => A_logic_31_port, A(30)
                           => A_logic_30_port, A(29) => A_logic_29_port, A(28) 
                           => A_logic_28_port, A(27) => A_logic_27_port, A(26) 
                           => A_logic_26_port, A(25) => A_logic_25_port, A(24) 
                           => A_logic_24_port, A(23) => A_logic_23_port, A(22) 
                           => A_logic_22_port, A(21) => A_logic_21_port, A(20) 
                           => A_logic_20_port, A(19) => A_logic_19_port, A(18) 
                           => A_logic_18_port, A(17) => A_logic_17_port, A(16) 
                           => A_logic_16_port, A(15) => A_logic_15_port, A(14) 
                           => A_logic_14_port, A(13) => A_logic_13_port, A(12) 
                           => A_logic_12_port, A(11) => A_logic_11_port, A(10) 
                           => A_logic_10_port, A(9) => A_logic_9_port, A(8) => 
                           A_logic_8_port, A(7) => A_logic_7_port, A(6) => 
                           A_logic_6_port, A(5) => A_logic_5_port, A(4) => 
                           A_logic_4_port, A(3) => A_logic_3_port, A(2) => 
                           A_logic_2_port, A(1) => A_logic_1_port, A(0) => 
                           A_logic_0_port, B(31) => B_logic_31_port, B(30) => 
                           B_logic_30_port, B(29) => B_logic_29_port, B(28) => 
                           B_logic_28_port, B(27) => B_logic_27_port, B(26) => 
                           B_logic_26_port, B(25) => B_logic_25_port, B(24) => 
                           B_logic_24_port, B(23) => B_logic_23_port, B(22) => 
                           B_logic_22_port, B(21) => B_logic_21_port, B(20) => 
                           B_logic_20_port, B(19) => B_logic_19_port, B(18) => 
                           B_logic_18_port, B(17) => B_logic_17_port, B(16) => 
                           B_logic_16_port, B(15) => B_logic_15_port, B(14) => 
                           B_logic_14_port, B(13) => B_logic_13_port, B(12) => 
                           B_logic_12_port, B(11) => B_logic_11_port, B(10) => 
                           B_logic_10_port, B(9) => B_logic_9_port, B(8) => 
                           B_logic_8_port, B(7) => B_logic_7_port, B(6) => 
                           B_logic_6_port, B(5) => B_logic_5_port, B(4) => 
                           B_logic_4_port, B(3) => B_logic_3_port, B(2) => 
                           B_logic_2_port, B(1) => B_logic_1_port, B(0) => 
                           B_logic_0_port, O(31) => out_logic_31_port, O(30) =>
                           out_logic_30_port, O(29) => out_logic_29_port, O(28)
                           => out_logic_28_port, O(27) => out_logic_27_port, 
                           O(26) => out_logic_26_port, O(25) => 
                           out_logic_25_port, O(24) => out_logic_24_port, O(23)
                           => out_logic_23_port, O(22) => out_logic_22_port, 
                           O(21) => out_logic_21_port, O(20) => 
                           out_logic_20_port, O(19) => out_logic_19_port, O(18)
                           => out_logic_18_port, O(17) => out_logic_17_port, 
                           O(16) => out_logic_16_port, O(15) => 
                           out_logic_15_port, O(14) => out_logic_14_port, O(13)
                           => out_logic_13_port, O(12) => out_logic_12_port, 
                           O(11) => out_logic_11_port, O(10) => 
                           out_logic_10_port, O(9) => out_logic_9_port, O(8) =>
                           out_logic_8_port, O(7) => out_logic_7_port, O(6) => 
                           out_logic_6_port, O(5) => out_logic_5_port, O(4) => 
                           out_logic_4_port, O(3) => out_logic_3_port, O(2) => 
                           out_logic_2_port, O(1) => out_logic_1_port, O(0) => 
                           out_logic_0_port);
   COMPARATOR : CMP_NBIT32 port map( SUM(31) => in_cmp_31_port, SUM(30) => 
                           in_cmp_30_port, SUM(29) => in_cmp_29_port, SUM(28) 
                           => in_cmp_28_port, SUM(27) => in_cmp_27_port, 
                           SUM(26) => in_cmp_26_port, SUM(25) => in_cmp_25_port
                           , SUM(24) => in_cmp_24_port, SUM(23) => 
                           in_cmp_23_port, SUM(22) => in_cmp_22_port, SUM(21) 
                           => in_cmp_21_port, SUM(20) => in_cmp_20_port, 
                           SUM(19) => in_cmp_19_port, SUM(18) => in_cmp_18_port
                           , SUM(17) => in_cmp_17_port, SUM(16) => 
                           in_cmp_16_port, SUM(15) => in_cmp_15_port, SUM(14) 
                           => in_cmp_14_port, SUM(13) => in_cmp_13_port, 
                           SUM(12) => in_cmp_12_port, SUM(11) => in_cmp_11_port
                           , SUM(10) => in_cmp_10_port, SUM(9) => in_cmp_9_port
                           , SUM(8) => in_cmp_8_port, SUM(7) => in_cmp_7_port, 
                           SUM(6) => in_cmp_6_port, SUM(5) => in_cmp_5_port, 
                           SUM(4) => in_cmp_4_port, SUM(3) => in_cmp_3_port, 
                           SUM(2) => in_cmp_2_port, SUM(1) => in_cmp_1_port, 
                           SUM(0) => in_cmp_0_port, Cout => Cout_port, A_L_B =>
                           COND(0), A_LE_B => COND(1), A_G_B => COND(2), A_GE_B
                           => COND(3), A_E_B => COND(4), A_NE_B => COND(5));
   MULTIPLIER : MUL port map( CLOCK => CLOCK, A(15) => A_mul_15_port, A(14) => 
                           A_mul_14_port, A(13) => A_mul_13_port, A(12) => 
                           A_mul_12_port, A(11) => A_mul_11_port, A(10) => 
                           A_mul_10_port, A(9) => A_mul_9_port, A(8) => 
                           A_mul_8_port, A(7) => A_mul_7_port, A(6) => 
                           A_mul_6_port, A(5) => A_mul_5_port, A(4) => 
                           A_mul_4_port, A(3) => A_mul_3_port, A(2) => 
                           A_mul_2_port, A(1) => A_mul_1_port, A(0) => 
                           A_mul_0_port, B(15) => B_mul_15_port, B(14) => 
                           B_mul_14_port, B(13) => B_mul_13_port, B(12) => 
                           B_mul_12_port, B(11) => B_mul_11_port, B(10) => 
                           B_mul_10_port, B(9) => B_mul_9_port, B(8) => 
                           B_mul_8_port, B(7) => B_mul_7_port, B(6) => 
                           B_mul_6_port, B(5) => B_mul_5_port, B(4) => 
                           B_mul_4_port, B(3) => B_mul_3_port, B(2) => 
                           B_mul_2_port, B(1) => B_mul_1_port, B(0) => 
                           B_mul_0_port, Y(31) => out_mul_31_port, Y(30) => 
                           out_mul_30_port, Y(29) => out_mul_29_port, Y(28) => 
                           out_mul_28_port, Y(27) => out_mul_27_port, Y(26) => 
                           out_mul_26_port, Y(25) => out_mul_25_port, Y(24) => 
                           out_mul_24_port, Y(23) => out_mul_23_port, Y(22) => 
                           out_mul_22_port, Y(21) => out_mul_21_port, Y(20) => 
                           out_mul_20_port, Y(19) => out_mul_19_port, Y(18) => 
                           out_mul_18_port, Y(17) => out_mul_17_port, Y(16) => 
                           out_mul_16_port, Y(15) => out_mul_15_port, Y(14) => 
                           out_mul_14_port, Y(13) => out_mul_13_port, Y(12) => 
                           out_mul_12_port, Y(11) => out_mul_11_port, Y(10) => 
                           out_mul_10_port, Y(9) => out_mul_9_port, Y(8) => 
                           out_mul_8_port, Y(7) => out_mul_7_port, Y(6) => 
                           out_mul_6_port, Y(5) => out_mul_5_port, Y(4) => 
                           out_mul_4_port, Y(3) => out_mul_3_port, Y(2) => 
                           out_mul_2_port, Y(1) => out_mul_1_port, Y(0) => 
                           out_mul_0_port);
   OUTPUT_SEL : MUX4to1_NBIT32_1 port map( A(31) => out_adder_31_port, A(30) =>
                           out_adder_30_port, A(29) => out_adder_29_port, A(28)
                           => out_adder_28_port, A(27) => out_adder_27_port, 
                           A(26) => out_adder_26_port, A(25) => 
                           out_adder_25_port, A(24) => out_adder_24_port, A(23)
                           => out_adder_23_port, A(22) => out_adder_22_port, 
                           A(21) => out_adder_21_port, A(20) => 
                           out_adder_20_port, A(19) => out_adder_19_port, A(18)
                           => out_adder_18_port, A(17) => out_adder_17_port, 
                           A(16) => out_adder_16_port, A(15) => 
                           out_adder_15_port, A(14) => out_adder_14_port, A(13)
                           => out_adder_13_port, A(12) => out_adder_12_port, 
                           A(11) => out_adder_11_port, A(10) => 
                           out_adder_10_port, A(9) => out_adder_9_port, A(8) =>
                           out_adder_8_port, A(7) => out_adder_7_port, A(6) => 
                           out_adder_6_port, A(5) => out_adder_5_port, A(4) => 
                           out_adder_4_port, A(3) => out_adder_3_port, A(2) => 
                           out_adder_2_port, A(1) => out_adder_1_port, A(0) => 
                           out_adder_0_port, B(31) => out_logic_31_port, B(30) 
                           => out_logic_30_port, B(29) => out_logic_29_port, 
                           B(28) => out_logic_28_port, B(27) => 
                           out_logic_27_port, B(26) => out_logic_26_port, B(25)
                           => out_logic_25_port, B(24) => out_logic_24_port, 
                           B(23) => out_logic_23_port, B(22) => 
                           out_logic_22_port, B(21) => out_logic_21_port, B(20)
                           => out_logic_20_port, B(19) => out_logic_19_port, 
                           B(18) => out_logic_18_port, B(17) => 
                           out_logic_17_port, B(16) => out_logic_16_port, B(15)
                           => out_logic_15_port, B(14) => out_logic_14_port, 
                           B(13) => out_logic_13_port, B(12) => 
                           out_logic_12_port, B(11) => out_logic_11_port, B(10)
                           => out_logic_10_port, B(9) => out_logic_9_port, B(8)
                           => out_logic_8_port, B(7) => out_logic_7_port, B(6) 
                           => out_logic_6_port, B(5) => out_logic_5_port, B(4) 
                           => out_logic_4_port, B(3) => out_logic_3_port, B(2) 
                           => out_logic_2_port, B(1) => out_logic_1_port, B(0) 
                           => out_logic_0_port, C(31) => out_shifter_31_port, 
                           C(30) => out_shifter_30_port, C(29) => 
                           out_shifter_29_port, C(28) => out_shifter_28_port, 
                           C(27) => out_shifter_27_port, C(26) => 
                           out_shifter_26_port, C(25) => out_shifter_25_port, 
                           C(24) => out_shifter_24_port, C(23) => 
                           out_shifter_23_port, C(22) => out_shifter_22_port, 
                           C(21) => out_shifter_21_port, C(20) => 
                           out_shifter_20_port, C(19) => out_shifter_19_port, 
                           C(18) => out_shifter_18_port, C(17) => 
                           out_shifter_17_port, C(16) => out_shifter_16_port, 
                           C(15) => out_shifter_15_port, C(14) => 
                           out_shifter_14_port, C(13) => out_shifter_13_port, 
                           C(12) => out_shifter_12_port, C(11) => 
                           out_shifter_11_port, C(10) => out_shifter_10_port, 
                           C(9) => out_shifter_9_port, C(8) => 
                           out_shifter_8_port, C(7) => out_shifter_7_port, C(6)
                           => out_shifter_6_port, C(5) => out_shifter_5_port, 
                           C(4) => out_shifter_4_port, C(3) => 
                           out_shifter_3_port, C(2) => out_shifter_2_port, C(1)
                           => out_shifter_1_port, C(0) => out_shifter_0_port, 
                           D(31) => out_mul_31_port, D(30) => out_mul_30_port, 
                           D(29) => out_mul_29_port, D(28) => out_mul_28_port, 
                           D(27) => out_mul_27_port, D(26) => out_mul_26_port, 
                           D(25) => out_mul_25_port, D(24) => out_mul_24_port, 
                           D(23) => out_mul_23_port, D(22) => out_mul_22_port, 
                           D(21) => out_mul_21_port, D(20) => out_mul_20_port, 
                           D(19) => out_mul_19_port, D(18) => out_mul_18_port, 
                           D(17) => out_mul_17_port, D(16) => out_mul_16_port, 
                           D(15) => out_mul_15_port, D(14) => out_mul_14_port, 
                           D(13) => out_mul_13_port, D(12) => out_mul_12_port, 
                           D(11) => out_mul_11_port, D(10) => out_mul_10_port, 
                           D(9) => out_mul_9_port, D(8) => out_mul_8_port, D(7)
                           => out_mul_7_port, D(6) => out_mul_6_port, D(5) => 
                           out_mul_5_port, D(4) => out_mul_4_port, D(3) => 
                           out_mul_3_port, D(2) => out_mul_2_port, D(1) => 
                           out_mul_1_port, D(0) => out_mul_0_port, SEL(1) => 
                           mux_out_1_port, SEL(0) => mux_out_0_port, Y(31) => 
                           ALU_out(31), Y(30) => ALU_out(30), Y(29) => 
                           ALU_out(29), Y(28) => ALU_out(28), Y(27) => 
                           ALU_out(27), Y(26) => ALU_out(26), Y(25) => 
                           ALU_out(25), Y(24) => ALU_out(24), Y(23) => 
                           ALU_out(23), Y(22) => ALU_out(22), Y(21) => 
                           ALU_out(21), Y(20) => ALU_out(20), Y(19) => 
                           ALU_out(19), Y(18) => ALU_out(18), Y(17) => 
                           ALU_out(17), Y(16) => ALU_out(16), Y(15) => 
                           ALU_out(15), Y(14) => ALU_out(14), Y(13) => 
                           ALU_out(13), Y(12) => ALU_out(12), Y(11) => 
                           ALU_out(11), Y(10) => ALU_out(10), Y(9) => 
                           ALU_out(9), Y(8) => ALU_out(8), Y(7) => ALU_out(7), 
                           Y(6) => ALU_out(6), Y(5) => ALU_out(5), Y(4) => 
                           ALU_out(4), Y(3) => ALU_out(3), Y(2) => ALU_out(2), 
                           Y(1) => ALU_out(1), Y(0) => ALU_out(0));
   U3 : BUF_X1 port map( A => n3, Z => n31);
   U4 : BUF_X1 port map( A => n18, Z => n14);
   U5 : BUF_X1 port map( A => en_adder, Z => n13);
   U6 : NAND2_X1 port map( A1 => n54, A2 => n48, ZN => n1);
   U7 : BUF_X1 port map( A => n31, Z => n30);
   U8 : BUF_X1 port map( A => n17, Z => n15);
   U9 : BUF_X1 port map( A => n69, Z => n24);
   U10 : BUF_X1 port map( A => n13, Z => n17);
   U11 : BUF_X1 port map( A => n69, Z => n22);
   U12 : BUF_X1 port map( A => n69, Z => n23);
   U13 : BUF_X1 port map( A => n70, Z => n26);
   U14 : BUF_X1 port map( A => n70, Z => n25);
   U15 : BUF_X1 port map( A => n70, Z => n27);
   U16 : BUF_X1 port map( A => n1, Z => n20);
   U17 : BUF_X1 port map( A => n1, Z => n19);
   U18 : INV_X1 port map( A => n30, ZN => n28);
   U19 : INV_X1 port map( A => n30, ZN => n29);
   U20 : AND2_X1 port map( A1 => n51, A2 => n46, ZN => n2);
   U21 : AOI211_X1 port map( C1 => n5, C2 => n63, A => n62, B => n61, ZN => N90
                           );
   U22 : INV_X1 port map( A => AluOpcode(0), ZN => n57);
   U23 : AND2_X1 port map( A1 => n55, A2 => n54, ZN => n8);
   U24 : BUF_X1 port map( A => AluOpcode(0), Z => n7);
   U25 : AND3_X1 port map( A1 => n64, A2 => n37, A3 => n36, ZN => n3);
   U26 : NAND2_X1 port map( A1 => n56, A2 => n8, ZN => en_adder);
   U27 : CLKBUF_X1 port map( A => n17, Z => n4);
   U28 : CLKBUF_X1 port map( A => n13, Z => n18);
   U29 : CLKBUF_X1 port map( A => n17, Z => n16);
   U30 : BUF_X1 port map( A => n6, Z => n5);
   U31 : BUF_X1 port map( A => AluOpcode(2), Z => n6);
   U32 : NAND2_X1 port map( A1 => AluOpcode(2), A2 => AluOpcode(3), ZN => n9);
   U33 : OR2_X1 port map( A1 => n9, A2 => n7, ZN => n10);
   U34 : CLKBUF_X1 port map( A => AluOpcode(3), Z => n11);
   U35 : NAND2_X1 port map( A1 => n56, A2 => n8, ZN => n67);
   U36 : NOR2_X1 port map( A1 => n32, A2 => n7, ZN => n12);
   U37 : XNOR2_X1 port map( A => n50, B => n58, ZN => n52);
   U38 : NOR2_X1 port map( A1 => n6, A2 => n53, ZN => n50);
   U39 : NOR2_X1 port map( A1 => n7, A2 => AluOpcode(1), ZN => n21);
   U40 : AND4_X1 port map( A1 => Cin, A2 => AluOpcode(3), A3 => n44, A4 => n57,
                           ZN => cin_internal);
   U41 : NAND2_X1 port map( A1 => n7, A2 => AluOpcode(3), ZN => n59);
   U42 : INV_X1 port map( A => AluOpcode(1), ZN => n51);
   U43 : INV_X1 port map( A => AluOpcode(2), ZN => n46);
   U44 : INV_X1 port map( A => AluOpcode(4), ZN => n53);
   U45 : NAND2_X1 port map( A1 => n2, A2 => n53, ZN => n33);
   U46 : NAND2_X1 port map( A1 => AluOpcode(2), A2 => AluOpcode(3), ZN => n32);
   U47 : INV_X1 port map( A => n9, ZN => n45);
   U48 : NAND2_X1 port map( A1 => AluOpcode(1), A2 => AluOpcode(4), ZN => n42);
   U49 : INV_X1 port map( A => AluOpcode(3), ZN => n58);
   U50 : NAND3_X1 port map( A1 => n6, A2 => n58, A3 => n57, ZN => n43);
   U51 : NAND2_X1 port map( A1 => AluOpcode(4), A2 => n51, ZN => n61);
   U52 : OAI222_X1 port map( A1 => n59, A2 => n33, B1 => n10, B2 => n42, C1 => 
                           n43, C2 => n61, ZN => N89);
   U53 : INV_X1 port map( A => n33, ZN => n44);
   U54 : NOR3_X1 port map( A1 => n5, A2 => AluOpcode(3), A3 => n61, ZN => n34);
   U55 : OAI21_X1 port map( B1 => n44, B2 => n34, A => n7, ZN => n64);
   U56 : INV_X1 port map( A => N89, ZN => n37);
   U57 : NAND2_X1 port map( A1 => n46, A2 => n57, ZN => n60);
   U58 : INV_X1 port map( A => n60, ZN => n35);
   U59 : INV_X1 port map( A => n61, ZN => n39);
   U60 : NAND3_X1 port map( A1 => n35, A2 => AluOpcode(3), A3 => n39, ZN => n36
                           );
   U61 : INV_X1 port map( A => n59, ZN => n38);
   U62 : NAND3_X1 port map( A1 => n39, A2 => n38, A3 => n46, ZN => n65);
   U63 : NAND2_X1 port map( A1 => n65, A2 => n31, ZN => mux_out_0_port);
   U64 : INV_X1 port map( A => n43, ZN => n40);
   U65 : NAND2_X1 port map( A1 => n40, A2 => n61, ZN => n49);
   U66 : NAND2_X1 port map( A1 => n49, A2 => n65, ZN => mux_out_1_port);
   U67 : AOI22_X1 port map( A1 => n21, A2 => n53, B1 => AluOpcode(1), B2 => n5,
                           ZN => n41);
   U68 : OAI22_X1 port map( A1 => n11, A2 => n41, B1 => n2, B2 => n57, ZN => 
                           N91);
   U69 : NOR2_X1 port map( A1 => n43, A2 => n42, ZN => N92);
   U70 : NOR3_X1 port map( A1 => AluOpcode(1), A2 => AluOpcode(4), A3 => n43, 
                           ZN => N93);
   U71 : NAND3_X1 port map( A1 => n53, A2 => n57, A3 => n45, ZN => n47);
   U72 : NAND3_X1 port map( A1 => AluOpcode(1), A2 => n46, A3 => n57, ZN => n54
                           );
   U73 : NAND2_X1 port map( A1 => n12, A2 => n51, ZN => n48);
   U74 : NAND3_X1 port map( A1 => n47, A2 => n54, A3 => n48, ZN => n68);
   U75 : INV_X1 port map( A => n49, ZN => n69);
   U76 : NAND3_X1 port map( A1 => n57, A2 => n52, A3 => n51, ZN => n56);
   U77 : NAND3_X1 port map( A1 => AluOpcode(3), A2 => n57, A3 => n53, ZN => n55
                           );
   U78 : NAND2_X1 port map( A1 => n56, A2 => n8, ZN => n66);
   U79 : NAND2_X1 port map( A1 => n58, A2 => n57, ZN => n63);
   U80 : OAI21_X1 port map( B1 => n11, B2 => n60, A => n59, ZN => n62);
   U81 : INV_X1 port map( A => n64, ZN => N88);
   U82 : INV_X1 port map( A => n65, ZN => n70);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT5 is

   port( A, B, C : in std_logic_vector (4 downto 0);  SEL : in std_logic_vector
         (1 downto 0);  Y : out std_logic_vector (4 downto 0));

end MUX3to1_NBIT5;

architecture SYN_Behavioral of MUX3to1_NBIT5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n7, n8, n9, n10, n11, n12_port, n13, n14, n1, n2, n3, n4, n5, n6
      : std_logic;

begin
   
   Y_reg_4_inst : DLH_X1 port map( G => N12, D => n1, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => N12, D => n2, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => N12, D => n3, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => n4, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => n5, Q => Y(0));
   U3 : NOR2_X1 port map( A1 => n6, A2 => SEL(0), ZN => n9);
   U4 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n8);
   U5 : AND2_X1 port map( A1 => SEL(0), A2 => n6, ZN => n10);
   U6 : NAND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => N12);
   U7 : INV_X1 port map( A => SEL(1), ZN => n6);
   U8 : INV_X1 port map( A => n14, ZN => n5);
   U9 : AOI222_X1 port map( A1 => A(0), A2 => n8, B1 => C(0), B2 => n9, C1 => 
                           B(0), C2 => n10, ZN => n14);
   U10 : INV_X1 port map( A => n13, ZN => n4);
   U11 : AOI222_X1 port map( A1 => A(1), A2 => n8, B1 => C(1), B2 => n9, C1 => 
                           B(1), C2 => n10, ZN => n13);
   U12 : INV_X1 port map( A => n12_port, ZN => n3);
   U13 : AOI222_X1 port map( A1 => A(2), A2 => n8, B1 => C(2), B2 => n9, C1 => 
                           B(2), C2 => n10, ZN => n12_port);
   U14 : INV_X1 port map( A => n11, ZN => n2);
   U15 : AOI222_X1 port map( A1 => A(3), A2 => n8, B1 => C(3), B2 => n9, C1 => 
                           B(3), C2 => n10, ZN => n11);
   U16 : INV_X1 port map( A => n7, ZN => n1);
   U17 : AOI222_X1 port map( A1 => A(4), A2 => n8, B1 => C(4), B2 => n9, C1 => 
                           B(4), C2 => n10, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX4to1_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX4to1_NBIT32_0;

architecture SYN_Behavioral of MUX4to1_NBIT32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n7, Z => n72);
   U2 : BUF_X1 port map( A => n6, Z => n76);
   U3 : BUF_X1 port map( A => n4, Z => n81);
   U4 : BUF_X1 port map( A => n5, Z => n77);
   U5 : BUF_X1 port map( A => n76, Z => n73);
   U6 : BUF_X1 port map( A => n76, Z => n74);
   U7 : BUF_X1 port map( A => n81, Z => n82);
   U8 : BUF_X1 port map( A => n81, Z => n83);
   U9 : BUF_X1 port map( A => n72, Z => n1);
   U10 : BUF_X1 port map( A => n72, Z => n70);
   U11 : BUF_X1 port map( A => n77, Z => n78);
   U12 : BUF_X1 port map( A => n77, Z => n79);
   U13 : BUF_X1 port map( A => n76, Z => n75);
   U14 : BUF_X1 port map( A => n81, Z => n84);
   U15 : BUF_X1 port map( A => n72, Z => n71);
   U16 : BUF_X1 port map( A => n77, Z => n80);
   U17 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(0));
   U18 : AOI22_X1 port map( A1 => D(0), A2 => n82, B1 => C(0), B2 => n78, ZN =>
                           n69);
   U19 : AOI22_X1 port map( A1 => B(0), A2 => n73, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U20 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(8));
   U21 : AOI22_X1 port map( A1 => D(8), A2 => n84, B1 => C(8), B2 => n80, ZN =>
                           n9);
   U22 : AOI22_X1 port map( A1 => B(8), A2 => n75, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U23 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(10));
   U24 : AOI22_X1 port map( A1 => D(10), A2 => n82, B1 => C(10), B2 => n78, ZN 
                           => n67);
   U25 : AOI22_X1 port map( A1 => B(10), A2 => n73, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U26 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(11));
   U27 : AOI22_X1 port map( A1 => D(11), A2 => n82, B1 => C(11), B2 => n78, ZN 
                           => n65);
   U28 : AOI22_X1 port map( A1 => B(11), A2 => n73, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U29 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(13));
   U30 : AOI22_X1 port map( A1 => D(13), A2 => n82, B1 => C(13), B2 => n78, ZN 
                           => n61);
   U31 : AOI22_X1 port map( A1 => B(13), A2 => n73, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U32 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(14));
   U33 : AOI22_X1 port map( A1 => D(14), A2 => n82, B1 => C(14), B2 => n78, ZN 
                           => n59);
   U34 : AOI22_X1 port map( A1 => B(14), A2 => n73, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U35 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(1));
   U36 : AOI22_X1 port map( A1 => D(1), A2 => n82, B1 => C(1), B2 => n78, ZN =>
                           n47);
   U37 : AOI22_X1 port map( A1 => B(1), A2 => n73, B1 => A(1), B2 => n1, ZN => 
                           n46);
   U38 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(2));
   U39 : AOI22_X1 port map( A1 => D(2), A2 => n83, B1 => C(2), B2 => n79, ZN =>
                           n25);
   U40 : AOI22_X1 port map( A1 => B(2), A2 => n74, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U41 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(3));
   U42 : AOI22_X1 port map( A1 => D(3), A2 => n84, B1 => C(3), B2 => n80, ZN =>
                           n19);
   U43 : AOI22_X1 port map( A1 => B(3), A2 => n75, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U44 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(4));
   U45 : AOI22_X1 port map( A1 => D(4), A2 => n84, B1 => C(4), B2 => n80, ZN =>
                           n17);
   U46 : AOI22_X1 port map( A1 => B(4), A2 => n75, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U47 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(5));
   U48 : AOI22_X1 port map( A1 => D(5), A2 => n84, B1 => C(5), B2 => n80, ZN =>
                           n15);
   U49 : AOI22_X1 port map( A1 => B(5), A2 => n75, B1 => A(5), B2 => n71, ZN =>
                           n14);
   U50 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(6));
   U51 : AOI22_X1 port map( A1 => D(6), A2 => n84, B1 => C(6), B2 => n80, ZN =>
                           n13);
   U52 : AOI22_X1 port map( A1 => B(6), A2 => n75, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U53 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(7));
   U54 : AOI22_X1 port map( A1 => D(7), A2 => n84, B1 => C(7), B2 => n80, ZN =>
                           n11);
   U55 : AOI22_X1 port map( A1 => B(7), A2 => n75, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U56 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(9));
   U57 : AOI22_X1 port map( A1 => D(9), A2 => n84, B1 => C(9), B2 => n80, ZN =>
                           n3);
   U58 : AOI22_X1 port map( A1 => B(9), A2 => n75, B1 => A(9), B2 => n71, ZN =>
                           n2);
   U59 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(12));
   U60 : AOI22_X1 port map( A1 => D(12), A2 => n82, B1 => C(12), B2 => n78, ZN 
                           => n63);
   U61 : AOI22_X1 port map( A1 => B(12), A2 => n73, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U62 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(15));
   U63 : AOI22_X1 port map( A1 => D(15), A2 => n82, B1 => C(15), B2 => n78, ZN 
                           => n57);
   U64 : AOI22_X1 port map( A1 => B(15), A2 => n73, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U65 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => D(28), A2 => n83, B1 => C(28), B2 => n79, ZN 
                           => n29);
   U67 : AOI22_X1 port map( A1 => B(28), A2 => n74, B1 => A(28), B2 => n70, ZN 
                           => n28);
   U68 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(16));
   U69 : AOI22_X1 port map( A1 => D(16), A2 => n82, B1 => C(16), B2 => n78, ZN 
                           => n55);
   U70 : AOI22_X1 port map( A1 => B(16), A2 => n73, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U71 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(17));
   U72 : AOI22_X1 port map( A1 => D(17), A2 => n82, B1 => C(17), B2 => n78, ZN 
                           => n53);
   U73 : AOI22_X1 port map( A1 => B(17), A2 => n73, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U74 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(18));
   U75 : AOI22_X1 port map( A1 => D(18), A2 => n82, B1 => C(18), B2 => n78, ZN 
                           => n51);
   U76 : AOI22_X1 port map( A1 => B(18), A2 => n73, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U77 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(19));
   U78 : AOI22_X1 port map( A1 => D(19), A2 => n82, B1 => C(19), B2 => n78, ZN 
                           => n49);
   U79 : AOI22_X1 port map( A1 => B(19), A2 => n73, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U80 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(20));
   U81 : AOI22_X1 port map( A1 => D(20), A2 => n83, B1 => C(20), B2 => n79, ZN 
                           => n45);
   U82 : AOI22_X1 port map( A1 => B(20), A2 => n74, B1 => A(20), B2 => n70, ZN 
                           => n44);
   U83 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(21));
   U84 : AOI22_X1 port map( A1 => D(21), A2 => n83, B1 => C(21), B2 => n79, ZN 
                           => n43);
   U85 : AOI22_X1 port map( A1 => B(21), A2 => n74, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U86 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(22));
   U87 : AOI22_X1 port map( A1 => D(22), A2 => n83, B1 => C(22), B2 => n79, ZN 
                           => n41);
   U88 : AOI22_X1 port map( A1 => B(22), A2 => n74, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U89 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(23));
   U90 : AOI22_X1 port map( A1 => D(23), A2 => n83, B1 => C(23), B2 => n79, ZN 
                           => n39);
   U91 : AOI22_X1 port map( A1 => B(23), A2 => n74, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U92 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(24));
   U93 : AOI22_X1 port map( A1 => D(24), A2 => n83, B1 => C(24), B2 => n79, ZN 
                           => n37);
   U94 : AOI22_X1 port map( A1 => B(24), A2 => n74, B1 => A(24), B2 => n70, ZN 
                           => n36);
   U95 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(25));
   U96 : AOI22_X1 port map( A1 => D(25), A2 => n83, B1 => C(25), B2 => n79, ZN 
                           => n35);
   U97 : AOI22_X1 port map( A1 => B(25), A2 => n74, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U98 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(26));
   U99 : AOI22_X1 port map( A1 => D(26), A2 => n83, B1 => C(26), B2 => n79, ZN 
                           => n33);
   U100 : AOI22_X1 port map( A1 => B(26), A2 => n74, B1 => A(26), B2 => n70, ZN
                           => n32);
   U101 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(27));
   U102 : AOI22_X1 port map( A1 => D(27), A2 => n83, B1 => C(27), B2 => n79, ZN
                           => n31);
   U103 : AOI22_X1 port map( A1 => B(27), A2 => n74, B1 => A(27), B2 => n70, ZN
                           => n30);
   U104 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(29));
   U105 : AOI22_X1 port map( A1 => D(29), A2 => n83, B1 => C(29), B2 => n79, ZN
                           => n27);
   U106 : AOI22_X1 port map( A1 => B(29), A2 => n74, B1 => A(29), B2 => n70, ZN
                           => n26);
   U107 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(30));
   U108 : AOI22_X1 port map( A1 => D(30), A2 => n83, B1 => C(30), B2 => n79, ZN
                           => n23);
   U109 : AOI22_X1 port map( A1 => B(30), A2 => n74, B1 => A(30), B2 => n70, ZN
                           => n22);
   U110 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(31));
   U111 : AOI22_X1 port map( A1 => D(31), A2 => n84, B1 => C(31), B2 => n80, ZN
                           => n21);
   U112 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n71, ZN
                           => n20);
   U113 : NOR2_X1 port map( A1 => n85, A2 => SEL(1), ZN => n6);
   U114 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n7);
   U115 : INV_X1 port map( A => SEL(0), ZN => n85);
   U116 : AND2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n4);
   U117 : AND2_X1 port map( A1 => SEL(1), A2 => n85, ZN => n5);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT2 is

   port( A, B, C, SEL : in std_logic_vector (1 downto 0);  Y : out 
         std_logic_vector (1 downto 0));

end MUX3to1_NBIT2;

architecture SYN_Behavioral of MUX3to1_NBIT2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, N13, N14, n2, n3, n4, n5, n1 : std_logic;

begin
   
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => N14, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => N13, Q => Y(0));
   U9 : NAND3_X1 port map( A1 => C(1), A2 => n1, A3 => SEL(1), ZN => n3);
   U10 : NAND3_X1 port map( A1 => SEL(1), A2 => n1, A3 => C(0), ZN => n5);
   U3 : INV_X1 port map( A => SEL(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => N12);
   U5 : OAI21_X1 port map( B1 => SEL(1), B2 => n4, A => n5, ZN => N13);
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => SEL(0), ZN 
                           => n4);
   U7 : OAI21_X1 port map( B1 => SEL(1), B2 => n2, A => n3, ZN => N14);
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => SEL(0), B2 => B(1), ZN 
                           => n2);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_0 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_0;

architecture SYN_Behavioral of MUX5to1_NBIT32_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n1, n2, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
      n94, n95, n96 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n91, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n92, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n92, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n93, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n93, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n94);
   U4 : BUF_X1 port map( A => n7, Z => n82);
   U5 : BUF_X1 port map( A => n5, Z => n90);
   U6 : BUF_X1 port map( A => n8, Z => n78);
   U7 : BUF_X1 port map( A => n9, Z => n74);
   U8 : BUF_X1 port map( A => n6, Z => n83);
   U9 : BUF_X1 port map( A => n94, Z => n92);
   U10 : BUF_X1 port map( A => n94, Z => n91);
   U11 : BUF_X1 port map( A => n94, Z => n93);
   U12 : OR4_X1 port map( A1 => n86, A2 => n81, A3 => n72, A4 => n89, ZN => N25
                           );
   U13 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n72);
   U14 : BUF_X1 port map( A => n78, Z => n76);
   U15 : BUF_X1 port map( A => n78, Z => n75);
   U16 : BUF_X1 port map( A => n74, Z => n2);
   U17 : BUF_X1 port map( A => n74, Z => n1);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n80);
   U21 : BUF_X1 port map( A => n82, Z => n79);
   U22 : BUF_X1 port map( A => n90, Z => n88);
   U23 : BUF_X1 port map( A => n90, Z => n87);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : BUF_X1 port map( A => n74, Z => n73);
   U26 : BUF_X1 port map( A => n83, Z => n86);
   U27 : BUF_X1 port map( A => n82, Z => n81);
   U28 : BUF_X1 port map( A => n90, Z => n89);
   U29 : INV_X1 port map( A => SEL(1), ZN => n96);
   U30 : INV_X1 port map( A => SEL(0), ZN => n95);
   U31 : NOR3_X1 port map( A1 => n95, A2 => SEL(2), A3 => n96, ZN => n7);
   U32 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n96, ZN => n5);
   U33 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n95, ZN => n8);
   U34 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n9);
   U35 : AND3_X1 port map( A1 => n95, A2 => n96, A3 => SEL(2), ZN => n6);
   U36 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U37 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN =>
                           n70);
   U38 : AOI222_X1 port map( A1 => C(0), A2 => n89, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n81, ZN => n71);
   U39 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U40 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN =>
                           n68);
   U41 : AOI222_X1 port map( A1 => C(1), A2 => n89, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n81, ZN => n69);
   U42 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U43 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN =>
                           n66);
   U44 : AOI222_X1 port map( A1 => C(2), A2 => n89, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n81, ZN => n67);
   U45 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U46 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN =>
                           n64);
   U47 : AOI222_X1 port map( A1 => C(3), A2 => n89, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n81, ZN => n65);
   U48 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U49 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN =>
                           n62);
   U50 : AOI222_X1 port map( A1 => C(4), A2 => n89, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n81, ZN => n63);
   U51 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U52 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n60);
   U53 : AOI222_X1 port map( A1 => C(5), A2 => n89, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n81, ZN => n61);
   U54 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U55 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n58);
   U56 : AOI222_X1 port map( A1 => C(6), A2 => n89, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n81, ZN => n59);
   U57 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U58 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n56_port);
   U59 : AOI222_X1 port map( A1 => C(7), A2 => n89, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n81, ZN => n57_port);
   U60 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U61 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n54_port);
   U62 : AOI222_X1 port map( A1 => C(8), A2 => n88, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n80, ZN => n55_port);
   U63 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U64 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n52_port);
   U65 : AOI222_X1 port map( A1 => C(9), A2 => n88, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n80, ZN => n53_port);
   U66 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U67 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n50_port);
   U68 : AOI222_X1 port map( A1 => C(10), A2 => n88, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n80, ZN => n51_port);
   U69 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U70 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n48_port);
   U71 : AOI222_X1 port map( A1 => C(11), A2 => n88, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n49_port);
   U72 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U73 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n46_port);
   U74 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n47_port);
   U75 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U76 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n44_port);
   U77 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n45_port);
   U78 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U79 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n42_port);
   U80 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n43_port);
   U81 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U82 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n40_port);
   U83 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n41_port);
   U84 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U85 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n38_port);
   U86 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n39_port);
   U87 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U88 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n36_port);
   U89 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n37_port);
   U90 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U91 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n34_port);
   U92 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n35_port);
   U93 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U94 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n32_port);
   U95 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n33_port);
   U96 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U97 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n30_port);
   U98 : AOI222_X1 port map( A1 => C(20), A2 => n87, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n79, ZN => n31_port);
   U99 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U100 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n28_port);
   U101 : AOI222_X1 port map( A1 => C(21), A2 => n87, B1 => E(21), B2 => n84, 
                           C1 => D(21), C2 => n79, ZN => n29_port);
   U102 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U103 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n26_port);
   U104 : AOI222_X1 port map( A1 => C(22), A2 => n87, B1 => E(22), B2 => n84, 
                           C1 => D(22), C2 => n79, ZN => n27_port);
   U105 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U106 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n24);
   U107 : AOI222_X1 port map( A1 => C(23), A2 => n87, B1 => E(23), B2 => n84, 
                           C1 => D(23), C2 => n79, ZN => n25_port);
   U108 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U109 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n22);
   U110 : AOI222_X1 port map( A1 => C(24), A2 => n87, B1 => E(24), B2 => n84, 
                           C1 => D(24), C2 => n79, ZN => n23);
   U111 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U112 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n20);
   U113 : AOI222_X1 port map( A1 => C(25), A2 => n87, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n79, ZN => n21);
   U114 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U115 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n18);
   U116 : AOI222_X1 port map( A1 => C(26), A2 => n87, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n79, ZN => n19);
   U117 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U118 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n16);
   U119 : AOI222_X1 port map( A1 => C(27), A2 => n87, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n79, ZN => n17);
   U120 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U121 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n14);
   U122 : AOI222_X1 port map( A1 => C(28), A2 => n87, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n79, ZN => n15);
   U123 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U124 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n12);
   U125 : AOI222_X1 port map( A1 => C(29), A2 => n87, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n79, ZN => n13);
   U126 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U127 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n10);
   U128 : AOI222_X1 port map( A1 => C(30), A2 => n87, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n79, ZN => n11);
   U129 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U130 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n3);
   U131 : AOI222_X1 port map( A1 => C(31), A2 => n87, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n79, ZN => n4);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_0;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : CLKBUF_X3 port map( A => SEL, Z => n1);
   U2 : BUF_X2 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U5 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U6 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U8 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U9 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U11 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U12 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U13 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U14 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U15 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U16 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U17 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U20 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U21 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U22 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U23 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U24 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U26 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U27 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U28 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U29 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U30 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U31 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U32 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U33 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U34 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U35 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_0 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_0;

architecture SYN_Behavioral of MUX3to1_NBIT32_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12_port, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
      , n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n16, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n17, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n18, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n27, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n28, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n73, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(0));
   U3 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U4 : BUF_X1 port map( A => n35, Z => n12_port);
   U5 : BUF_X1 port map( A => n36, Z => n8);
   U6 : BUF_X1 port map( A => n37, Z => n1);
   U7 : BUF_X1 port map( A => N12, Z => n14);
   U8 : BUF_X1 port map( A => N12, Z => n13);
   U9 : BUF_X1 port map( A => N12, Z => n15);
   U10 : BUF_X1 port map( A => n8, Z => n6);
   U11 : BUF_X1 port map( A => n8, Z => n5);
   U12 : BUF_X1 port map( A => n1, Z => n2);
   U13 : BUF_X1 port map( A => n1, Z => n3);
   U14 : BUF_X1 port map( A => n12_port, Z => n9);
   U15 : BUF_X1 port map( A => n12_port, Z => n10);
   U16 : BUF_X1 port map( A => n8, Z => n7);
   U17 : BUF_X1 port map( A => n1, Z => n4);
   U18 : BUF_X1 port map( A => n12_port, Z => n11);
   U19 : INV_X1 port map( A => SEL(1), ZN => n83);
   U20 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n35);
   U21 : NOR2_X1 port map( A1 => n83, A2 => SEL(0), ZN => n36);
   U22 : AND2_X1 port map( A1 => SEL(0), A2 => n83, ZN => n37);
   U23 : INV_X1 port map( A => n68, ZN => n82);
   U24 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n68);
   U25 : INV_X1 port map( A => n67, ZN => n81);
   U26 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n67);
   U27 : INV_X1 port map( A => n66, ZN => n80);
   U28 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n66);
   U29 : INV_X1 port map( A => n65, ZN => n79);
   U30 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n65);
   U31 : INV_X1 port map( A => n64, ZN => n78);
   U32 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n64);
   U33 : INV_X1 port map( A => n63, ZN => n77);
   U34 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n63);
   U35 : INV_X1 port map( A => n62, ZN => n76);
   U36 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n62);
   U37 : INV_X1 port map( A => n61, ZN => n75);
   U38 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n61);
   U39 : INV_X1 port map( A => n60, ZN => n74);
   U40 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n60);
   U41 : INV_X1 port map( A => n59, ZN => n73);
   U42 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n59);
   U43 : INV_X1 port map( A => n58, ZN => n72);
   U44 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n58);
   U45 : INV_X1 port map( A => n57, ZN => n71);
   U46 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n57);
   U47 : INV_X1 port map( A => n56, ZN => n70);
   U48 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n56);
   U49 : INV_X1 port map( A => n55, ZN => n69);
   U50 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n55);
   U51 : INV_X1 port map( A => n54, ZN => n33);
   U52 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n54);
   U53 : INV_X1 port map( A => n53, ZN => n32);
   U54 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n53);
   U55 : INV_X1 port map( A => n52, ZN => n31);
   U56 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n52);
   U57 : INV_X1 port map( A => n51, ZN => n30);
   U58 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n51);
   U59 : INV_X1 port map( A => n50, ZN => n29);
   U60 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n50);
   U61 : INV_X1 port map( A => n49, ZN => n28);
   U62 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n49);
   U63 : INV_X1 port map( A => n48, ZN => n27);
   U64 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n48);
   U65 : INV_X1 port map( A => n47, ZN => n26);
   U66 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n47);
   U67 : INV_X1 port map( A => n46, ZN => n25);
   U68 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n46);
   U69 : INV_X1 port map( A => n45, ZN => n24);
   U70 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n45);
   U71 : INV_X1 port map( A => n44, ZN => n23);
   U72 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n44);
   U73 : INV_X1 port map( A => n43, ZN => n22);
   U74 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n43);
   U75 : INV_X1 port map( A => n42, ZN => n21);
   U76 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n42);
   U77 : INV_X1 port map( A => n41, ZN => n20);
   U78 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n41);
   U79 : INV_X1 port map( A => n40, ZN => n19);
   U80 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n40);
   U81 : INV_X1 port map( A => n39, ZN => n18);
   U82 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n39);
   U83 : INV_X1 port map( A => n38, ZN => n17);
   U84 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n38);
   U85 : INV_X1 port map( A => n34, ZN => n16);
   U86 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n34);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Sum : out std_logic_vector 
         (31 downto 0));

end PC_adder_0;

architecture SYN_Behavioral of PC_adder_0 is

   component PC_adder_0_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1734 : std_logic;

begin
   
   n1 <= '0';
   add_16 : PC_adder_0_DW01_add_1 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(31) => Sum(31), 
                           SUM(30) => Sum(30), SUM(29) => Sum(29), SUM(28) => 
                           Sum(28), SUM(27) => Sum(27), SUM(26) => Sum(26), 
                           SUM(25) => Sum(25), SUM(24) => Sum(24), SUM(23) => 
                           Sum(23), SUM(22) => Sum(22), SUM(21) => Sum(21), 
                           SUM(20) => Sum(20), SUM(19) => Sum(19), SUM(18) => 
                           Sum(18), SUM(17) => Sum(17), SUM(16) => Sum(16), 
                           SUM(15) => Sum(15), SUM(14) => Sum(14), SUM(13) => 
                           Sum(13), SUM(12) => Sum(12), SUM(11) => Sum(11), 
                           SUM(10) => Sum(10), SUM(9) => Sum(9), SUM(8) => 
                           Sum(8), SUM(7) => Sum(7), SUM(6) => Sum(6), SUM(5) 
                           => Sum(5), SUM(4) => Sum(4), SUM(3) => Sum(3), 
                           SUM(2) => Sum(2), SUM(1) => Sum(1), SUM(0) => Sum(0)
                           , CO => n_1734);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT7 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (6 
         downto 0);  data_out : out std_logic_vector (6 downto 0));

end REG_NBIT7;

architecture SYN_Behavioral of REG_NBIT7 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n8, n9, n10, n11, n12, n15, n16, n17, n18, n19, n20, n22
      , n1, n2, n3, n4, n5, n6, n7, data_out_5_port, data_out_6_port, n21, 
      n_1735, n_1736 : std_logic;

begin
   data_out <= ( data_out_6_port, data_out_5_port, data_out_4_port, 
      data_out_3_port, data_out_2_port, data_out_1_port, data_out_0_port );
   
   reg_reg_6_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n3, Q => 
                           data_out_6_port, QN => n_1735);
   reg_reg_5_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n3, Q => 
                           data_out_5_port, QN => n_1736);
   reg_reg_4_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n3, Q => 
                           data_out_4_port, QN => n12);
   reg_reg_3_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n3, Q => 
                           data_out_3_port, QN => n11);
   reg_reg_2_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n3, Q => 
                           data_out_2_port, QN => n10);
   reg_reg_1_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n3, Q => 
                           data_out_1_port, QN => n9);
   reg_reg_0_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n3, Q => 
                           data_out_0_port, QN => n8);
   U2 : INV_X1 port map( A => reset, ZN => n3);
   U3 : INV_X1 port map( A => n2, ZN => n1);
   U4 : INV_X1 port map( A => enable, ZN => n2);
   U5 : OAI22_X1 port map( A1 => n2, A2 => n4, B1 => n8, B2 => n1, ZN => n15);
   U6 : INV_X1 port map( A => data_in(0), ZN => n4);
   U7 : NAND2_X1 port map( A1 => data_in(1), A2 => n1, ZN => n5);
   U8 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n5, ZN => n16);
   U9 : NAND2_X1 port map( A1 => data_in(2), A2 => n1, ZN => n6);
   U10 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U11 : NAND2_X1 port map( A1 => data_in(3), A2 => n1, ZN => n7);
   U12 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n7, ZN => n18);
   U13 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n1, Z =>
                           n20);
   U14 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n1, Z =>
                           n22);
   U15 : NAND2_X1 port map( A1 => data_in(4), A2 => n1, ZN => n21);
   U16 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n21, ZN => n19);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FFD_0;

architecture SYN_BEHAVIORAL of FFD_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2, n4, n1, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n1, Q => Q, QN => n2);
   U2 : INV_X1 port map( A => RESET, ZN => n1);
   U3 : INV_X1 port map( A => n2, ZN => n3);
   U4 : MUX2_X1 port map( A => n3, B => D, S => ENABLE, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_0 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_0;

architecture SYN_Behavioral of REG_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n97, n1, n2, n3, n4, n5, data_out_0_port, data_out_1_port, 
      data_out_2_port, data_out_3_port, data_out_4_port, data_out_5_port, 
      data_out_6_port, data_out_7_port, data_out_8_port, data_out_9_port, 
      data_out_10_port, data_out_11_port, data_out_12_port, data_out_13_port, 
      data_out_14_port, data_out_15_port, data_out_16_port, data_out_17_port, 
      data_out_18_port, data_out_19_port, data_out_20_port, data_out_21_port, 
      data_out_22_port, data_out_23_port, data_out_24_port, data_out_25_port, 
      data_out_26_port, data_out_27_port, data_out_28_port, data_out_29_port, 
      data_out_30_port, data_out_31_port, n_1737, n_1738, n_1739, n_1740, 
      n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, 
      n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, 
      n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, 
      n_1768 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n5, Q => 
                           data_out_0_port, QN => n_1737);
   reg_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n5, Q => 
                           data_out_1_port, QN => n_1738);
   reg_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n5, Q => 
                           data_out_2_port, QN => n_1739);
   reg_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n5, Q => 
                           data_out_3_port, QN => n_1740);
   reg_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n5, Q => 
                           data_out_4_port, QN => n_1741);
   reg_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n5, Q => 
                           data_out_5_port, QN => n_1742);
   reg_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n5, Q => 
                           data_out_8_port, QN => n_1743);
   reg_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n5, Q => 
                           data_out_9_port, QN => n_1744);
   reg_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n5, Q => 
                           data_out_12_port, QN => n_1745);
   reg_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n5, Q => 
                           data_out_6_port, QN => n_1746);
   reg_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n5, Q => 
                           data_out_13_port, QN => n_1747);
   reg_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n5, Q => 
                           data_out_16_port, QN => n_1748);
   reg_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n5, Q => 
                           data_out_10_port, QN => n_1749);
   reg_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n5, Q => 
                           data_out_11_port, QN => n_1750);
   reg_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n5, Q => 
                           data_out_7_port, QN => n_1751);
   reg_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n5, Q => 
                           data_out_14_port, QN => n_1752);
   reg_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n5, Q => 
                           data_out_15_port, QN => n_1753);
   reg_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n5, Q => 
                           data_out_21_port, QN => n_1754);
   reg_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n5, Q => 
                           data_out_24_port, QN => n_1755);
   reg_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n5, Q => 
                           data_out_28_port, QN => n_1756);
   reg_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n5, Q => 
                           data_out_17_port, QN => n_1757);
   reg_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n5, Q => 
                           data_out_20_port, QN => n_1758);
   reg_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n5, Q => 
                           data_out_18_port, QN => n_1759);
   reg_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n5, Q => 
                           data_out_25_port, QN => n_1760);
   reg_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n5, Q => 
                           data_out_26_port, QN => n_1761);
   reg_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n5, Q => 
                           data_out_29_port, QN => n_1762);
   reg_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n5, Q => 
                           data_out_23_port, QN => n_1763);
   reg_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n5, Q => 
                           data_out_27_port, QN => n_1764);
   reg_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n5, Q => 
                           data_out_31_port, QN => n_1765);
   reg_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n5, Q => 
                           data_out_22_port, QN => n_1766);
   reg_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n5, Q => 
                           data_out_19_port, QN => n_1767);
   reg_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n5, Q => 
                           data_out_30_port, QN => n_1768);
   U2 : INV_X2 port map( A => reset, ZN => n5);
   U3 : BUF_X1 port map( A => enable, Z => n4);
   U4 : BUF_X1 port map( A => n4, Z => n3);
   U5 : BUF_X1 port map( A => n4, Z => n1);
   U6 : BUF_X1 port map( A => n4, Z => n2);
   U7 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => n1, Z => 
                           n65);
   U8 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n1, Z => 
                           n66);
   U9 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => n1, Z => 
                           n67);
   U10 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => n1, Z =>
                           n68);
   U11 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => n1, Z =>
                           n69);
   U12 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n1, Z =>
                           n70);
   U13 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n1, Z =>
                           n71);
   U14 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => n1, Z =>
                           n72);
   U15 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => n1, Z =>
                           n73);
   U16 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n1, Z =>
                           n74);
   U17 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => n1, Z 
                           => n75);
   U18 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => n1, Z 
                           => n76);
   U19 : MUX2_X1 port map( A => data_out_12_port, B => data_in(12), S => n2, Z 
                           => n77);
   U20 : MUX2_X1 port map( A => data_out_13_port, B => data_in(13), S => n2, Z 
                           => n78);
   U21 : MUX2_X1 port map( A => data_out_14_port, B => data_in(14), S => n2, Z 
                           => n79);
   U22 : MUX2_X1 port map( A => data_out_15_port, B => data_in(15), S => n2, Z 
                           => n80);
   U23 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => n2, Z 
                           => n81);
   U24 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => n2, Z 
                           => n82);
   U25 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => n2, Z 
                           => n83);
   U26 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => n2, Z 
                           => n84);
   U27 : MUX2_X1 port map( A => data_out_20_port, B => data_in(20), S => n2, Z 
                           => n85);
   U28 : MUX2_X1 port map( A => data_out_21_port, B => data_in(21), S => n2, Z 
                           => n86);
   U29 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => n2, Z 
                           => n87);
   U30 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => n2, Z 
                           => n88);
   U31 : MUX2_X1 port map( A => data_out_24_port, B => data_in(24), S => n3, Z 
                           => n89);
   U32 : MUX2_X1 port map( A => data_out_25_port, B => data_in(25), S => n3, Z 
                           => n90);
   U33 : MUX2_X1 port map( A => data_out_26_port, B => data_in(26), S => n3, Z 
                           => n91);
   U34 : MUX2_X1 port map( A => data_out_27_port, B => data_in(27), S => n3, Z 
                           => n92);
   U35 : MUX2_X1 port map( A => data_out_28_port, B => data_in(28), S => n3, Z 
                           => n93);
   U36 : MUX2_X1 port map( A => data_out_29_port, B => data_in(29), S => n3, Z 
                           => n94);
   U37 : MUX2_X1 port map( A => data_out_30_port, B => data_in(30), S => n3, Z 
                           => n95);
   U38 : MUX2_X1 port map( A => data_out_31_port, B => data_in(31), S => n3, Z 
                           => n97);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector (31 
         downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out std_logic_vector (31 
         downto 0);  BMP : inout std_logic;  STALL : out std_logic_vector (1 
         downto 0);  ID_EN, RF_RD, SIGND, IMM_SEL, BPR_EN : in std_logic;  
         ALU_OPCODE : in std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, ALUB_SEL,
         UCB_EN, MEM_EN, MEM_DATA_SEL : in std_logic;  LD_SEL : in 
         std_logic_vector (2 downto 0);  ALR2_SEL : in std_logic;  CWB_SEL : in
         std_logic_vector (1 downto 0);  WB_SEL, RF_WR : in std_logic;  
         RF_MUX_SEL : in std_logic_vector (1 downto 0));

end Datapath;

architecture SYN_BEHAVIORAL of Datapath is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RF_NBIT32_NREG32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component CWBU
      port( CLOCK : in std_logic;  ALU_OP : in std_logic_vector (0 to 4);  PSW 
            : in std_logic_vector (6 downto 0);  COND_SEL : out 
            std_logic_vector (1 downto 0);  CWB_SEL : in std_logic_vector (1 
            downto 0);  CWB_MUW_SEL : out std_logic_vector (1 downto 0));
   end component;
   
   component BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0
      port( clock, rst : in std_logic;  address : in std_logic_vector (31 
            downto 0);  d_in, w_en : in std_logic;  d_out : out std_logic);
   end component;
   
   component HDU_IR_SIZE32
      port( clk, rst : in std_logic;  IR : in std_logic_vector (31 downto 0);  
            STALL_CODE : out std_logic_vector (1 downto 0);  IF_STALL, ID_STALL
            , EX_STALL, MEM_STALL, WB_STALL : out std_logic);
   end component;
   
   component FWDU_IR_SIZE32
      port( CLOCK, RESET, EN : in std_logic;  IR : in std_logic_vector (31 
            downto 0);  FWD_A, FWD_B : out std_logic_vector (1 downto 0);  
            FWD_B2 : out std_logic;  ZDU_SEL : out std_logic_vector (1 downto 
            0));
   end component;
   
   component ALU_NBIT32
      port( CLOCK : in std_logic;  AluOpcode : in std_logic_vector (0 to 4);  A
            , B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            ALU_out : out std_logic_vector (31 downto 0);  Cout : out std_logic
            ;  COND : out std_logic_vector (5 downto 0));
   end component;
   
   component MUX3to1_NBIT5
      port( A, B, C : in std_logic_vector (4 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (4 downto 
            0));
   end component;
   
   component MUX2to1_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX4to1_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT2
      port( A, B, C, SEL : in std_logic_vector (1 downto 0);  Y : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component MUX2to1_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX5to1_NBIT32_0
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX2to1_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX3to1_NBIT32_1
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT32_2
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT32_3
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX2to1_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_8
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX3to1_NBIT32_0
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component PC_adder_1
      port( A, B : in std_logic_vector (31 downto 0);  Sum : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component PC_adder_0
      port( A, B : in std_logic_vector (31 downto 0);  Sum : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_4
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_5
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT7
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (6 downto 0);  data_out : out std_logic_vector (6 downto 0));
   end component;
   
   component REG_NBIT32_6
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_7
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_8
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_9
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_10
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component FFD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component REG_NBIT32_11
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_12
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component FFD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component REG_NBIT32_13
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_14
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_15
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_16
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_17
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_0
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IRAM_ADDR_31_port, IRAM_ADDR_30_port, 
      IRAM_ADDR_29_port, IRAM_ADDR_28_port, IRAM_ADDR_27_port, 
      IRAM_ADDR_26_port, IRAM_ADDR_25_port, IRAM_ADDR_24_port, 
      IRAM_ADDR_23_port, IRAM_ADDR_22_port, IRAM_ADDR_21_port, 
      IRAM_ADDR_20_port, IRAM_ADDR_19_port, IRAM_ADDR_18_port, 
      IRAM_ADDR_17_port, IRAM_ADDR_16_port, IRAM_ADDR_15_port, 
      IRAM_ADDR_14_port, IRAM_ADDR_13_port, IRAM_ADDR_12_port, 
      IRAM_ADDR_11_port, IRAM_ADDR_10_port, IRAM_ADDR_9_port, IRAM_ADDR_8_port,
      IRAM_ADDR_7_port, IRAM_ADDR_6_port, IRAM_ADDR_5_port, IRAM_ADDR_4_port, 
      IRAM_ADDR_3_port, IRAM_ADDR_2_port, IRAM_ADDR_1_port, IRAM_ADDR_0_port, 
      DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port, NPC_in_31_port, 
      NPC_in_30_port, NPC_in_29_port, NPC_in_28_port, NPC_in_27_port, 
      NPC_in_26_port, NPC_in_25_port, NPC_in_24_port, NPC_in_23_port, 
      NPC_in_22_port, NPC_in_21_port, NPC_in_20_port, NPC_in_19_port, 
      NPC_in_18_port, NPC_in_17_port, NPC_in_16_port, NPC_in_15_port, 
      NPC_in_14_port, NPC_in_13_port, NPC_in_12_port, NPC_in_11_port, 
      NPC_in_10_port, NPC_in_9_port, NPC_in_8_port, NPC_in_7_port, 
      NPC_in_6_port, NPC_in_5_port, NPC_in_4_port, NPC_in_3_port, NPC_in_2_port
      , NPC_in_1_port, NPC_in_0_port, PC_out_31_port, PC_out_30_port, 
      PC_out_29_port, PC_out_28_port, PC_out_27_port, PC_out_26_port, 
      PC_out_25_port, PC_out_24_port, PC_out_23_port, PC_out_22_port, 
      PC_out_21_port, PC_out_20_port, PC_out_19_port, PC_out_18_port, 
      PC_out_17_port, PC_out_16_port, PC_out_15_port, PC_out_14_port, 
      PC_out_13_port, PC_out_12_port, PC_out_11_port, PC_out_10_port, 
      PC_out_9_port, PC_out_8_port, PC_out_7_port, PC_out_6_port, PC_out_5_port
      , PC_out_4_port, PC_out_3_port, PC_out_2_port, PC_out_1_port, 
      PC_out_0_port, IR_out_31_port, IR_out_30_port, IR_out_29_port, 
      IR_out_28_port, IR_out_27_port, IR_out_26_port, IR_out_25_port, 
      IR_out_24_port, IR_out_23_port, IR_out_22_port, IR_out_21_port, 
      IR_out_20_port, IR_out_19_port, IR_out_18_port, IR_out_17_port, 
      IR_out_16_port, IR_out_15_port, IR_out_14_port, IR_out_13_port, 
      IR_out_12_port, IR_out_11_port, IR_out_10_port, IR_out_9_port, 
      IR_out_8_port, IR_out_7_port, IR_out_6_port, IR_out_5_port, IR_out_4_port
      , IR_out_3_port, IR_out_2_port, IR_out_1_port, IR_out_0_port, 
      NPC_out_31_port, NPC_out_30_port, NPC_out_29_port, NPC_out_28_port, 
      NPC_out_27_port, NPC_out_26_port, NPC_out_25_port, NPC_out_24_port, 
      NPC_out_23_port, NPC_out_22_port, NPC_out_21_port, NPC_out_20_port, 
      NPC_out_19_port, NPC_out_18_port, NPC_out_17_port, NPC_out_16_port, 
      NPC_out_15_port, NPC_out_14_port, NPC_out_13_port, NPC_out_12_port, 
      NPC_out_11_port, NPC_out_10_port, NPC_out_9_port, NPC_out_8_port, 
      NPC_out_7_port, NPC_out_6_port, NPC_out_5_port, NPC_out_4_port, 
      NPC_out_3_port, NPC_out_2_port, NPC_out_1_port, NPC_out_0_port, 
      PC2_out_31_port, PC2_out_30_port, PC2_out_29_port, PC2_out_28_port, 
      PC2_out_27_port, PC2_out_26_port, PC2_out_25_port, PC2_out_24_port, 
      PC2_out_23_port, PC2_out_22_port, PC2_out_21_port, PC2_out_20_port, 
      PC2_out_19_port, PC2_out_18_port, PC2_out_17_port, PC2_out_16_port, 
      PC2_out_15_port, PC2_out_14_port, PC2_out_13_port, PC2_out_12_port, 
      PC2_out_11_port, PC2_out_10_port, PC2_out_9_port, PC2_out_8_port, 
      PC2_out_7_port, PC2_out_6_port, PC2_out_5_port, PC2_out_4_port, 
      PC2_out_3_port, PC2_out_2_port, PC2_out_1_port, PC2_out_0_port, 
      RIMM_out_31_port, RIMM_out_30_port, RIMM_out_29_port, RIMM_out_28_port, 
      RIMM_out_27_port, RIMM_out_26_port, RIMM_out_25_port, RIMM_out_24_port, 
      RIMM_out_23_port, RIMM_out_22_port, RIMM_out_21_port, RIMM_out_20_port, 
      RIMM_out_19_port, RIMM_out_18_port, RIMM_out_17_port, RIMM_out_16_port, 
      RIMM_out_15_port, RIMM_out_14_port, RIMM_out_13_port, RIMM_out_12_port, 
      RIMM_out_11_port, RIMM_out_10_port, RIMM_out_9_port, RIMM_out_8_port, 
      RIMM_out_7_port, RIMM_out_6_port, RIMM_out_5_port, RIMM_out_4_port, 
      RIMM_out_3_port, RIMM_out_2_port, RIMM_out_1_port, RIMM_out_0_port, 
      RWB1_out_31_port, RWB1_out_30_port, RWB1_out_29_port, RWB1_out_28_port, 
      RWB1_out_27_port, RWB1_out_26_port, RWB1_out_25_port, RWB1_out_24_port, 
      RWB1_out_23_port, RWB1_out_22_port, RWB1_out_21_port, RWB1_out_20_port, 
      RWB1_out_19_port, RWB1_out_18_port, RWB1_out_17_port, RWB1_out_16_port, 
      RWB1_out_15_port, RWB1_out_14_port, RWB1_out_13_port, RWB1_out_12_port, 
      RWB1_out_11_port, RWB1_out_10_port, RWB1_out_9_port, RWB1_out_8_port, 
      RWB1_out_7_port, RWB1_out_6_port, RWB1_out_5_port, RWB1_out_4_port, 
      RWB1_out_3_port, RWB1_out_2_port, RWB1_out_1_port, RWB1_out_0_port, 
      BHT_out, PRD_OUT, NPC2_out_31_port, NPC2_out_30_port, NPC2_out_29_port, 
      NPC2_out_28_port, NPC2_out_27_port, NPC2_out_26_port, NPC2_out_25_port, 
      NPC2_out_24_port, NPC2_out_23_port, NPC2_out_22_port, NPC2_out_21_port, 
      NPC2_out_20_port, NPC2_out_19_port, NPC2_out_18_port, NPC2_out_17_port, 
      NPC2_out_16_port, NPC2_out_15_port, NPC2_out_14_port, NPC2_out_13_port, 
      NPC2_out_12_port, NPC2_out_11_port, NPC2_out_10_port, NPC2_out_9_port, 
      NPC2_out_8_port, NPC2_out_7_port, NPC2_out_6_port, NPC2_out_5_port, 
      NPC2_out_4_port, NPC2_out_3_port, NPC2_out_2_port, NPC2_out_1_port, 
      NPC2_out_0_port, JADDER_out_31_port, JADDER_out_30_port, 
      JADDER_out_29_port, JADDER_out_28_port, JADDER_out_27_port, 
      JADDER_out_26_port, JADDER_out_25_port, JADDER_out_24_port, 
      JADDER_out_23_port, JADDER_out_22_port, JADDER_out_21_port, 
      JADDER_out_20_port, JADDER_out_19_port, JADDER_out_18_port, 
      JADDER_out_17_port, JADDER_out_16_port, JADDER_out_15_port, 
      JADDER_out_14_port, JADDER_out_13_port, JADDER_out_12_port, 
      JADDER_out_11_port, JADDER_out_10_port, JADDER_out_9_port, 
      JADDER_out_8_port, JADDER_out_7_port, JADDER_out_6_port, 
      JADDER_out_5_port, JADDER_out_4_port, JADDER_out_3_port, 
      JADDER_out_2_port, JADDER_out_1_port, JADDER_out_0_port, 
      JADDER2_out_31_port, JADDER2_out_30_port, JADDER2_out_29_port, 
      JADDER2_out_28_port, JADDER2_out_27_port, JADDER2_out_26_port, 
      JADDER2_out_25_port, JADDER2_out_24_port, JADDER2_out_23_port, 
      JADDER2_out_22_port, JADDER2_out_21_port, JADDER2_out_20_port, 
      JADDER2_out_19_port, JADDER2_out_18_port, JADDER2_out_17_port, 
      JADDER2_out_16_port, JADDER2_out_15_port, JADDER2_out_14_port, 
      JADDER2_out_13_port, JADDER2_out_12_port, JADDER2_out_11_port, 
      JADDER2_out_10_port, JADDER2_out_9_port, JADDER2_out_8_port, 
      JADDER2_out_7_port, JADDER2_out_6_port, JADDER2_out_5_port, 
      JADDER2_out_4_port, JADDER2_out_3_port, JADDER2_out_2_port, 
      JADDER2_out_1_port, JADDER2_out_0_port, BPR_EN2, EX_ENABLE, 
      PC3_out_31_port, PC3_out_30_port, PC3_out_29_port, PC3_out_28_port, 
      PC3_out_27_port, PC3_out_26_port, PC3_out_25_port, PC3_out_24_port, 
      PC3_out_23_port, PC3_out_22_port, PC3_out_21_port, PC3_out_20_port, 
      PC3_out_19_port, PC3_out_18_port, PC3_out_17_port, PC3_out_16_port, 
      PC3_out_15_port, PC3_out_14_port, PC3_out_13_port, PC3_out_12_port, 
      PC3_out_11_port, PC3_out_10_port, PC3_out_9_port, PC3_out_8_port, 
      PC3_out_7_port, PC3_out_6_port, PC3_out_5_port, PC3_out_4_port, 
      PC3_out_3_port, PC3_out_2_port, PC3_out_1_port, PC3_out_0_port, 
      RWB2_out_31_port, RWB2_out_30_port, RWB2_out_29_port, RWB2_out_28_port, 
      RWB2_out_27_port, RWB2_out_26_port, RWB2_out_25_port, RWB2_out_24_port, 
      RWB2_out_23_port, RWB2_out_22_port, RWB2_out_21_port, RWB2_out_20_port, 
      RWB2_out_19_port, RWB2_out_18_port, RWB2_out_17_port, RWB2_out_16_port, 
      RWB2_out_15_port, RWB2_out_14_port, RWB2_out_13_port, RWB2_out_12_port, 
      RWB2_out_11_port, RWB2_out_10_port, RWB2_out_9_port, RWB2_out_8_port, 
      RWB2_out_7_port, RWB2_out_6_port, RWB2_out_5_port, RWB2_out_4_port, 
      RWB2_out_3_port, RWB2_out_2_port, RWB2_out_1_port, RWB2_out_0_port, 
      RB_out_31_port, RB_out_30_port, RB_out_29_port, RB_out_28_port, 
      RB_out_27_port, RB_out_26_port, RB_out_25_port, RB_out_24_port, 
      RB_out_23_port, RB_out_22_port, RB_out_21_port, RB_out_20_port, 
      RB_out_19_port, RB_out_18_port, RB_out_17_port, RB_out_16_port, 
      RB_out_15_port, RB_out_14_port, RB_out_13_port, RB_out_12_port, 
      RB_out_11_port, RB_out_10_port, RB_out_9_port, RB_out_8_port, 
      RB_out_7_port, RB_out_6_port, RB_out_5_port, RB_out_4_port, RB_out_3_port
      , RB_out_2_port, RB_out_1_port, RB_out_0_port, B2_out_31_port, 
      B2_out_30_port, B2_out_29_port, B2_out_28_port, B2_out_27_port, 
      B2_out_26_port, B2_out_25_port, B2_out_24_port, B2_out_23_port, 
      B2_out_22_port, B2_out_21_port, B2_out_20_port, B2_out_19_port, 
      B2_out_18_port, B2_out_17_port, B2_out_16_port, B2_out_15_port, 
      B2_out_14_port, B2_out_13_port, B2_out_12_port, B2_out_11_port, 
      B2_out_10_port, B2_out_9_port, B2_out_8_port, B2_out_7_port, 
      B2_out_6_port, B2_out_5_port, B2_out_4_port, B2_out_3_port, B2_out_2_port
      , B2_out_1_port, B2_out_0_port, ALR_in_31_port, ALR_in_30_port, 
      ALR_in_29_port, ALR_in_28_port, ALR_in_27_port, ALR_in_26_port, 
      ALR_in_25_port, ALR_in_24_port, ALR_in_23_port, ALR_in_22_port, 
      ALR_in_21_port, ALR_in_20_port, ALR_in_19_port, ALR_in_18_port, 
      ALR_in_17_port, ALR_in_16_port, ALR_in_15_port, ALR_in_14_port, 
      ALR_in_13_port, ALR_in_12_port, ALR_in_11_port, ALR_in_10_port, 
      ALR_in_9_port, ALR_in_8_port, ALR_in_7_port, ALR_in_6_port, ALR_in_5_port
      , ALR_in_4_port, ALR_in_3_port, ALR_in_2_port, ALR_in_1_port, 
      ALR_in_0_port, NPC3_out_31_port, NPC3_out_30_port, NPC3_out_29_port, 
      NPC3_out_28_port, NPC3_out_27_port, NPC3_out_26_port, NPC3_out_25_port, 
      NPC3_out_24_port, NPC3_out_23_port, NPC3_out_22_port, NPC3_out_21_port, 
      NPC3_out_20_port, NPC3_out_19_port, NPC3_out_18_port, NPC3_out_17_port, 
      NPC3_out_16_port, NPC3_out_15_port, NPC3_out_14_port, NPC3_out_13_port, 
      NPC3_out_12_port, NPC3_out_11_port, NPC3_out_10_port, NPC3_out_9_port, 
      NPC3_out_8_port, NPC3_out_7_port, NPC3_out_6_port, NPC3_out_5_port, 
      NPC3_out_4_port, NPC3_out_3_port, NPC3_out_2_port, NPC3_out_1_port, 
      NPC3_out_0_port, PSW_in_6_port, PSW_in_5_port, PSW_in_4_port, 
      PSW_in_3_port, PSW_in_2_port, PSW_in_1_port, PSW_in_0_port, 
      PSW_out_6_port, PSW_out_5_port, PSW_out_4_port, PSW_out_3_port, 
      PSW_out_2_port, PSW_out_1_port, PSW_out_0_port, MEM_ENABLE, 
      ALR2_in_31_port, ALR2_in_30_port, ALR2_in_29_port, ALR2_in_28_port, 
      ALR2_in_27_port, ALR2_in_26_port, ALR2_in_25_port, ALR2_in_24_port, 
      ALR2_in_23_port, ALR2_in_22_port, ALR2_in_21_port, ALR2_in_20_port, 
      ALR2_in_19_port, ALR2_in_18_port, ALR2_in_17_port, ALR2_in_16_port, 
      ALR2_in_15_port, ALR2_in_14_port, ALR2_in_13_port, ALR2_in_12_port, 
      ALR2_in_11_port, ALR2_in_10_port, ALR2_in_9_port, ALR2_in_8_port, 
      ALR2_in_7_port, ALR2_in_6_port, ALR2_in_5_port, ALR2_in_4_port, 
      ALR2_in_3_port, ALR2_in_2_port, ALR2_in_1_port, ALR2_in_0_port, 
      ALR2_out_31_port, ALR2_out_30_port, ALR2_out_29_port, ALR2_out_28_port, 
      ALR2_out_27_port, ALR2_out_26_port, ALR2_out_25_port, ALR2_out_24_port, 
      ALR2_out_23_port, ALR2_out_22_port, ALR2_out_21_port, ALR2_out_20_port, 
      ALR2_out_19_port, ALR2_out_18_port, ALR2_out_17_port, ALR2_out_16_port, 
      ALR2_out_15_port, ALR2_out_14_port, ALR2_out_13_port, ALR2_out_12_port, 
      ALR2_out_11_port, ALR2_out_10_port, ALR2_out_9_port, ALR2_out_8_port, 
      ALR2_out_7_port, ALR2_out_6_port, ALR2_out_5_port, ALR2_out_4_port, 
      ALR2_out_3_port, ALR2_out_2_port, ALR2_out_1_port, ALR2_out_0_port, 
      RWB3_out_20_port, RWB3_out_19_port, RWB3_out_18_port, RWB3_out_17_port, 
      RWB3_out_16_port, RWB3_out_15_port, RWB3_out_14_port, RWB3_out_13_port, 
      RWB3_out_12_port, RWB3_out_11_port, IMM_out_31_port, IMM_out_30_port, 
      IMM_out_29_port, IMM_out_28_port, IMM_out_27_port, IMM_out_26_port, 
      IMM_out_25_port, IMM_out_24_port, IMM_out_23_port, IMM_out_22_port, 
      IMM_out_21_port, IMM_out_20_port, IMM_out_19_port, IMM_out_18_port, 
      IMM_out_17_port, IMM_out_16_port, IMM_out_15_port, IMM_out_14_port, 
      IMM_out_13_port, IMM_out_12_port, IMM_out_11_port, IMM_out_10_port, 
      IMM_out_9_port, IMM_out_8_port, IMM_out_7_port, IMM_out_6_port, 
      IMM_out_5_port, IMM_out_4_port, IMM_out_3_port, IMM_out_2_port, 
      IMM_out_1_port, IMM_out_0_port, PC_SEL_1_port, PC_MUX_out_31_port, 
      PC_MUX_out_30_port, PC_MUX_out_29_port, PC_MUX_out_28_port, 
      PC_MUX_out_27_port, PC_MUX_out_26_port, PC_MUX_out_25_port, 
      PC_MUX_out_24_port, PC_MUX_out_23_port, PC_MUX_out_22_port, 
      PC_MUX_out_21_port, PC_MUX_out_20_port, PC_MUX_out_19_port, 
      PC_MUX_out_18_port, PC_MUX_out_17_port, PC_MUX_out_16_port, 
      PC_MUX_out_15_port, PC_MUX_out_14_port, PC_MUX_out_13_port, 
      PC_MUX_out_12_port, PC_MUX_out_11_port, PC_MUX_out_10_port, 
      PC_MUX_out_9_port, PC_MUX_out_8_port, PC_MUX_out_7_port, 
      PC_MUX_out_6_port, PC_MUX_out_5_port, PC_MUX_out_4_port, 
      PC_MUX_out_3_port, PC_MUX_out_2_port, PC_MUX_out_1_port, 
      PC_MUX_out_0_port, IRAMMUX_SEL, BHT_in_31_port, BHT_in_30_port, 
      BHT_in_29_port, BHT_in_28_port, BHT_in_27_port, BHT_in_26_port, 
      BHT_in_25_port, BHT_in_24_port, BHT_in_23_port, BHT_in_22_port, 
      BHT_in_21_port, BHT_in_20_port, BHT_in_19_port, BHT_in_18_port, 
      BHT_in_17_port, BHT_in_16_port, BHT_in_15_port, BHT_in_14_port, 
      BHT_in_13_port, BHT_in_12_port, BHT_in_11_port, BHT_in_10_port, 
      BHT_in_9_port, BHT_in_8_port, BHT_in_7_port, BHT_in_6_port, BHT_in_5_port
      , BHT_in_4_port, BHT_in_3_port, BHT_in_2_port, BHT_in_1_port, 
      BHT_in_0_port, FWDA_OUT_31_port, FWDA_OUT_30_port, FWDA_OUT_29_port, 
      FWDA_OUT_28_port, FWDA_OUT_27_port, FWDA_OUT_26_port, FWDA_OUT_25_port, 
      FWDA_OUT_24_port, FWDA_OUT_23_port, FWDA_OUT_22_port, FWDA_OUT_21_port, 
      FWDA_OUT_20_port, FWDA_OUT_19_port, FWDA_OUT_18_port, FWDA_OUT_17_port, 
      FWDA_OUT_16_port, FWDA_OUT_15_port, FWDA_OUT_14_port, FWDA_OUT_13_port, 
      FWDA_OUT_12_port, FWDA_OUT_11_port, FWDA_OUT_10_port, FWDA_OUT_9_port, 
      FWDA_OUT_8_port, FWDA_OUT_7_port, FWDA_OUT_6_port, FWDA_OUT_5_port, 
      FWDA_OUT_4_port, FWDA_OUT_3_port, FWDA_OUT_2_port, FWDA_OUT_1_port, 
      FWDA_OUT_0_port, A_in_31_port, A_in_30_port, A_in_29_port, A_in_28_port, 
      A_in_27_port, A_in_26_port, A_in_25_port, A_in_24_port, A_in_23_port, 
      A_in_22_port, A_in_21_port, A_in_20_port, A_in_19_port, A_in_18_port, 
      A_in_17_port, A_in_16_port, A_in_15_port, A_in_14_port, A_in_13_port, 
      A_in_12_port, A_in_11_port, A_in_10_port, A_in_9_port, A_in_8_port, 
      A_in_7_port, A_in_6_port, A_in_5_port, A_in_4_port, A_in_3_port, 
      A_in_2_port, A_in_1_port, A_in_0_port, FWDB_OUT_31_port, FWDB_OUT_30_port
      , FWDB_OUT_29_port, FWDB_OUT_28_port, FWDB_OUT_27_port, FWDB_OUT_26_port,
      FWDB_OUT_25_port, FWDB_OUT_24_port, FWDB_OUT_23_port, FWDB_OUT_22_port, 
      FWDB_OUT_21_port, FWDB_OUT_20_port, FWDB_OUT_19_port, FWDB_OUT_18_port, 
      FWDB_OUT_17_port, FWDB_OUT_16_port, FWDB_OUT_15_port, FWDB_OUT_14_port, 
      FWDB_OUT_13_port, FWDB_OUT_12_port, FWDB_OUT_11_port, FWDB_OUT_10_port, 
      FWDB_OUT_9_port, FWDB_OUT_8_port, FWDB_OUT_7_port, FWDB_OUT_6_port, 
      FWDB_OUT_5_port, FWDB_OUT_4_port, FWDB_OUT_3_port, FWDB_OUT_2_port, 
      FWDB_OUT_1_port, FWDB_OUT_0_port, B_in_31_port, B_in_30_port, 
      B_in_29_port, B_in_28_port, B_in_27_port, B_in_26_port, B_in_25_port, 
      B_in_24_port, B_in_23_port, B_in_22_port, B_in_21_port, B_in_20_port, 
      B_in_19_port, B_in_18_port, B_in_17_port, B_in_16_port, B_in_15_port, 
      B_in_14_port, B_in_13_port, B_in_12_port, B_in_11_port, B_in_10_port, 
      B_in_9_port, B_in_8_port, B_in_7_port, B_in_6_port, B_in_5_port, 
      B_in_4_port, B_in_3_port, B_in_2_port, B_in_1_port, B_in_0_port, 
      RA_out_31_port, RA_out_30_port, RA_out_29_port, RA_out_28_port, 
      RA_out_27_port, RA_out_26_port, RA_out_25_port, RA_out_24_port, 
      RA_out_23_port, RA_out_22_port, RA_out_21_port, RA_out_20_port, 
      RA_out_19_port, RA_out_18_port, RA_out_17_port, RA_out_16_port, 
      RA_out_15_port, RA_out_14_port, RA_out_13_port, RA_out_12_port, 
      RA_out_11_port, RA_out_10_port, RA_out_9_port, RA_out_8_port, 
      RA_out_7_port, RA_out_6_port, RA_out_5_port, RA_out_4_port, RA_out_3_port
      , RA_out_2_port, RA_out_1_port, RA_out_0_port, WB_in_31_port, 
      WB_in_30_port, WB_in_29_port, WB_in_28_port, WB_in_27_port, WB_in_26_port
      , WB_in_25_port, WB_in_24_port, WB_in_23_port, WB_in_22_port, 
      WB_in_21_port, WB_in_20_port, WB_in_19_port, WB_in_18_port, WB_in_17_port
      , WB_in_16_port, WB_in_15_port, WB_in_14_port, WB_in_13_port, 
      WB_in_12_port, WB_in_11_port, WB_in_10_port, WB_in_9_port, WB_in_8_port, 
      WB_in_7_port, WB_in_6_port, WB_in_5_port, WB_in_4_port, WB_in_3_port, 
      WB_in_2_port, WB_in_1_port, WB_in_0_port, FWDA_SEL_1_port, 
      FWDA_SEL_0_port, FWDB_SEL_1_port, FWDB_SEL_0_port, CWB_MUX2_out_31_port, 
      CWB_MUX2_out_30_port, CWB_MUX2_out_29_port, CWB_MUX2_out_28_port, 
      CWB_MUX2_out_27_port, CWB_MUX2_out_26_port, CWB_MUX2_out_25_port, 
      CWB_MUX2_out_24_port, CWB_MUX2_out_23_port, CWB_MUX2_out_22_port, 
      CWB_MUX2_out_21_port, CWB_MUX2_out_20_port, CWB_MUX2_out_19_port, 
      CWB_MUX2_out_18_port, CWB_MUX2_out_17_port, CWB_MUX2_out_16_port, 
      CWB_MUX2_out_15_port, CWB_MUX2_out_14_port, CWB_MUX2_out_13_port, 
      CWB_MUX2_out_12_port, CWB_MUX2_out_11_port, CWB_MUX2_out_10_port, 
      CWB_MUX2_out_9_port, CWB_MUX2_out_8_port, CWB_MUX2_out_7_port, 
      CWB_MUX2_out_6_port, CWB_MUX2_out_5_port, CWB_MUX2_out_4_port, 
      CWB_MUX2_out_3_port, CWB_MUX2_out_2_port, CWB_MUX2_out_1_port, 
      CWB_MUX2_out_0_port, ZDU_SEL_1_port, ZDU_SEL_0_port, ZDU_MUX_out_30_port,
      ZDU_MUX_out_29_port, ZDU_MUX_out_28_port, ZDU_MUX_out_27_port, 
      ZDU_MUX_out_26_port, ZDU_MUX_out_25_port, ZDU_MUX_out_24_port, 
      ZDU_MUX_out_23_port, ZDU_MUX_out_22_port, ZDU_MUX_out_21_port, 
      ZDU_MUX_out_20_port, ZDU_MUX_out_19_port, ZDU_MUX_out_18_port, 
      ZDU_MUX_out_17_port, ZDU_MUX_out_16_port, ZDU_MUX_out_15_port, 
      ZDU_MUX_out_14_port, ZDU_MUX_out_13_port, ZDU_MUX_out_12_port, 
      ZDU_MUX_out_11_port, ZDU_MUX_out_10_port, ZDU_MUX_out_9_port, 
      ZDU_MUX_out_8_port, ZDU_MUX_out_7_port, ZDU_MUX_out_6_port, 
      ZDU_MUX_out_5_port, ZDU_MUX_out_4_port, ZDU_MUX_out_3_port, 
      ZDU_MUX_out_2_port, ZDU_MUX_out_1_port, ZDU_MUX_out_0_port, 
      B2_MUX_out_31_port, B2_MUX_out_30_port, B2_MUX_out_29_port, 
      B2_MUX_out_28_port, B2_MUX_out_27_port, B2_MUX_out_26_port, 
      B2_MUX_out_25_port, B2_MUX_out_24_port, B2_MUX_out_23_port, 
      B2_MUX_out_22_port, B2_MUX_out_21_port, B2_MUX_out_20_port, 
      B2_MUX_out_19_port, B2_MUX_out_18_port, B2_MUX_out_17_port, 
      B2_MUX_out_16_port, B2_MUX_out_15_port, B2_MUX_out_14_port, 
      B2_MUX_out_13_port, B2_MUX_out_12_port, B2_MUX_out_11_port, 
      B2_MUX_out_10_port, B2_MUX_out_9_port, B2_MUX_out_8_port, 
      B2_MUX_out_7_port, B2_MUX_out_6_port, B2_MUX_out_5_port, 
      B2_MUX_out_4_port, B2_MUX_out_3_port, B2_MUX_out_2_port, 
      B2_MUX_out_1_port, B2_MUX_out_0_port, LMD_out_31_port, LMD_out_30_port, 
      LMD_out_29_port, LMD_out_28_port, LMD_out_27_port, LMD_out_26_port, 
      LMD_out_25_port, LMD_out_24_port, LMD_out_23_port, LMD_out_22_port, 
      LMD_out_21_port, LMD_out_20_port, LMD_out_19_port, LMD_out_18_port, 
      LMD_out_17_port, LMD_out_16_port, LMD_out_15_port, LMD_out_14_port, 
      LMD_out_13_port, LMD_out_12_port, LMD_out_11_port, LMD_out_10_port, 
      LMD_out_9_port, LMD_out_8_port, LMD_out_7_port, LMD_out_6_port, 
      LMD_out_5_port, LMD_out_4_port, LMD_out_3_port, LMD_out_2_port, 
      LMD_out_1_port, LMD_out_0_port, CWB_out_1_port, CWB_out_0_port, 
      CWB_MUX_SEL_1_port, CWB_MUX_SEL_0_port, CWB2_SEL_1_port, CWB2_SEL_0_port,
      FWDB2_SEL, RF_MUX_out_4_port, RF_MUX_out_3_port, RF_MUX_out_2_port, 
      RF_MUX_out_1_port, RF_MUX_out_0_port, IF_STALL, ID_STALL, EX_STALL, 
      MEM_STALL, ZDU_out, N14, n13, n14_port, n15, n16, n17, n18, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n25,
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792 : std_logic;

begin
   IRAM_ADDR <= ( IRAM_ADDR_31_port, IRAM_ADDR_30_port, IRAM_ADDR_29_port, 
      IRAM_ADDR_28_port, IRAM_ADDR_27_port, IRAM_ADDR_26_port, 
      IRAM_ADDR_25_port, IRAM_ADDR_24_port, IRAM_ADDR_23_port, 
      IRAM_ADDR_22_port, IRAM_ADDR_21_port, IRAM_ADDR_20_port, 
      IRAM_ADDR_19_port, IRAM_ADDR_18_port, IRAM_ADDR_17_port, 
      IRAM_ADDR_16_port, IRAM_ADDR_15_port, IRAM_ADDR_14_port, 
      IRAM_ADDR_13_port, IRAM_ADDR_12_port, IRAM_ADDR_11_port, 
      IRAM_ADDR_10_port, IRAM_ADDR_9_port, IRAM_ADDR_8_port, IRAM_ADDR_7_port, 
      IRAM_ADDR_6_port, IRAM_ADDR_5_port, IRAM_ADDR_4_port, IRAM_ADDR_3_port, 
      IRAM_ADDR_2_port, IRAM_ADDR_1_port, IRAM_ADDR_0_port );
   DATA_ADDR <= ( DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RegPC : REG_NBIT32_0 port map( clk => CLK, reset => n23, enable => n33, 
                           data_in(31) => NPC_in_31_port, data_in(30) => 
                           NPC_in_30_port, data_in(29) => NPC_in_29_port, 
                           data_in(28) => NPC_in_28_port, data_in(27) => 
                           NPC_in_27_port, data_in(26) => NPC_in_26_port, 
                           data_in(25) => NPC_in_25_port, data_in(24) => 
                           NPC_in_24_port, data_in(23) => NPC_in_23_port, 
                           data_in(22) => NPC_in_22_port, data_in(21) => 
                           NPC_in_21_port, data_in(20) => NPC_in_20_port, 
                           data_in(19) => NPC_in_19_port, data_in(18) => 
                           NPC_in_18_port, data_in(17) => NPC_in_17_port, 
                           data_in(16) => NPC_in_16_port, data_in(15) => 
                           NPC_in_15_port, data_in(14) => NPC_in_14_port, 
                           data_in(13) => NPC_in_13_port, data_in(12) => 
                           NPC_in_12_port, data_in(11) => NPC_in_11_port, 
                           data_in(10) => NPC_in_10_port, data_in(9) => 
                           NPC_in_9_port, data_in(8) => NPC_in_8_port, 
                           data_in(7) => NPC_in_7_port, data_in(6) => 
                           NPC_in_6_port, data_in(5) => NPC_in_5_port, 
                           data_in(4) => NPC_in_4_port, data_in(3) => 
                           NPC_in_3_port, data_in(2) => NPC_in_2_port, 
                           data_in(1) => NPC_in_1_port, data_in(0) => 
                           NPC_in_0_port, data_out(31) => PC_out_31_port, 
                           data_out(30) => PC_out_30_port, data_out(29) => 
                           PC_out_29_port, data_out(28) => PC_out_28_port, 
                           data_out(27) => PC_out_27_port, data_out(26) => 
                           PC_out_26_port, data_out(25) => PC_out_25_port, 
                           data_out(24) => PC_out_24_port, data_out(23) => 
                           PC_out_23_port, data_out(22) => PC_out_22_port, 
                           data_out(21) => PC_out_21_port, data_out(20) => 
                           PC_out_20_port, data_out(19) => PC_out_19_port, 
                           data_out(18) => PC_out_18_port, data_out(17) => 
                           PC_out_17_port, data_out(16) => PC_out_16_port, 
                           data_out(15) => PC_out_15_port, data_out(14) => 
                           PC_out_14_port, data_out(13) => PC_out_13_port, 
                           data_out(12) => PC_out_12_port, data_out(11) => 
                           PC_out_11_port, data_out(10) => PC_out_10_port, 
                           data_out(9) => PC_out_9_port, data_out(8) => 
                           PC_out_8_port, data_out(7) => PC_out_7_port, 
                           data_out(6) => PC_out_6_port, data_out(5) => 
                           PC_out_5_port, data_out(4) => PC_out_4_port, 
                           data_out(3) => PC_out_3_port, data_out(2) => 
                           PC_out_2_port, data_out(1) => PC_out_1_port, 
                           data_out(0) => PC_out_0_port);
   RegIR : REG_NBIT32_17 port map( clk => CLK, reset => n24, enable => n33, 
                           data_in(31) => IRAM_OUT(31), data_in(30) => 
                           IRAM_OUT(30), data_in(29) => IRAM_OUT(29), 
                           data_in(28) => IRAM_OUT(28), data_in(27) => 
                           IRAM_OUT(27), data_in(26) => IRAM_OUT(26), 
                           data_in(25) => IRAM_OUT(25), data_in(24) => 
                           IRAM_OUT(24), data_in(23) => IRAM_OUT(23), 
                           data_in(22) => IRAM_OUT(22), data_in(21) => 
                           IRAM_OUT(21), data_in(20) => IRAM_OUT(20), 
                           data_in(19) => IRAM_OUT(19), data_in(18) => 
                           IRAM_OUT(18), data_in(17) => IRAM_OUT(17), 
                           data_in(16) => IRAM_OUT(16), data_in(15) => 
                           IRAM_OUT(15), data_in(14) => IRAM_OUT(14), 
                           data_in(13) => IRAM_OUT(13), data_in(12) => 
                           IRAM_OUT(12), data_in(11) => IRAM_OUT(11), 
                           data_in(10) => IRAM_OUT(10), data_in(9) => 
                           IRAM_OUT(9), data_in(8) => IRAM_OUT(8), data_in(7) 
                           => IRAM_OUT(7), data_in(6) => IRAM_OUT(6), 
                           data_in(5) => IRAM_OUT(5), data_in(4) => IRAM_OUT(4)
                           , data_in(3) => IRAM_OUT(3), data_in(2) => 
                           IRAM_OUT(2), data_in(1) => IRAM_OUT(1), data_in(0) 
                           => IRAM_OUT(0), data_out(31) => IR_out_31_port, 
                           data_out(30) => IR_out_30_port, data_out(29) => 
                           IR_out_29_port, data_out(28) => IR_out_28_port, 
                           data_out(27) => IR_out_27_port, data_out(26) => 
                           IR_out_26_port, data_out(25) => IR_out_25_port, 
                           data_out(24) => IR_out_24_port, data_out(23) => 
                           IR_out_23_port, data_out(22) => IR_out_22_port, 
                           data_out(21) => IR_out_21_port, data_out(20) => 
                           IR_out_20_port, data_out(19) => IR_out_19_port, 
                           data_out(18) => IR_out_18_port, data_out(17) => 
                           IR_out_17_port, data_out(16) => IR_out_16_port, 
                           data_out(15) => IR_out_15_port, data_out(14) => 
                           IR_out_14_port, data_out(13) => IR_out_13_port, 
                           data_out(12) => IR_out_12_port, data_out(11) => 
                           IR_out_11_port, data_out(10) => IR_out_10_port, 
                           data_out(9) => IR_out_9_port, data_out(8) => 
                           IR_out_8_port, data_out(7) => IR_out_7_port, 
                           data_out(6) => IR_out_6_port, data_out(5) => 
                           IR_out_5_port, data_out(4) => IR_out_4_port, 
                           data_out(3) => IR_out_3_port, data_out(2) => 
                           IR_out_2_port, data_out(1) => IR_out_1_port, 
                           data_out(0) => IR_out_0_port);
   RegNPC : REG_NBIT32_16 port map( clk => CLK, reset => n24, enable => n33, 
                           data_in(31) => NPC_in_31_port, data_in(30) => 
                           NPC_in_30_port, data_in(29) => NPC_in_29_port, 
                           data_in(28) => NPC_in_28_port, data_in(27) => 
                           NPC_in_27_port, data_in(26) => NPC_in_26_port, 
                           data_in(25) => NPC_in_25_port, data_in(24) => 
                           NPC_in_24_port, data_in(23) => NPC_in_23_port, 
                           data_in(22) => NPC_in_22_port, data_in(21) => 
                           NPC_in_21_port, data_in(20) => NPC_in_20_port, 
                           data_in(19) => NPC_in_19_port, data_in(18) => 
                           NPC_in_18_port, data_in(17) => NPC_in_17_port, 
                           data_in(16) => NPC_in_16_port, data_in(15) => 
                           NPC_in_15_port, data_in(14) => NPC_in_14_port, 
                           data_in(13) => NPC_in_13_port, data_in(12) => 
                           NPC_in_12_port, data_in(11) => NPC_in_11_port, 
                           data_in(10) => NPC_in_10_port, data_in(9) => 
                           NPC_in_9_port, data_in(8) => NPC_in_8_port, 
                           data_in(7) => NPC_in_7_port, data_in(6) => 
                           NPC_in_6_port, data_in(5) => NPC_in_5_port, 
                           data_in(4) => NPC_in_4_port, data_in(3) => 
                           NPC_in_3_port, data_in(2) => NPC_in_2_port, 
                           data_in(1) => NPC_in_1_port, data_in(0) => 
                           NPC_in_0_port, data_out(31) => NPC_out_31_port, 
                           data_out(30) => NPC_out_30_port, data_out(29) => 
                           NPC_out_29_port, data_out(28) => NPC_out_28_port, 
                           data_out(27) => NPC_out_27_port, data_out(26) => 
                           NPC_out_26_port, data_out(25) => NPC_out_25_port, 
                           data_out(24) => NPC_out_24_port, data_out(23) => 
                           NPC_out_23_port, data_out(22) => NPC_out_22_port, 
                           data_out(21) => NPC_out_21_port, data_out(20) => 
                           NPC_out_20_port, data_out(19) => NPC_out_19_port, 
                           data_out(18) => NPC_out_18_port, data_out(17) => 
                           NPC_out_17_port, data_out(16) => NPC_out_16_port, 
                           data_out(15) => NPC_out_15_port, data_out(14) => 
                           NPC_out_14_port, data_out(13) => NPC_out_13_port, 
                           data_out(12) => NPC_out_12_port, data_out(11) => 
                           NPC_out_11_port, data_out(10) => NPC_out_10_port, 
                           data_out(9) => NPC_out_9_port, data_out(8) => 
                           NPC_out_8_port, data_out(7) => NPC_out_7_port, 
                           data_out(6) => NPC_out_6_port, data_out(5) => 
                           NPC_out_5_port, data_out(4) => NPC_out_4_port, 
                           data_out(3) => NPC_out_3_port, data_out(2) => 
                           NPC_out_2_port, data_out(1) => NPC_out_1_port, 
                           data_out(0) => NPC_out_0_port);
   RegPC2 : REG_NBIT32_15 port map( clk => CLK, reset => n24, enable => n1, 
                           data_in(31) => PC_out_31_port, data_in(30) => 
                           PC_out_30_port, data_in(29) => PC_out_29_port, 
                           data_in(28) => PC_out_28_port, data_in(27) => 
                           PC_out_27_port, data_in(26) => PC_out_26_port, 
                           data_in(25) => PC_out_25_port, data_in(24) => 
                           PC_out_24_port, data_in(23) => PC_out_23_port, 
                           data_in(22) => PC_out_22_port, data_in(21) => 
                           PC_out_21_port, data_in(20) => PC_out_20_port, 
                           data_in(19) => PC_out_19_port, data_in(18) => 
                           PC_out_18_port, data_in(17) => PC_out_17_port, 
                           data_in(16) => PC_out_16_port, data_in(15) => 
                           PC_out_15_port, data_in(14) => PC_out_14_port, 
                           data_in(13) => PC_out_13_port, data_in(12) => 
                           PC_out_12_port, data_in(11) => PC_out_11_port, 
                           data_in(10) => PC_out_10_port, data_in(9) => 
                           PC_out_9_port, data_in(8) => PC_out_8_port, 
                           data_in(7) => PC_out_7_port, data_in(6) => 
                           PC_out_6_port, data_in(5) => PC_out_5_port, 
                           data_in(4) => PC_out_4_port, data_in(3) => 
                           PC_out_3_port, data_in(2) => PC_out_2_port, 
                           data_in(1) => PC_out_1_port, data_in(0) => 
                           PC_out_0_port, data_out(31) => PC2_out_31_port, 
                           data_out(30) => PC2_out_30_port, data_out(29) => 
                           PC2_out_29_port, data_out(28) => PC2_out_28_port, 
                           data_out(27) => PC2_out_27_port, data_out(26) => 
                           PC2_out_26_port, data_out(25) => PC2_out_25_port, 
                           data_out(24) => PC2_out_24_port, data_out(23) => 
                           PC2_out_23_port, data_out(22) => PC2_out_22_port, 
                           data_out(21) => PC2_out_21_port, data_out(20) => 
                           PC2_out_20_port, data_out(19) => PC2_out_19_port, 
                           data_out(18) => PC2_out_18_port, data_out(17) => 
                           PC2_out_17_port, data_out(16) => PC2_out_16_port, 
                           data_out(15) => PC2_out_15_port, data_out(14) => 
                           PC2_out_14_port, data_out(13) => PC2_out_13_port, 
                           data_out(12) => PC2_out_12_port, data_out(11) => 
                           PC2_out_11_port, data_out(10) => PC2_out_10_port, 
                           data_out(9) => PC2_out_9_port, data_out(8) => 
                           PC2_out_8_port, data_out(7) => PC2_out_7_port, 
                           data_out(6) => PC2_out_6_port, data_out(5) => 
                           PC2_out_5_port, data_out(4) => PC2_out_4_port, 
                           data_out(3) => PC2_out_3_port, data_out(2) => 
                           PC2_out_2_port, data_out(1) => PC2_out_1_port, 
                           data_out(0) => PC2_out_0_port);
   RegIMM : REG_NBIT32_14 port map( clk => CLK, reset => n24, enable => n1, 
                           data_in(31) => N14, data_in(30) => N14, data_in(29) 
                           => N14, data_in(28) => N14, data_in(27) => N14, 
                           data_in(26) => N14, data_in(25) => N14, data_in(24) 
                           => N14, data_in(23) => N14, data_in(22) => N14, 
                           data_in(21) => N14, data_in(20) => N14, data_in(19) 
                           => N14, data_in(18) => N14, data_in(17) => N14, 
                           data_in(16) => N14, data_in(15) => IR_out_15_port, 
                           data_in(14) => IR_out_14_port, data_in(13) => 
                           IR_out_13_port, data_in(12) => IR_out_12_port, 
                           data_in(11) => IR_out_11_port, data_in(10) => 
                           IR_out_10_port, data_in(9) => IR_out_9_port, 
                           data_in(8) => IR_out_8_port, data_in(7) => 
                           IR_out_7_port, data_in(6) => IR_out_6_port, 
                           data_in(5) => IR_out_5_port, data_in(4) => 
                           IR_out_4_port, data_in(3) => IR_out_3_port, 
                           data_in(2) => IR_out_2_port, data_in(1) => 
                           IR_out_1_port, data_in(0) => IR_out_0_port, 
                           data_out(31) => RIMM_out_31_port, data_out(30) => 
                           RIMM_out_30_port, data_out(29) => RIMM_out_29_port, 
                           data_out(28) => RIMM_out_28_port, data_out(27) => 
                           RIMM_out_27_port, data_out(26) => RIMM_out_26_port, 
                           data_out(25) => RIMM_out_25_port, data_out(24) => 
                           RIMM_out_24_port, data_out(23) => RIMM_out_23_port, 
                           data_out(22) => RIMM_out_22_port, data_out(21) => 
                           RIMM_out_21_port, data_out(20) => RIMM_out_20_port, 
                           data_out(19) => RIMM_out_19_port, data_out(18) => 
                           RIMM_out_18_port, data_out(17) => RIMM_out_17_port, 
                           data_out(16) => RIMM_out_16_port, data_out(15) => 
                           RIMM_out_15_port, data_out(14) => RIMM_out_14_port, 
                           data_out(13) => RIMM_out_13_port, data_out(12) => 
                           RIMM_out_12_port, data_out(11) => RIMM_out_11_port, 
                           data_out(10) => RIMM_out_10_port, data_out(9) => 
                           RIMM_out_9_port, data_out(8) => RIMM_out_8_port, 
                           data_out(7) => RIMM_out_7_port, data_out(6) => 
                           RIMM_out_6_port, data_out(5) => RIMM_out_5_port, 
                           data_out(4) => RIMM_out_4_port, data_out(3) => 
                           RIMM_out_3_port, data_out(2) => RIMM_out_2_port, 
                           data_out(1) => RIMM_out_1_port, data_out(0) => 
                           RIMM_out_0_port);
   RegWB1 : REG_NBIT32_13 port map( clk => CLK, reset => n24, enable => n1, 
                           data_in(31) => IR_out_31_port, data_in(30) => 
                           IR_out_30_port, data_in(29) => IR_out_29_port, 
                           data_in(28) => IR_out_28_port, data_in(27) => 
                           IR_out_27_port, data_in(26) => IR_out_26_port, 
                           data_in(25) => IR_out_25_port, data_in(24) => 
                           IR_out_24_port, data_in(23) => IR_out_23_port, 
                           data_in(22) => IR_out_22_port, data_in(21) => 
                           IR_out_21_port, data_in(20) => IR_out_20_port, 
                           data_in(19) => IR_out_19_port, data_in(18) => 
                           IR_out_18_port, data_in(17) => IR_out_17_port, 
                           data_in(16) => IR_out_16_port, data_in(15) => 
                           IR_out_15_port, data_in(14) => IR_out_14_port, 
                           data_in(13) => IR_out_13_port, data_in(12) => 
                           IR_out_12_port, data_in(11) => IR_out_11_port, 
                           data_in(10) => IR_out_10_port, data_in(9) => 
                           IR_out_9_port, data_in(8) => IR_out_8_port, 
                           data_in(7) => IR_out_7_port, data_in(6) => 
                           IR_out_6_port, data_in(5) => IR_out_5_port, 
                           data_in(4) => IR_out_4_port, data_in(3) => 
                           IR_out_3_port, data_in(2) => IR_out_2_port, 
                           data_in(1) => IR_out_1_port, data_in(0) => 
                           IR_out_0_port, data_out(31) => RWB1_out_31_port, 
                           data_out(30) => RWB1_out_30_port, data_out(29) => 
                           RWB1_out_29_port, data_out(28) => RWB1_out_28_port, 
                           data_out(27) => RWB1_out_27_port, data_out(26) => 
                           RWB1_out_26_port, data_out(25) => RWB1_out_25_port, 
                           data_out(24) => RWB1_out_24_port, data_out(23) => 
                           RWB1_out_23_port, data_out(22) => RWB1_out_22_port, 
                           data_out(21) => RWB1_out_21_port, data_out(20) => 
                           RWB1_out_20_port, data_out(19) => RWB1_out_19_port, 
                           data_out(18) => RWB1_out_18_port, data_out(17) => 
                           RWB1_out_17_port, data_out(16) => RWB1_out_16_port, 
                           data_out(15) => RWB1_out_15_port, data_out(14) => 
                           RWB1_out_14_port, data_out(13) => RWB1_out_13_port, 
                           data_out(12) => RWB1_out_12_port, data_out(11) => 
                           RWB1_out_11_port, data_out(10) => RWB1_out_10_port, 
                           data_out(9) => RWB1_out_9_port, data_out(8) => 
                           RWB1_out_8_port, data_out(7) => RWB1_out_7_port, 
                           data_out(6) => RWB1_out_6_port, data_out(5) => 
                           RWB1_out_5_port, data_out(4) => RWB1_out_4_port, 
                           data_out(3) => RWB1_out_3_port, data_out(2) => 
                           RWB1_out_2_port, data_out(1) => RWB1_out_1_port, 
                           data_out(0) => RWB1_out_0_port);
   F_PRD : FFD_0 port map( D => BHT_out, CK => CLK, RESET => n23, ENABLE => n1,
                           Q => PRD_OUT);
   RegNPC2 : REG_NBIT32_12 port map( clk => CLK, reset => n24, enable => n1, 
                           data_in(31) => NPC_out_31_port, data_in(30) => 
                           NPC_out_30_port, data_in(29) => NPC_out_29_port, 
                           data_in(28) => NPC_out_28_port, data_in(27) => 
                           NPC_out_27_port, data_in(26) => NPC_out_26_port, 
                           data_in(25) => NPC_out_25_port, data_in(24) => 
                           NPC_out_24_port, data_in(23) => NPC_out_23_port, 
                           data_in(22) => NPC_out_22_port, data_in(21) => 
                           NPC_out_21_port, data_in(20) => NPC_out_20_port, 
                           data_in(19) => NPC_out_19_port, data_in(18) => 
                           NPC_out_18_port, data_in(17) => NPC_out_17_port, 
                           data_in(16) => NPC_out_16_port, data_in(15) => 
                           NPC_out_15_port, data_in(14) => NPC_out_14_port, 
                           data_in(13) => NPC_out_13_port, data_in(12) => 
                           NPC_out_12_port, data_in(11) => NPC_out_11_port, 
                           data_in(10) => NPC_out_10_port, data_in(9) => 
                           NPC_out_9_port, data_in(8) => NPC_out_8_port, 
                           data_in(7) => NPC_out_7_port, data_in(6) => 
                           NPC_out_6_port, data_in(5) => NPC_out_5_port, 
                           data_in(4) => NPC_out_4_port, data_in(3) => 
                           NPC_out_3_port, data_in(2) => NPC_out_2_port, 
                           data_in(1) => NPC_out_1_port, data_in(0) => 
                           NPC_out_0_port, data_out(31) => NPC2_out_31_port, 
                           data_out(30) => NPC2_out_30_port, data_out(29) => 
                           NPC2_out_29_port, data_out(28) => NPC2_out_28_port, 
                           data_out(27) => NPC2_out_27_port, data_out(26) => 
                           NPC2_out_26_port, data_out(25) => NPC2_out_25_port, 
                           data_out(24) => NPC2_out_24_port, data_out(23) => 
                           NPC2_out_23_port, data_out(22) => NPC2_out_22_port, 
                           data_out(21) => NPC2_out_21_port, data_out(20) => 
                           NPC2_out_20_port, data_out(19) => NPC2_out_19_port, 
                           data_out(18) => NPC2_out_18_port, data_out(17) => 
                           NPC2_out_17_port, data_out(16) => NPC2_out_16_port, 
                           data_out(15) => NPC2_out_15_port, data_out(14) => 
                           NPC2_out_14_port, data_out(13) => NPC2_out_13_port, 
                           data_out(12) => NPC2_out_12_port, data_out(11) => 
                           NPC2_out_11_port, data_out(10) => NPC2_out_10_port, 
                           data_out(9) => NPC2_out_9_port, data_out(8) => 
                           NPC2_out_8_port, data_out(7) => NPC2_out_7_port, 
                           data_out(6) => NPC2_out_6_port, data_out(5) => 
                           NPC2_out_5_port, data_out(4) => NPC2_out_4_port, 
                           data_out(3) => NPC2_out_3_port, data_out(2) => 
                           NPC2_out_2_port, data_out(1) => NPC2_out_1_port, 
                           data_out(0) => NPC2_out_0_port);
   RegJADD2 : REG_NBIT32_11 port map( clk => CLK, reset => n24, enable => n1, 
                           data_in(31) => JADDER_out_31_port, data_in(30) => 
                           JADDER_out_30_port, data_in(29) => 
                           JADDER_out_29_port, data_in(28) => 
                           JADDER_out_28_port, data_in(27) => 
                           JADDER_out_27_port, data_in(26) => 
                           JADDER_out_26_port, data_in(25) => 
                           JADDER_out_25_port, data_in(24) => 
                           JADDER_out_24_port, data_in(23) => 
                           JADDER_out_23_port, data_in(22) => 
                           JADDER_out_22_port, data_in(21) => 
                           JADDER_out_21_port, data_in(20) => 
                           JADDER_out_20_port, data_in(19) => 
                           JADDER_out_19_port, data_in(18) => 
                           JADDER_out_18_port, data_in(17) => 
                           JADDER_out_17_port, data_in(16) => 
                           JADDER_out_16_port, data_in(15) => 
                           JADDER_out_15_port, data_in(14) => 
                           JADDER_out_14_port, data_in(13) => 
                           JADDER_out_13_port, data_in(12) => 
                           JADDER_out_12_port, data_in(11) => 
                           JADDER_out_11_port, data_in(10) => 
                           JADDER_out_10_port, data_in(9) => JADDER_out_9_port,
                           data_in(8) => JADDER_out_8_port, data_in(7) => 
                           JADDER_out_7_port, data_in(6) => JADDER_out_6_port, 
                           data_in(5) => JADDER_out_5_port, data_in(4) => 
                           JADDER_out_4_port, data_in(3) => JADDER_out_3_port, 
                           data_in(2) => JADDER_out_2_port, data_in(1) => 
                           JADDER_out_1_port, data_in(0) => JADDER_out_0_port, 
                           data_out(31) => JADDER2_out_31_port, data_out(30) =>
                           JADDER2_out_30_port, data_out(29) => 
                           JADDER2_out_29_port, data_out(28) => 
                           JADDER2_out_28_port, data_out(27) => 
                           JADDER2_out_27_port, data_out(26) => 
                           JADDER2_out_26_port, data_out(25) => 
                           JADDER2_out_25_port, data_out(24) => 
                           JADDER2_out_24_port, data_out(23) => 
                           JADDER2_out_23_port, data_out(22) => 
                           JADDER2_out_22_port, data_out(21) => 
                           JADDER2_out_21_port, data_out(20) => 
                           JADDER2_out_20_port, data_out(19) => 
                           JADDER2_out_19_port, data_out(18) => 
                           JADDER2_out_18_port, data_out(17) => 
                           JADDER2_out_17_port, data_out(16) => 
                           JADDER2_out_16_port, data_out(15) => 
                           JADDER2_out_15_port, data_out(14) => 
                           JADDER2_out_14_port, data_out(13) => 
                           JADDER2_out_13_port, data_out(12) => 
                           JADDER2_out_12_port, data_out(11) => 
                           JADDER2_out_11_port, data_out(10) => 
                           JADDER2_out_10_port, data_out(9) => 
                           JADDER2_out_9_port, data_out(8) => 
                           JADDER2_out_8_port, data_out(7) => 
                           JADDER2_out_7_port, data_out(6) => 
                           JADDER2_out_6_port, data_out(5) => 
                           JADDER2_out_5_port, data_out(4) => 
                           JADDER2_out_4_port, data_out(3) => 
                           JADDER2_out_3_port, data_out(2) => 
                           JADDER2_out_2_port, data_out(1) => 
                           JADDER2_out_1_port, data_out(0) => 
                           JADDER2_out_0_port);
   F_JR : FFD_1 port map( D => BPR_EN, CK => CLK, RESET => n23, ENABLE => n1, Q
                           => BPR_EN2);
   RegPC3 : REG_NBIT32_10 port map( clk => CLK, reset => n24, enable => n6, 
                           data_in(31) => PC2_out_31_port, data_in(30) => 
                           PC2_out_30_port, data_in(29) => PC2_out_29_port, 
                           data_in(28) => PC2_out_28_port, data_in(27) => 
                           PC2_out_27_port, data_in(26) => PC2_out_26_port, 
                           data_in(25) => PC2_out_25_port, data_in(24) => 
                           PC2_out_24_port, data_in(23) => PC2_out_23_port, 
                           data_in(22) => PC2_out_22_port, data_in(21) => 
                           PC2_out_21_port, data_in(20) => PC2_out_20_port, 
                           data_in(19) => PC2_out_19_port, data_in(18) => 
                           PC2_out_18_port, data_in(17) => PC2_out_17_port, 
                           data_in(16) => PC2_out_16_port, data_in(15) => 
                           PC2_out_15_port, data_in(14) => PC2_out_14_port, 
                           data_in(13) => PC2_out_13_port, data_in(12) => 
                           PC2_out_12_port, data_in(11) => PC2_out_11_port, 
                           data_in(10) => PC2_out_10_port, data_in(9) => 
                           PC2_out_9_port, data_in(8) => PC2_out_8_port, 
                           data_in(7) => PC2_out_7_port, data_in(6) => 
                           PC2_out_6_port, data_in(5) => PC2_out_5_port, 
                           data_in(4) => PC2_out_4_port, data_in(3) => 
                           PC2_out_3_port, data_in(2) => PC2_out_2_port, 
                           data_in(1) => PC2_out_1_port, data_in(0) => 
                           PC2_out_0_port, data_out(31) => PC3_out_31_port, 
                           data_out(30) => PC3_out_30_port, data_out(29) => 
                           PC3_out_29_port, data_out(28) => PC3_out_28_port, 
                           data_out(27) => PC3_out_27_port, data_out(26) => 
                           PC3_out_26_port, data_out(25) => PC3_out_25_port, 
                           data_out(24) => PC3_out_24_port, data_out(23) => 
                           PC3_out_23_port, data_out(22) => PC3_out_22_port, 
                           data_out(21) => PC3_out_21_port, data_out(20) => 
                           PC3_out_20_port, data_out(19) => PC3_out_19_port, 
                           data_out(18) => PC3_out_18_port, data_out(17) => 
                           PC3_out_17_port, data_out(16) => PC3_out_16_port, 
                           data_out(15) => PC3_out_15_port, data_out(14) => 
                           PC3_out_14_port, data_out(13) => PC3_out_13_port, 
                           data_out(12) => PC3_out_12_port, data_out(11) => 
                           PC3_out_11_port, data_out(10) => PC3_out_10_port, 
                           data_out(9) => PC3_out_9_port, data_out(8) => 
                           PC3_out_8_port, data_out(7) => PC3_out_7_port, 
                           data_out(6) => PC3_out_6_port, data_out(5) => 
                           PC3_out_5_port, data_out(4) => PC3_out_4_port, 
                           data_out(3) => PC3_out_3_port, data_out(2) => 
                           PC3_out_2_port, data_out(1) => PC3_out_1_port, 
                           data_out(0) => PC3_out_0_port);
   RegWB2 : REG_NBIT32_9 port map( clk => CLK, reset => n23, enable => n6, 
                           data_in(31) => RWB1_out_31_port, data_in(30) => 
                           RWB1_out_30_port, data_in(29) => RWB1_out_29_port, 
                           data_in(28) => RWB1_out_28_port, data_in(27) => 
                           RWB1_out_27_port, data_in(26) => RWB1_out_26_port, 
                           data_in(25) => RWB1_out_25_port, data_in(24) => 
                           RWB1_out_24_port, data_in(23) => RWB1_out_23_port, 
                           data_in(22) => RWB1_out_22_port, data_in(21) => 
                           RWB1_out_21_port, data_in(20) => RWB1_out_20_port, 
                           data_in(19) => RWB1_out_19_port, data_in(18) => 
                           RWB1_out_18_port, data_in(17) => RWB1_out_17_port, 
                           data_in(16) => RWB1_out_16_port, data_in(15) => 
                           RWB1_out_15_port, data_in(14) => RWB1_out_14_port, 
                           data_in(13) => RWB1_out_13_port, data_in(12) => 
                           RWB1_out_12_port, data_in(11) => RWB1_out_11_port, 
                           data_in(10) => RWB1_out_10_port, data_in(9) => 
                           RWB1_out_9_port, data_in(8) => RWB1_out_8_port, 
                           data_in(7) => RWB1_out_7_port, data_in(6) => 
                           RWB1_out_6_port, data_in(5) => RWB1_out_5_port, 
                           data_in(4) => RWB1_out_4_port, data_in(3) => 
                           RWB1_out_3_port, data_in(2) => RWB1_out_2_port, 
                           data_in(1) => RWB1_out_1_port, data_in(0) => 
                           RWB1_out_0_port, data_out(31) => RWB2_out_31_port, 
                           data_out(30) => RWB2_out_30_port, data_out(29) => 
                           RWB2_out_29_port, data_out(28) => RWB2_out_28_port, 
                           data_out(27) => RWB2_out_27_port, data_out(26) => 
                           RWB2_out_26_port, data_out(25) => RWB2_out_25_port, 
                           data_out(24) => RWB2_out_24_port, data_out(23) => 
                           RWB2_out_23_port, data_out(22) => RWB2_out_22_port, 
                           data_out(21) => RWB2_out_21_port, data_out(20) => 
                           RWB2_out_20_port, data_out(19) => RWB2_out_19_port, 
                           data_out(18) => RWB2_out_18_port, data_out(17) => 
                           RWB2_out_17_port, data_out(16) => RWB2_out_16_port, 
                           data_out(15) => RWB2_out_15_port, data_out(14) => 
                           RWB2_out_14_port, data_out(13) => RWB2_out_13_port, 
                           data_out(12) => RWB2_out_12_port, data_out(11) => 
                           RWB2_out_11_port, data_out(10) => RWB2_out_10_port, 
                           data_out(9) => RWB2_out_9_port, data_out(8) => 
                           RWB2_out_8_port, data_out(7) => RWB2_out_7_port, 
                           data_out(6) => RWB2_out_6_port, data_out(5) => 
                           RWB2_out_5_port, data_out(4) => RWB2_out_4_port, 
                           data_out(3) => RWB2_out_3_port, data_out(2) => 
                           RWB2_out_2_port, data_out(1) => RWB2_out_1_port, 
                           data_out(0) => RWB2_out_0_port);
   RegB2 : REG_NBIT32_8 port map( clk => CLK, reset => n23, enable => n6, 
                           data_in(31) => RB_out_31_port, data_in(30) => 
                           RB_out_30_port, data_in(29) => RB_out_29_port, 
                           data_in(28) => RB_out_28_port, data_in(27) => 
                           RB_out_27_port, data_in(26) => RB_out_26_port, 
                           data_in(25) => RB_out_25_port, data_in(24) => 
                           RB_out_24_port, data_in(23) => RB_out_23_port, 
                           data_in(22) => RB_out_22_port, data_in(21) => 
                           RB_out_21_port, data_in(20) => RB_out_20_port, 
                           data_in(19) => RB_out_19_port, data_in(18) => 
                           RB_out_18_port, data_in(17) => RB_out_17_port, 
                           data_in(16) => RB_out_16_port, data_in(15) => 
                           RB_out_15_port, data_in(14) => RB_out_14_port, 
                           data_in(13) => RB_out_13_port, data_in(12) => 
                           RB_out_12_port, data_in(11) => RB_out_11_port, 
                           data_in(10) => RB_out_10_port, data_in(9) => 
                           RB_out_9_port, data_in(8) => RB_out_8_port, 
                           data_in(7) => RB_out_7_port, data_in(6) => 
                           RB_out_6_port, data_in(5) => RB_out_5_port, 
                           data_in(4) => RB_out_4_port, data_in(3) => 
                           RB_out_3_port, data_in(2) => RB_out_2_port, 
                           data_in(1) => RB_out_1_port, data_in(0) => 
                           RB_out_0_port, data_out(31) => B2_out_31_port, 
                           data_out(30) => B2_out_30_port, data_out(29) => 
                           B2_out_29_port, data_out(28) => B2_out_28_port, 
                           data_out(27) => B2_out_27_port, data_out(26) => 
                           B2_out_26_port, data_out(25) => B2_out_25_port, 
                           data_out(24) => B2_out_24_port, data_out(23) => 
                           B2_out_23_port, data_out(22) => B2_out_22_port, 
                           data_out(21) => B2_out_21_port, data_out(20) => 
                           B2_out_20_port, data_out(19) => B2_out_19_port, 
                           data_out(18) => B2_out_18_port, data_out(17) => 
                           B2_out_17_port, data_out(16) => B2_out_16_port, 
                           data_out(15) => B2_out_15_port, data_out(14) => 
                           B2_out_14_port, data_out(13) => B2_out_13_port, 
                           data_out(12) => B2_out_12_port, data_out(11) => 
                           B2_out_11_port, data_out(10) => B2_out_10_port, 
                           data_out(9) => B2_out_9_port, data_out(8) => 
                           B2_out_8_port, data_out(7) => B2_out_7_port, 
                           data_out(6) => B2_out_6_port, data_out(5) => 
                           B2_out_5_port, data_out(4) => B2_out_4_port, 
                           data_out(3) => B2_out_3_port, data_out(2) => 
                           B2_out_2_port, data_out(1) => B2_out_1_port, 
                           data_out(0) => B2_out_0_port);
   RegALR : REG_NBIT32_7 port map( clk => CLK, reset => n23, enable => n6, 
                           data_in(31) => ALR_in_31_port, data_in(30) => 
                           ALR_in_30_port, data_in(29) => ALR_in_29_port, 
                           data_in(28) => ALR_in_28_port, data_in(27) => 
                           ALR_in_27_port, data_in(26) => ALR_in_26_port, 
                           data_in(25) => ALR_in_25_port, data_in(24) => 
                           ALR_in_24_port, data_in(23) => ALR_in_23_port, 
                           data_in(22) => ALR_in_22_port, data_in(21) => 
                           ALR_in_21_port, data_in(20) => ALR_in_20_port, 
                           data_in(19) => ALR_in_19_port, data_in(18) => 
                           ALR_in_18_port, data_in(17) => ALR_in_17_port, 
                           data_in(16) => ALR_in_16_port, data_in(15) => 
                           ALR_in_15_port, data_in(14) => ALR_in_14_port, 
                           data_in(13) => ALR_in_13_port, data_in(12) => 
                           ALR_in_12_port, data_in(11) => ALR_in_11_port, 
                           data_in(10) => ALR_in_10_port, data_in(9) => 
                           ALR_in_9_port, data_in(8) => ALR_in_8_port, 
                           data_in(7) => ALR_in_7_port, data_in(6) => 
                           ALR_in_6_port, data_in(5) => ALR_in_5_port, 
                           data_in(4) => ALR_in_4_port, data_in(3) => 
                           ALR_in_3_port, data_in(2) => ALR_in_2_port, 
                           data_in(1) => ALR_in_1_port, data_in(0) => 
                           ALR_in_0_port, data_out(31) => DATA_ADDR_31_port, 
                           data_out(30) => DATA_ADDR_30_port, data_out(29) => 
                           DATA_ADDR_29_port, data_out(28) => DATA_ADDR_28_port
                           , data_out(27) => DATA_ADDR_27_port, data_out(26) =>
                           DATA_ADDR_26_port, data_out(25) => DATA_ADDR_25_port
                           , data_out(24) => DATA_ADDR_24_port, data_out(23) =>
                           DATA_ADDR_23_port, data_out(22) => DATA_ADDR_22_port
                           , data_out(21) => DATA_ADDR_21_port, data_out(20) =>
                           DATA_ADDR_20_port, data_out(19) => DATA_ADDR_19_port
                           , data_out(18) => DATA_ADDR_18_port, data_out(17) =>
                           DATA_ADDR_17_port, data_out(16) => DATA_ADDR_16_port
                           , data_out(15) => DATA_ADDR_15_port, data_out(14) =>
                           DATA_ADDR_14_port, data_out(13) => DATA_ADDR_13_port
                           , data_out(12) => DATA_ADDR_12_port, data_out(11) =>
                           DATA_ADDR_11_port, data_out(10) => DATA_ADDR_10_port
                           , data_out(9) => DATA_ADDR_9_port, data_out(8) => 
                           DATA_ADDR_8_port, data_out(7) => DATA_ADDR_7_port, 
                           data_out(6) => DATA_ADDR_6_port, data_out(5) => 
                           DATA_ADDR_5_port, data_out(4) => DATA_ADDR_4_port, 
                           data_out(3) => DATA_ADDR_3_port, data_out(2) => 
                           DATA_ADDR_2_port, data_out(1) => DATA_ADDR_1_port, 
                           data_out(0) => DATA_ADDR_0_port);
   RegNPC3 : REG_NBIT32_6 port map( clk => CLK, reset => n23, enable => n6, 
                           data_in(31) => NPC2_out_31_port, data_in(30) => 
                           NPC2_out_30_port, data_in(29) => NPC2_out_29_port, 
                           data_in(28) => NPC2_out_28_port, data_in(27) => 
                           NPC2_out_27_port, data_in(26) => NPC2_out_26_port, 
                           data_in(25) => NPC2_out_25_port, data_in(24) => 
                           NPC2_out_24_port, data_in(23) => NPC2_out_23_port, 
                           data_in(22) => NPC2_out_22_port, data_in(21) => 
                           NPC2_out_21_port, data_in(20) => NPC2_out_20_port, 
                           data_in(19) => NPC2_out_19_port, data_in(18) => 
                           NPC2_out_18_port, data_in(17) => NPC2_out_17_port, 
                           data_in(16) => NPC2_out_16_port, data_in(15) => 
                           NPC2_out_15_port, data_in(14) => NPC2_out_14_port, 
                           data_in(13) => NPC2_out_13_port, data_in(12) => 
                           NPC2_out_12_port, data_in(11) => NPC2_out_11_port, 
                           data_in(10) => NPC2_out_10_port, data_in(9) => 
                           NPC2_out_9_port, data_in(8) => NPC2_out_8_port, 
                           data_in(7) => NPC2_out_7_port, data_in(6) => 
                           NPC2_out_6_port, data_in(5) => NPC2_out_5_port, 
                           data_in(4) => NPC2_out_4_port, data_in(3) => 
                           NPC2_out_3_port, data_in(2) => NPC2_out_2_port, 
                           data_in(1) => NPC2_out_1_port, data_in(0) => 
                           NPC2_out_0_port, data_out(31) => NPC3_out_31_port, 
                           data_out(30) => NPC3_out_30_port, data_out(29) => 
                           NPC3_out_29_port, data_out(28) => NPC3_out_28_port, 
                           data_out(27) => NPC3_out_27_port, data_out(26) => 
                           NPC3_out_26_port, data_out(25) => NPC3_out_25_port, 
                           data_out(24) => NPC3_out_24_port, data_out(23) => 
                           NPC3_out_23_port, data_out(22) => NPC3_out_22_port, 
                           data_out(21) => NPC3_out_21_port, data_out(20) => 
                           NPC3_out_20_port, data_out(19) => NPC3_out_19_port, 
                           data_out(18) => NPC3_out_18_port, data_out(17) => 
                           NPC3_out_17_port, data_out(16) => NPC3_out_16_port, 
                           data_out(15) => NPC3_out_15_port, data_out(14) => 
                           NPC3_out_14_port, data_out(13) => NPC3_out_13_port, 
                           data_out(12) => NPC3_out_12_port, data_out(11) => 
                           NPC3_out_11_port, data_out(10) => NPC3_out_10_port, 
                           data_out(9) => NPC3_out_9_port, data_out(8) => 
                           NPC3_out_8_port, data_out(7) => NPC3_out_7_port, 
                           data_out(6) => NPC3_out_6_port, data_out(5) => 
                           NPC3_out_5_port, data_out(4) => NPC3_out_4_port, 
                           data_out(3) => NPC3_out_3_port, data_out(2) => 
                           NPC3_out_2_port, data_out(1) => NPC3_out_1_port, 
                           data_out(0) => NPC3_out_0_port);
   RegPSW : REG_NBIT7 port map( clk => CLK, reset => n23, enable => n6, 
                           data_in(6) => PSW_in_6_port, data_in(5) => 
                           PSW_in_5_port, data_in(4) => PSW_in_4_port, 
                           data_in(3) => PSW_in_3_port, data_in(2) => 
                           PSW_in_2_port, data_in(1) => PSW_in_1_port, 
                           data_in(0) => PSW_in_0_port, data_out(6) => 
                           PSW_out_6_port, data_out(5) => PSW_out_5_port, 
                           data_out(4) => PSW_out_4_port, data_out(3) => 
                           PSW_out_3_port, data_out(2) => PSW_out_2_port, 
                           data_out(1) => PSW_out_1_port, data_out(0) => 
                           PSW_out_0_port);
   RegALR2 : REG_NBIT32_5 port map( clk => CLK, reset => n23, enable => n5, 
                           data_in(31) => ALR2_in_31_port, data_in(30) => 
                           ALR2_in_30_port, data_in(29) => ALR2_in_29_port, 
                           data_in(28) => ALR2_in_28_port, data_in(27) => 
                           ALR2_in_27_port, data_in(26) => ALR2_in_26_port, 
                           data_in(25) => ALR2_in_25_port, data_in(24) => 
                           ALR2_in_24_port, data_in(23) => ALR2_in_23_port, 
                           data_in(22) => ALR2_in_22_port, data_in(21) => 
                           ALR2_in_21_port, data_in(20) => ALR2_in_20_port, 
                           data_in(19) => ALR2_in_19_port, data_in(18) => 
                           ALR2_in_18_port, data_in(17) => ALR2_in_17_port, 
                           data_in(16) => ALR2_in_16_port, data_in(15) => 
                           ALR2_in_15_port, data_in(14) => ALR2_in_14_port, 
                           data_in(13) => ALR2_in_13_port, data_in(12) => 
                           ALR2_in_12_port, data_in(11) => ALR2_in_11_port, 
                           data_in(10) => ALR2_in_10_port, data_in(9) => 
                           ALR2_in_9_port, data_in(8) => ALR2_in_8_port, 
                           data_in(7) => ALR2_in_7_port, data_in(6) => 
                           ALR2_in_6_port, data_in(5) => ALR2_in_5_port, 
                           data_in(4) => ALR2_in_4_port, data_in(3) => 
                           ALR2_in_3_port, data_in(2) => ALR2_in_2_port, 
                           data_in(1) => ALR2_in_1_port, data_in(0) => 
                           ALR2_in_0_port, data_out(31) => ALR2_out_31_port, 
                           data_out(30) => ALR2_out_30_port, data_out(29) => 
                           ALR2_out_29_port, data_out(28) => ALR2_out_28_port, 
                           data_out(27) => ALR2_out_27_port, data_out(26) => 
                           ALR2_out_26_port, data_out(25) => ALR2_out_25_port, 
                           data_out(24) => ALR2_out_24_port, data_out(23) => 
                           ALR2_out_23_port, data_out(22) => ALR2_out_22_port, 
                           data_out(21) => ALR2_out_21_port, data_out(20) => 
                           ALR2_out_20_port, data_out(19) => ALR2_out_19_port, 
                           data_out(18) => ALR2_out_18_port, data_out(17) => 
                           ALR2_out_17_port, data_out(16) => ALR2_out_16_port, 
                           data_out(15) => ALR2_out_15_port, data_out(14) => 
                           ALR2_out_14_port, data_out(13) => ALR2_out_13_port, 
                           data_out(12) => ALR2_out_12_port, data_out(11) => 
                           ALR2_out_11_port, data_out(10) => ALR2_out_10_port, 
                           data_out(9) => ALR2_out_9_port, data_out(8) => 
                           ALR2_out_8_port, data_out(7) => ALR2_out_7_port, 
                           data_out(6) => ALR2_out_6_port, data_out(5) => 
                           ALR2_out_5_port, data_out(4) => ALR2_out_4_port, 
                           data_out(3) => ALR2_out_3_port, data_out(2) => 
                           ALR2_out_2_port, data_out(1) => ALR2_out_1_port, 
                           data_out(0) => ALR2_out_0_port);
   RegWB3 : REG_NBIT32_4 port map( clk => CLK, reset => n23, enable => n5, 
                           data_in(31) => RWB2_out_31_port, data_in(30) => 
                           RWB2_out_30_port, data_in(29) => RWB2_out_29_port, 
                           data_in(28) => RWB2_out_28_port, data_in(27) => 
                           RWB2_out_27_port, data_in(26) => RWB2_out_26_port, 
                           data_in(25) => RWB2_out_25_port, data_in(24) => 
                           RWB2_out_24_port, data_in(23) => RWB2_out_23_port, 
                           data_in(22) => RWB2_out_22_port, data_in(21) => 
                           RWB2_out_21_port, data_in(20) => RWB2_out_20_port, 
                           data_in(19) => RWB2_out_19_port, data_in(18) => 
                           RWB2_out_18_port, data_in(17) => RWB2_out_17_port, 
                           data_in(16) => RWB2_out_16_port, data_in(15) => 
                           RWB2_out_15_port, data_in(14) => RWB2_out_14_port, 
                           data_in(13) => RWB2_out_13_port, data_in(12) => 
                           RWB2_out_12_port, data_in(11) => RWB2_out_11_port, 
                           data_in(10) => RWB2_out_10_port, data_in(9) => 
                           RWB2_out_9_port, data_in(8) => RWB2_out_8_port, 
                           data_in(7) => RWB2_out_7_port, data_in(6) => 
                           RWB2_out_6_port, data_in(5) => RWB2_out_5_port, 
                           data_in(4) => RWB2_out_4_port, data_in(3) => 
                           RWB2_out_3_port, data_in(2) => RWB2_out_2_port, 
                           data_in(1) => RWB2_out_1_port, data_in(0) => 
                           RWB2_out_0_port, data_out(31) => n_1769, 
                           data_out(30) => n_1770, data_out(29) => n_1771, 
                           data_out(28) => n_1772, data_out(27) => n_1773, 
                           data_out(26) => n_1774, data_out(25) => n_1775, 
                           data_out(24) => n_1776, data_out(23) => n_1777, 
                           data_out(22) => n_1778, data_out(21) => n_1779, 
                           data_out(20) => RWB3_out_20_port, data_out(19) => 
                           RWB3_out_19_port, data_out(18) => RWB3_out_18_port, 
                           data_out(17) => RWB3_out_17_port, data_out(16) => 
                           RWB3_out_16_port, data_out(15) => RWB3_out_15_port, 
                           data_out(14) => RWB3_out_14_port, data_out(13) => 
                           RWB3_out_13_port, data_out(12) => RWB3_out_12_port, 
                           data_out(11) => RWB3_out_11_port, data_out(10) => 
                           n_1780, data_out(9) => n_1781, data_out(8) => n_1782
                           , data_out(7) => n_1783, data_out(6) => n_1784, 
                           data_out(5) => n_1785, data_out(4) => n_1786, 
                           data_out(3) => n_1787, data_out(2) => n_1788, 
                           data_out(1) => n_1789, data_out(0) => n_1790);
   AdderPC : PC_adder_0 port map( A(31) => IRAM_ADDR_31_port, A(30) => 
                           IRAM_ADDR_30_port, A(29) => IRAM_ADDR_29_port, A(28)
                           => IRAM_ADDR_28_port, A(27) => IRAM_ADDR_27_port, 
                           A(26) => IRAM_ADDR_26_port, A(25) => 
                           IRAM_ADDR_25_port, A(24) => IRAM_ADDR_24_port, A(23)
                           => IRAM_ADDR_23_port, A(22) => IRAM_ADDR_22_port, 
                           A(21) => IRAM_ADDR_21_port, A(20) => 
                           IRAM_ADDR_20_port, A(19) => IRAM_ADDR_19_port, A(18)
                           => IRAM_ADDR_18_port, A(17) => IRAM_ADDR_17_port, 
                           A(16) => IRAM_ADDR_16_port, A(15) => 
                           IRAM_ADDR_15_port, A(14) => IRAM_ADDR_14_port, A(13)
                           => IRAM_ADDR_13_port, A(12) => IRAM_ADDR_12_port, 
                           A(11) => IRAM_ADDR_11_port, A(10) => 
                           IRAM_ADDR_10_port, A(9) => IRAM_ADDR_9_port, A(8) =>
                           IRAM_ADDR_8_port, A(7) => IRAM_ADDR_7_port, A(6) => 
                           IRAM_ADDR_6_port, A(5) => IRAM_ADDR_5_port, A(4) => 
                           IRAM_ADDR_4_port, A(3) => IRAM_ADDR_3_port, A(2) => 
                           IRAM_ADDR_2_port, A(1) => IRAM_ADDR_1_port, A(0) => 
                           IRAM_ADDR_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, Sum(31) => NPC_in_31_port, Sum(30) =>
                           NPC_in_30_port, Sum(29) => NPC_in_29_port, Sum(28) 
                           => NPC_in_28_port, Sum(27) => NPC_in_27_port, 
                           Sum(26) => NPC_in_26_port, Sum(25) => NPC_in_25_port
                           , Sum(24) => NPC_in_24_port, Sum(23) => 
                           NPC_in_23_port, Sum(22) => NPC_in_22_port, Sum(21) 
                           => NPC_in_21_port, Sum(20) => NPC_in_20_port, 
                           Sum(19) => NPC_in_19_port, Sum(18) => NPC_in_18_port
                           , Sum(17) => NPC_in_17_port, Sum(16) => 
                           NPC_in_16_port, Sum(15) => NPC_in_15_port, Sum(14) 
                           => NPC_in_14_port, Sum(13) => NPC_in_13_port, 
                           Sum(12) => NPC_in_12_port, Sum(11) => NPC_in_11_port
                           , Sum(10) => NPC_in_10_port, Sum(9) => NPC_in_9_port
                           , Sum(8) => NPC_in_8_port, Sum(7) => NPC_in_7_port, 
                           Sum(6) => NPC_in_6_port, Sum(5) => NPC_in_5_port, 
                           Sum(4) => NPC_in_4_port, Sum(3) => NPC_in_3_port, 
                           Sum(2) => NPC_in_2_port, Sum(1) => NPC_in_1_port, 
                           Sum(0) => NPC_in_0_port);
   J_Adder : PC_adder_1 port map( A(31) => PC2_out_31_port, A(30) => 
                           PC2_out_30_port, A(29) => PC2_out_29_port, A(28) => 
                           PC2_out_28_port, A(27) => PC2_out_27_port, A(26) => 
                           PC2_out_26_port, A(25) => PC2_out_25_port, A(24) => 
                           PC2_out_24_port, A(23) => PC2_out_23_port, A(22) => 
                           PC2_out_22_port, A(21) => PC2_out_21_port, A(20) => 
                           PC2_out_20_port, A(19) => PC2_out_19_port, A(18) => 
                           PC2_out_18_port, A(17) => PC2_out_17_port, A(16) => 
                           PC2_out_16_port, A(15) => PC2_out_15_port, A(14) => 
                           PC2_out_14_port, A(13) => PC2_out_13_port, A(12) => 
                           PC2_out_12_port, A(11) => PC2_out_11_port, A(10) => 
                           PC2_out_10_port, A(9) => PC2_out_9_port, A(8) => 
                           PC2_out_8_port, A(7) => PC2_out_7_port, A(6) => 
                           PC2_out_6_port, A(5) => PC2_out_5_port, A(4) => 
                           PC2_out_4_port, A(3) => PC2_out_3_port, A(2) => 
                           PC2_out_2_port, A(1) => PC2_out_1_port, A(0) => 
                           PC2_out_0_port, B(31) => IMM_out_31_port, B(30) => 
                           IMM_out_30_port, B(29) => IMM_out_29_port, B(28) => 
                           IMM_out_28_port, B(27) => IMM_out_27_port, B(26) => 
                           IMM_out_26_port, B(25) => IMM_out_25_port, B(24) => 
                           IMM_out_24_port, B(23) => IMM_out_23_port, B(22) => 
                           IMM_out_22_port, B(21) => IMM_out_21_port, B(20) => 
                           IMM_out_20_port, B(19) => IMM_out_19_port, B(18) => 
                           IMM_out_18_port, B(17) => IMM_out_17_port, B(16) => 
                           IMM_out_16_port, B(15) => IMM_out_15_port, B(14) => 
                           IMM_out_14_port, B(13) => IMM_out_13_port, B(12) => 
                           IMM_out_12_port, B(11) => IMM_out_11_port, B(10) => 
                           IMM_out_10_port, B(9) => IMM_out_9_port, B(8) => 
                           IMM_out_8_port, B(7) => IMM_out_7_port, B(6) => 
                           IMM_out_6_port, B(5) => IMM_out_5_port, B(4) => 
                           IMM_out_4_port, B(3) => IMM_out_3_port, B(2) => 
                           IMM_out_2_port, B(1) => IMM_out_1_port, B(0) => 
                           IMM_out_0_port, Sum(31) => JADDER_out_31_port, 
                           Sum(30) => JADDER_out_30_port, Sum(29) => 
                           JADDER_out_29_port, Sum(28) => JADDER_out_28_port, 
                           Sum(27) => JADDER_out_27_port, Sum(26) => 
                           JADDER_out_26_port, Sum(25) => JADDER_out_25_port, 
                           Sum(24) => JADDER_out_24_port, Sum(23) => 
                           JADDER_out_23_port, Sum(22) => JADDER_out_22_port, 
                           Sum(21) => JADDER_out_21_port, Sum(20) => 
                           JADDER_out_20_port, Sum(19) => JADDER_out_19_port, 
                           Sum(18) => JADDER_out_18_port, Sum(17) => 
                           JADDER_out_17_port, Sum(16) => JADDER_out_16_port, 
                           Sum(15) => JADDER_out_15_port, Sum(14) => 
                           JADDER_out_14_port, Sum(13) => JADDER_out_13_port, 
                           Sum(12) => JADDER_out_12_port, Sum(11) => 
                           JADDER_out_11_port, Sum(10) => JADDER_out_10_port, 
                           Sum(9) => JADDER_out_9_port, Sum(8) => 
                           JADDER_out_8_port, Sum(7) => JADDER_out_7_port, 
                           Sum(6) => JADDER_out_6_port, Sum(5) => 
                           JADDER_out_5_port, Sum(4) => JADDER_out_4_port, 
                           Sum(3) => JADDER_out_3_port, Sum(2) => 
                           JADDER_out_2_port, Sum(1) => JADDER_out_1_port, 
                           Sum(0) => JADDER_out_0_port);
   PCMUX : MUX3to1_NBIT32_0 port map( A(31) => PC_out_31_port, A(30) => 
                           PC_out_30_port, A(29) => PC_out_29_port, A(28) => 
                           PC_out_28_port, A(27) => PC_out_27_port, A(26) => 
                           PC_out_26_port, A(25) => PC_out_25_port, A(24) => 
                           PC_out_24_port, A(23) => PC_out_23_port, A(22) => 
                           PC_out_22_port, A(21) => PC_out_21_port, A(20) => 
                           PC_out_20_port, A(19) => PC_out_19_port, A(18) => 
                           PC_out_18_port, A(17) => PC_out_17_port, A(16) => 
                           PC_out_16_port, A(15) => PC_out_15_port, A(14) => 
                           PC_out_14_port, A(13) => PC_out_13_port, A(12) => 
                           PC_out_12_port, A(11) => PC_out_11_port, A(10) => 
                           PC_out_10_port, A(9) => PC_out_9_port, A(8) => 
                           PC_out_8_port, A(7) => PC_out_7_port, A(6) => 
                           PC_out_6_port, A(5) => PC_out_5_port, A(4) => 
                           PC_out_4_port, A(3) => PC_out_3_port, A(2) => 
                           PC_out_2_port, A(1) => PC_out_1_port, A(0) => 
                           PC_out_0_port, B(31) => JADDER_out_31_port, B(30) =>
                           JADDER_out_30_port, B(29) => JADDER_out_29_port, 
                           B(28) => JADDER_out_28_port, B(27) => 
                           JADDER_out_27_port, B(26) => JADDER_out_26_port, 
                           B(25) => JADDER_out_25_port, B(24) => 
                           JADDER_out_24_port, B(23) => JADDER_out_23_port, 
                           B(22) => JADDER_out_22_port, B(21) => 
                           JADDER_out_21_port, B(20) => JADDER_out_20_port, 
                           B(19) => JADDER_out_19_port, B(18) => 
                           JADDER_out_18_port, B(17) => JADDER_out_17_port, 
                           B(16) => JADDER_out_16_port, B(15) => 
                           JADDER_out_15_port, B(14) => JADDER_out_14_port, 
                           B(13) => JADDER_out_13_port, B(12) => 
                           JADDER_out_12_port, B(11) => JADDER_out_11_port, 
                           B(10) => JADDER_out_10_port, B(9) => 
                           JADDER_out_9_port, B(8) => JADDER_out_8_port, B(7) 
                           => JADDER_out_7_port, B(6) => JADDER_out_6_port, 
                           B(5) => JADDER_out_5_port, B(4) => JADDER_out_4_port
                           , B(3) => JADDER_out_3_port, B(2) => 
                           JADDER_out_2_port, B(1) => JADDER_out_1_port, B(0) 
                           => JADDER_out_0_port, C(31) => JADDER2_out_31_port, 
                           C(30) => JADDER2_out_30_port, C(29) => 
                           JADDER2_out_29_port, C(28) => JADDER2_out_28_port, 
                           C(27) => JADDER2_out_27_port, C(26) => 
                           JADDER2_out_26_port, C(25) => JADDER2_out_25_port, 
                           C(24) => JADDER2_out_24_port, C(23) => 
                           JADDER2_out_23_port, C(22) => JADDER2_out_22_port, 
                           C(21) => JADDER2_out_21_port, C(20) => 
                           JADDER2_out_20_port, C(19) => JADDER2_out_19_port, 
                           C(18) => JADDER2_out_18_port, C(17) => 
                           JADDER2_out_17_port, C(16) => JADDER2_out_16_port, 
                           C(15) => JADDER2_out_15_port, C(14) => 
                           JADDER2_out_14_port, C(13) => JADDER2_out_13_port, 
                           C(12) => JADDER2_out_12_port, C(11) => 
                           JADDER2_out_11_port, C(10) => JADDER2_out_10_port, 
                           C(9) => JADDER2_out_9_port, C(8) => 
                           JADDER2_out_8_port, C(7) => JADDER2_out_7_port, C(6)
                           => JADDER2_out_6_port, C(5) => JADDER2_out_5_port, 
                           C(4) => JADDER2_out_4_port, C(3) => 
                           JADDER2_out_3_port, C(2) => JADDER2_out_2_port, C(1)
                           => JADDER2_out_1_port, C(0) => JADDER2_out_0_port, 
                           SEL(1) => PC_SEL_1_port, SEL(0) => n34, Y(31) => 
                           PC_MUX_out_31_port, Y(30) => PC_MUX_out_30_port, 
                           Y(29) => PC_MUX_out_29_port, Y(28) => 
                           PC_MUX_out_28_port, Y(27) => PC_MUX_out_27_port, 
                           Y(26) => PC_MUX_out_26_port, Y(25) => 
                           PC_MUX_out_25_port, Y(24) => PC_MUX_out_24_port, 
                           Y(23) => PC_MUX_out_23_port, Y(22) => 
                           PC_MUX_out_22_port, Y(21) => PC_MUX_out_21_port, 
                           Y(20) => PC_MUX_out_20_port, Y(19) => 
                           PC_MUX_out_19_port, Y(18) => PC_MUX_out_18_port, 
                           Y(17) => PC_MUX_out_17_port, Y(16) => 
                           PC_MUX_out_16_port, Y(15) => PC_MUX_out_15_port, 
                           Y(14) => PC_MUX_out_14_port, Y(13) => 
                           PC_MUX_out_13_port, Y(12) => PC_MUX_out_12_port, 
                           Y(11) => PC_MUX_out_11_port, Y(10) => 
                           PC_MUX_out_10_port, Y(9) => PC_MUX_out_9_port, Y(8) 
                           => PC_MUX_out_8_port, Y(7) => PC_MUX_out_7_port, 
                           Y(6) => PC_MUX_out_6_port, Y(5) => PC_MUX_out_5_port
                           , Y(4) => PC_MUX_out_4_port, Y(3) => 
                           PC_MUX_out_3_port, Y(2) => PC_MUX_out_2_port, Y(1) 
                           => PC_MUX_out_1_port, Y(0) => PC_MUX_out_0_port);
   IRAMMUX : MUX2to1_NBIT32_0 port map( A(31) => PC_MUX_out_31_port, A(30) => 
                           PC_MUX_out_30_port, A(29) => PC_MUX_out_29_port, 
                           A(28) => PC_MUX_out_28_port, A(27) => 
                           PC_MUX_out_27_port, A(26) => PC_MUX_out_26_port, 
                           A(25) => PC_MUX_out_25_port, A(24) => 
                           PC_MUX_out_24_port, A(23) => PC_MUX_out_23_port, 
                           A(22) => PC_MUX_out_22_port, A(21) => 
                           PC_MUX_out_21_port, A(20) => PC_MUX_out_20_port, 
                           A(19) => PC_MUX_out_19_port, A(18) => 
                           PC_MUX_out_18_port, A(17) => PC_MUX_out_17_port, 
                           A(16) => PC_MUX_out_16_port, A(15) => 
                           PC_MUX_out_15_port, A(14) => PC_MUX_out_14_port, 
                           A(13) => PC_MUX_out_13_port, A(12) => 
                           PC_MUX_out_12_port, A(11) => PC_MUX_out_11_port, 
                           A(10) => PC_MUX_out_10_port, A(9) => 
                           PC_MUX_out_9_port, A(8) => PC_MUX_out_8_port, A(7) 
                           => PC_MUX_out_7_port, A(6) => PC_MUX_out_6_port, 
                           A(5) => PC_MUX_out_5_port, A(4) => PC_MUX_out_4_port
                           , A(3) => PC_MUX_out_3_port, A(2) => 
                           PC_MUX_out_2_port, A(1) => PC_MUX_out_1_port, A(0) 
                           => PC_MUX_out_0_port, B(31) => NPC2_out_31_port, 
                           B(30) => NPC2_out_30_port, B(29) => NPC2_out_29_port
                           , B(28) => NPC2_out_28_port, B(27) => 
                           NPC2_out_27_port, B(26) => NPC2_out_26_port, B(25) 
                           => NPC2_out_25_port, B(24) => NPC2_out_24_port, 
                           B(23) => NPC2_out_23_port, B(22) => NPC2_out_22_port
                           , B(21) => NPC2_out_21_port, B(20) => 
                           NPC2_out_20_port, B(19) => NPC2_out_19_port, B(18) 
                           => NPC2_out_18_port, B(17) => NPC2_out_17_port, 
                           B(16) => NPC2_out_16_port, B(15) => NPC2_out_15_port
                           , B(14) => NPC2_out_14_port, B(13) => 
                           NPC2_out_13_port, B(12) => NPC2_out_12_port, B(11) 
                           => NPC2_out_11_port, B(10) => NPC2_out_10_port, B(9)
                           => NPC2_out_9_port, B(8) => NPC2_out_8_port, B(7) =>
                           NPC2_out_7_port, B(6) => NPC2_out_6_port, B(5) => 
                           NPC2_out_5_port, B(4) => NPC2_out_4_port, B(3) => 
                           NPC2_out_3_port, B(2) => NPC2_out_2_port, B(1) => 
                           NPC2_out_1_port, B(0) => NPC2_out_0_port, SEL => 
                           IRAMMUX_SEL, Y(31) => IRAM_ADDR_31_port, Y(30) => 
                           IRAM_ADDR_30_port, Y(29) => IRAM_ADDR_29_port, Y(28)
                           => IRAM_ADDR_28_port, Y(27) => IRAM_ADDR_27_port, 
                           Y(26) => IRAM_ADDR_26_port, Y(25) => 
                           IRAM_ADDR_25_port, Y(24) => IRAM_ADDR_24_port, Y(23)
                           => IRAM_ADDR_23_port, Y(22) => IRAM_ADDR_22_port, 
                           Y(21) => IRAM_ADDR_21_port, Y(20) => 
                           IRAM_ADDR_20_port, Y(19) => IRAM_ADDR_19_port, Y(18)
                           => IRAM_ADDR_18_port, Y(17) => IRAM_ADDR_17_port, 
                           Y(16) => IRAM_ADDR_16_port, Y(15) => 
                           IRAM_ADDR_15_port, Y(14) => IRAM_ADDR_14_port, Y(13)
                           => IRAM_ADDR_13_port, Y(12) => IRAM_ADDR_12_port, 
                           Y(11) => IRAM_ADDR_11_port, Y(10) => 
                           IRAM_ADDR_10_port, Y(9) => IRAM_ADDR_9_port, Y(8) =>
                           IRAM_ADDR_8_port, Y(7) => IRAM_ADDR_7_port, Y(6) => 
                           IRAM_ADDR_6_port, Y(5) => IRAM_ADDR_5_port, Y(4) => 
                           IRAM_ADDR_4_port, Y(3) => IRAM_ADDR_3_port, Y(2) => 
                           IRAM_ADDR_2_port, Y(1) => IRAM_ADDR_1_port, Y(0) => 
                           IRAM_ADDR_0_port);
   IMMMUX : MUX2to1_NBIT32_8 port map( A(31) => IR_out_15_port, A(30) => 
                           IR_out_15_port, A(29) => IR_out_15_port, A(28) => 
                           IR_out_15_port, A(27) => IR_out_15_port, A(26) => 
                           IR_out_15_port, A(25) => IR_out_15_port, A(24) => 
                           IR_out_15_port, A(23) => IR_out_15_port, A(22) => 
                           IR_out_15_port, A(21) => IR_out_15_port, A(20) => 
                           IR_out_15_port, A(19) => IR_out_15_port, A(18) => 
                           IR_out_15_port, A(17) => IR_out_15_port, A(16) => 
                           IR_out_15_port, A(15) => IR_out_15_port, A(14) => 
                           IR_out_14_port, A(13) => IR_out_13_port, A(12) => 
                           IR_out_12_port, A(11) => IR_out_11_port, A(10) => 
                           IR_out_10_port, A(9) => IR_out_9_port, A(8) => 
                           IR_out_8_port, A(7) => IR_out_7_port, A(6) => 
                           IR_out_6_port, A(5) => IR_out_5_port, A(4) => 
                           IR_out_4_port, A(3) => IR_out_3_port, A(2) => 
                           IR_out_2_port, A(1) => IR_out_1_port, A(0) => 
                           IR_out_0_port, B(31) => IR_out_25_port, B(30) => 
                           IR_out_25_port, B(29) => IR_out_25_port, B(28) => 
                           IR_out_25_port, B(27) => IR_out_25_port, B(26) => 
                           IR_out_25_port, B(25) => IR_out_25_port, B(24) => 
                           IR_out_24_port, B(23) => IR_out_23_port, B(22) => 
                           IR_out_22_port, B(21) => IR_out_21_port, B(20) => 
                           IR_out_20_port, B(19) => IR_out_19_port, B(18) => 
                           IR_out_18_port, B(17) => IR_out_17_port, B(16) => 
                           IR_out_16_port, B(15) => IR_out_15_port, B(14) => 
                           IR_out_14_port, B(13) => IR_out_13_port, B(12) => 
                           IR_out_12_port, B(11) => IR_out_11_port, B(10) => 
                           IR_out_10_port, B(9) => IR_out_9_port, B(8) => 
                           IR_out_8_port, B(7) => IR_out_7_port, B(6) => 
                           IR_out_6_port, B(5) => IR_out_5_port, B(4) => 
                           IR_out_4_port, B(3) => IR_out_3_port, B(2) => 
                           IR_out_2_port, B(1) => IR_out_1_port, B(0) => 
                           IR_out_0_port, SEL => IMM_SEL, Y(31) => 
                           IMM_out_31_port, Y(30) => IMM_out_30_port, Y(29) => 
                           IMM_out_29_port, Y(28) => IMM_out_28_port, Y(27) => 
                           IMM_out_27_port, Y(26) => IMM_out_26_port, Y(25) => 
                           IMM_out_25_port, Y(24) => IMM_out_24_port, Y(23) => 
                           IMM_out_23_port, Y(22) => IMM_out_22_port, Y(21) => 
                           IMM_out_21_port, Y(20) => IMM_out_20_port, Y(19) => 
                           IMM_out_19_port, Y(18) => IMM_out_18_port, Y(17) => 
                           IMM_out_17_port, Y(16) => IMM_out_16_port, Y(15) => 
                           IMM_out_15_port, Y(14) => IMM_out_14_port, Y(13) => 
                           IMM_out_13_port, Y(12) => IMM_out_12_port, Y(11) => 
                           IMM_out_11_port, Y(10) => IMM_out_10_port, Y(9) => 
                           IMM_out_9_port, Y(8) => IMM_out_8_port, Y(7) => 
                           IMM_out_7_port, Y(6) => IMM_out_6_port, Y(5) => 
                           IMM_out_5_port, Y(4) => IMM_out_4_port, Y(3) => 
                           IMM_out_3_port, Y(2) => IMM_out_2_port, Y(1) => 
                           IMM_out_1_port, Y(0) => IMM_out_0_port);
   BHTMUX : MUX2to1_NBIT32_7 port map( A(31) => PC2_out_31_port, A(30) => 
                           PC2_out_30_port, A(29) => PC2_out_29_port, A(28) => 
                           PC2_out_28_port, A(27) => PC2_out_27_port, A(26) => 
                           PC2_out_26_port, A(25) => PC2_out_25_port, A(24) => 
                           PC2_out_24_port, A(23) => PC2_out_23_port, A(22) => 
                           PC2_out_22_port, A(21) => PC2_out_21_port, A(20) => 
                           PC2_out_20_port, A(19) => PC2_out_19_port, A(18) => 
                           PC2_out_18_port, A(17) => PC2_out_17_port, A(16) => 
                           PC2_out_16_port, A(15) => PC2_out_15_port, A(14) => 
                           PC2_out_14_port, A(13) => PC2_out_13_port, A(12) => 
                           PC2_out_12_port, A(11) => PC2_out_11_port, A(10) => 
                           PC2_out_10_port, A(9) => PC2_out_9_port, A(8) => 
                           PC2_out_8_port, A(7) => PC2_out_7_port, A(6) => 
                           PC2_out_6_port, A(5) => PC2_out_5_port, A(4) => 
                           PC2_out_4_port, A(3) => PC2_out_3_port, A(2) => 
                           PC2_out_2_port, A(1) => PC2_out_1_port, A(0) => 
                           PC2_out_0_port, B(31) => PC3_out_31_port, B(30) => 
                           PC3_out_30_port, B(29) => PC3_out_29_port, B(28) => 
                           PC3_out_28_port, B(27) => PC3_out_27_port, B(26) => 
                           PC3_out_26_port, B(25) => PC3_out_25_port, B(24) => 
                           PC3_out_24_port, B(23) => PC3_out_23_port, B(22) => 
                           PC3_out_22_port, B(21) => PC3_out_21_port, B(20) => 
                           PC3_out_20_port, B(19) => PC3_out_19_port, B(18) => 
                           PC3_out_18_port, B(17) => PC3_out_17_port, B(16) => 
                           PC3_out_16_port, B(15) => PC3_out_15_port, B(14) => 
                           PC3_out_14_port, B(13) => PC3_out_13_port, B(12) => 
                           PC3_out_12_port, B(11) => PC3_out_11_port, B(10) => 
                           PC3_out_10_port, B(9) => PC3_out_9_port, B(8) => 
                           PC3_out_8_port, B(7) => PC3_out_7_port, B(6) => 
                           PC3_out_6_port, B(5) => PC3_out_5_port, B(4) => 
                           PC3_out_4_port, B(3) => PC3_out_3_port, B(2) => 
                           PC3_out_2_port, B(1) => PC3_out_1_port, B(0) => 
                           PC3_out_0_port, SEL => n7, Y(31) => BHT_in_31_port, 
                           Y(30) => BHT_in_30_port, Y(29) => BHT_in_29_port, 
                           Y(28) => BHT_in_28_port, Y(27) => BHT_in_27_port, 
                           Y(26) => BHT_in_26_port, Y(25) => BHT_in_25_port, 
                           Y(24) => BHT_in_24_port, Y(23) => BHT_in_23_port, 
                           Y(22) => BHT_in_22_port, Y(21) => BHT_in_21_port, 
                           Y(20) => BHT_in_20_port, Y(19) => BHT_in_19_port, 
                           Y(18) => BHT_in_18_port, Y(17) => BHT_in_17_port, 
                           Y(16) => BHT_in_16_port, Y(15) => BHT_in_15_port, 
                           Y(14) => BHT_in_14_port, Y(13) => BHT_in_13_port, 
                           Y(12) => BHT_in_12_port, Y(11) => BHT_in_11_port, 
                           Y(10) => BHT_in_10_port, Y(9) => BHT_in_9_port, Y(8)
                           => BHT_in_8_port, Y(7) => BHT_in_7_port, Y(6) => 
                           BHT_in_6_port, Y(5) => BHT_in_5_port, Y(4) => 
                           BHT_in_4_port, Y(3) => BHT_in_3_port, Y(2) => 
                           BHT_in_2_port, Y(1) => BHT_in_1_port, Y(0) => 
                           BHT_in_0_port);
   RegAMUX : MUX2to1_NBIT32_6 port map( A(31) => FWDA_OUT_31_port, A(30) => 
                           FWDA_OUT_30_port, A(29) => FWDA_OUT_29_port, A(28) 
                           => FWDA_OUT_28_port, A(27) => FWDA_OUT_27_port, 
                           A(26) => FWDA_OUT_26_port, A(25) => FWDA_OUT_25_port
                           , A(24) => FWDA_OUT_24_port, A(23) => 
                           FWDA_OUT_23_port, A(22) => FWDA_OUT_22_port, A(21) 
                           => FWDA_OUT_21_port, A(20) => FWDA_OUT_20_port, 
                           A(19) => FWDA_OUT_19_port, A(18) => FWDA_OUT_18_port
                           , A(17) => FWDA_OUT_17_port, A(16) => 
                           FWDA_OUT_16_port, A(15) => FWDA_OUT_15_port, A(14) 
                           => FWDA_OUT_14_port, A(13) => FWDA_OUT_13_port, 
                           A(12) => FWDA_OUT_12_port, A(11) => FWDA_OUT_11_port
                           , A(10) => FWDA_OUT_10_port, A(9) => FWDA_OUT_9_port
                           , A(8) => FWDA_OUT_8_port, A(7) => FWDA_OUT_7_port, 
                           A(6) => FWDA_OUT_6_port, A(5) => FWDA_OUT_5_port, 
                           A(4) => FWDA_OUT_4_port, A(3) => FWDA_OUT_3_port, 
                           A(2) => FWDA_OUT_2_port, A(1) => FWDA_OUT_1_port, 
                           A(0) => FWDA_OUT_0_port, B(31) => X_Logic0_port, 
                           B(30) => X_Logic0_port, B(29) => X_Logic0_port, 
                           B(28) => X_Logic0_port, B(27) => X_Logic0_port, 
                           B(26) => X_Logic0_port, B(25) => X_Logic0_port, 
                           B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
                           B(22) => X_Logic0_port, B(21) => X_Logic0_port, 
                           B(20) => X_Logic0_port, B(19) => X_Logic0_port, 
                           B(18) => X_Logic0_port, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => X_Logic0_port, 
                           B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
                           B(12) => X_Logic0_port, B(11) => X_Logic0_port, 
                           B(10) => X_Logic0_port, B(9) => X_Logic0_port, B(8) 
                           => X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => ALUA_SEL, Y(31) => 
                           A_in_31_port, Y(30) => A_in_30_port, Y(29) => 
                           A_in_29_port, Y(28) => A_in_28_port, Y(27) => 
                           A_in_27_port, Y(26) => A_in_26_port, Y(25) => 
                           A_in_25_port, Y(24) => A_in_24_port, Y(23) => 
                           A_in_23_port, Y(22) => A_in_22_port, Y(21) => 
                           A_in_21_port, Y(20) => A_in_20_port, Y(19) => 
                           A_in_19_port, Y(18) => A_in_18_port, Y(17) => 
                           A_in_17_port, Y(16) => A_in_16_port, Y(15) => 
                           A_in_15_port, Y(14) => A_in_14_port, Y(13) => 
                           A_in_13_port, Y(12) => A_in_12_port, Y(11) => 
                           A_in_11_port, Y(10) => A_in_10_port, Y(9) => 
                           A_in_9_port, Y(8) => A_in_8_port, Y(7) => 
                           A_in_7_port, Y(6) => A_in_6_port, Y(5) => 
                           A_in_5_port, Y(4) => A_in_4_port, Y(3) => 
                           A_in_3_port, Y(2) => A_in_2_port, Y(1) => 
                           A_in_1_port, Y(0) => A_in_0_port);
   RegBMUX : MUX2to1_NBIT32_5 port map( A(31) => FWDB_OUT_31_port, A(30) => 
                           FWDB_OUT_30_port, A(29) => FWDB_OUT_29_port, A(28) 
                           => FWDB_OUT_28_port, A(27) => FWDB_OUT_27_port, 
                           A(26) => FWDB_OUT_26_port, A(25) => FWDB_OUT_25_port
                           , A(24) => FWDB_OUT_24_port, A(23) => 
                           FWDB_OUT_23_port, A(22) => FWDB_OUT_22_port, A(21) 
                           => FWDB_OUT_21_port, A(20) => FWDB_OUT_20_port, 
                           A(19) => FWDB_OUT_19_port, A(18) => FWDB_OUT_18_port
                           , A(17) => FWDB_OUT_17_port, A(16) => 
                           FWDB_OUT_16_port, A(15) => FWDB_OUT_15_port, A(14) 
                           => FWDB_OUT_14_port, A(13) => FWDB_OUT_13_port, 
                           A(12) => FWDB_OUT_12_port, A(11) => FWDB_OUT_11_port
                           , A(10) => FWDB_OUT_10_port, A(9) => FWDB_OUT_9_port
                           , A(8) => FWDB_OUT_8_port, A(7) => FWDB_OUT_7_port, 
                           A(6) => FWDB_OUT_6_port, A(5) => FWDB_OUT_5_port, 
                           A(4) => FWDB_OUT_4_port, A(3) => FWDB_OUT_3_port, 
                           A(2) => FWDB_OUT_2_port, A(1) => FWDB_OUT_1_port, 
                           A(0) => FWDB_OUT_0_port, B(31) => RIMM_out_31_port, 
                           B(30) => RIMM_out_30_port, B(29) => RIMM_out_29_port
                           , B(28) => RIMM_out_28_port, B(27) => 
                           RIMM_out_27_port, B(26) => RIMM_out_26_port, B(25) 
                           => RIMM_out_25_port, B(24) => RIMM_out_24_port, 
                           B(23) => RIMM_out_23_port, B(22) => RIMM_out_22_port
                           , B(21) => RIMM_out_21_port, B(20) => 
                           RIMM_out_20_port, B(19) => RIMM_out_19_port, B(18) 
                           => RIMM_out_18_port, B(17) => RIMM_out_17_port, 
                           B(16) => RIMM_out_16_port, B(15) => RIMM_out_15_port
                           , B(14) => RIMM_out_14_port, B(13) => 
                           RIMM_out_13_port, B(12) => RIMM_out_12_port, B(11) 
                           => RIMM_out_11_port, B(10) => RIMM_out_10_port, B(9)
                           => RIMM_out_9_port, B(8) => RIMM_out_8_port, B(7) =>
                           RIMM_out_7_port, B(6) => RIMM_out_6_port, B(5) => 
                           RIMM_out_5_port, B(4) => RIMM_out_4_port, B(3) => 
                           RIMM_out_3_port, B(2) => RIMM_out_2_port, B(1) => 
                           RIMM_out_1_port, B(0) => RIMM_out_0_port, SEL => 
                           ALUB_SEL, Y(31) => B_in_31_port, Y(30) => 
                           B_in_30_port, Y(29) => B_in_29_port, Y(28) => 
                           B_in_28_port, Y(27) => B_in_27_port, Y(26) => 
                           B_in_26_port, Y(25) => B_in_25_port, Y(24) => 
                           B_in_24_port, Y(23) => B_in_23_port, Y(22) => 
                           B_in_22_port, Y(21) => B_in_21_port, Y(20) => 
                           B_in_20_port, Y(19) => B_in_19_port, Y(18) => 
                           B_in_18_port, Y(17) => B_in_17_port, Y(16) => 
                           B_in_16_port, Y(15) => B_in_15_port, Y(14) => 
                           B_in_14_port, Y(13) => B_in_13_port, Y(12) => 
                           B_in_12_port, Y(11) => B_in_11_port, Y(10) => 
                           B_in_10_port, Y(9) => B_in_9_port, Y(8) => 
                           B_in_8_port, Y(7) => B_in_7_port, Y(6) => 
                           B_in_6_port, Y(5) => B_in_5_port, Y(4) => 
                           B_in_4_port, Y(3) => B_in_3_port, Y(2) => 
                           B_in_2_port, Y(1) => B_in_1_port, Y(0) => 
                           B_in_0_port);
   FWDA_MUX : MUX3to1_NBIT32_3 port map( A(31) => RA_out_31_port, A(30) => 
                           RA_out_30_port, A(29) => RA_out_29_port, A(28) => 
                           RA_out_28_port, A(27) => RA_out_27_port, A(26) => 
                           RA_out_26_port, A(25) => RA_out_25_port, A(24) => 
                           RA_out_24_port, A(23) => RA_out_23_port, A(22) => 
                           RA_out_22_port, A(21) => RA_out_21_port, A(20) => 
                           RA_out_20_port, A(19) => RA_out_19_port, A(18) => 
                           RA_out_18_port, A(17) => RA_out_17_port, A(16) => 
                           RA_out_16_port, A(15) => RA_out_15_port, A(14) => 
                           RA_out_14_port, A(13) => RA_out_13_port, A(12) => 
                           RA_out_12_port, A(11) => RA_out_11_port, A(10) => 
                           RA_out_10_port, A(9) => RA_out_9_port, A(8) => 
                           RA_out_8_port, A(7) => RA_out_7_port, A(6) => 
                           RA_out_6_port, A(5) => RA_out_5_port, A(4) => 
                           RA_out_4_port, A(3) => RA_out_3_port, A(2) => 
                           RA_out_2_port, A(1) => RA_out_1_port, A(0) => 
                           RA_out_0_port, B(31) => DATA_ADDR_31_port, B(30) => 
                           DATA_ADDR_30_port, B(29) => DATA_ADDR_29_port, B(28)
                           => DATA_ADDR_28_port, B(27) => DATA_ADDR_27_port, 
                           B(26) => DATA_ADDR_26_port, B(25) => 
                           DATA_ADDR_25_port, B(24) => DATA_ADDR_24_port, B(23)
                           => DATA_ADDR_23_port, B(22) => DATA_ADDR_22_port, 
                           B(21) => DATA_ADDR_21_port, B(20) => 
                           DATA_ADDR_20_port, B(19) => DATA_ADDR_19_port, B(18)
                           => DATA_ADDR_18_port, B(17) => DATA_ADDR_17_port, 
                           B(16) => DATA_ADDR_16_port, B(15) => 
                           DATA_ADDR_15_port, B(14) => DATA_ADDR_14_port, B(13)
                           => DATA_ADDR_13_port, B(12) => DATA_ADDR_12_port, 
                           B(11) => DATA_ADDR_11_port, B(10) => 
                           DATA_ADDR_10_port, B(9) => DATA_ADDR_9_port, B(8) =>
                           DATA_ADDR_8_port, B(7) => DATA_ADDR_7_port, B(6) => 
                           DATA_ADDR_6_port, B(5) => DATA_ADDR_5_port, B(4) => 
                           DATA_ADDR_4_port, B(3) => DATA_ADDR_3_port, B(2) => 
                           DATA_ADDR_2_port, B(1) => DATA_ADDR_1_port, B(0) => 
                           DATA_ADDR_0_port, C(31) => WB_in_31_port, C(30) => 
                           WB_in_30_port, C(29) => WB_in_29_port, C(28) => 
                           WB_in_28_port, C(27) => WB_in_27_port, C(26) => 
                           WB_in_26_port, C(25) => WB_in_25_port, C(24) => 
                           WB_in_24_port, C(23) => WB_in_23_port, C(22) => 
                           WB_in_22_port, C(21) => WB_in_21_port, C(20) => 
                           WB_in_20_port, C(19) => WB_in_19_port, C(18) => 
                           WB_in_18_port, C(17) => WB_in_17_port, C(16) => 
                           WB_in_16_port, C(15) => WB_in_15_port, C(14) => 
                           WB_in_14_port, C(13) => WB_in_13_port, C(12) => 
                           WB_in_12_port, C(11) => WB_in_11_port, C(10) => 
                           WB_in_10_port, C(9) => WB_in_9_port, C(8) => 
                           WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => FWDA_SEL_1_port, SEL(0) => 
                           FWDA_SEL_0_port, Y(31) => FWDA_OUT_31_port, Y(30) =>
                           FWDA_OUT_30_port, Y(29) => FWDA_OUT_29_port, Y(28) 
                           => FWDA_OUT_28_port, Y(27) => FWDA_OUT_27_port, 
                           Y(26) => FWDA_OUT_26_port, Y(25) => FWDA_OUT_25_port
                           , Y(24) => FWDA_OUT_24_port, Y(23) => 
                           FWDA_OUT_23_port, Y(22) => FWDA_OUT_22_port, Y(21) 
                           => FWDA_OUT_21_port, Y(20) => FWDA_OUT_20_port, 
                           Y(19) => FWDA_OUT_19_port, Y(18) => FWDA_OUT_18_port
                           , Y(17) => FWDA_OUT_17_port, Y(16) => 
                           FWDA_OUT_16_port, Y(15) => FWDA_OUT_15_port, Y(14) 
                           => FWDA_OUT_14_port, Y(13) => FWDA_OUT_13_port, 
                           Y(12) => FWDA_OUT_12_port, Y(11) => FWDA_OUT_11_port
                           , Y(10) => FWDA_OUT_10_port, Y(9) => FWDA_OUT_9_port
                           , Y(8) => FWDA_OUT_8_port, Y(7) => FWDA_OUT_7_port, 
                           Y(6) => FWDA_OUT_6_port, Y(5) => FWDA_OUT_5_port, 
                           Y(4) => FWDA_OUT_4_port, Y(3) => FWDA_OUT_3_port, 
                           Y(2) => FWDA_OUT_2_port, Y(1) => FWDA_OUT_1_port, 
                           Y(0) => FWDA_OUT_0_port);
   FWDB_MUX : MUX3to1_NBIT32_2 port map( A(31) => RB_out_31_port, A(30) => 
                           RB_out_30_port, A(29) => RB_out_29_port, A(28) => 
                           RB_out_28_port, A(27) => RB_out_27_port, A(26) => 
                           RB_out_26_port, A(25) => RB_out_25_port, A(24) => 
                           RB_out_24_port, A(23) => RB_out_23_port, A(22) => 
                           RB_out_22_port, A(21) => RB_out_21_port, A(20) => 
                           RB_out_20_port, A(19) => RB_out_19_port, A(18) => 
                           RB_out_18_port, A(17) => RB_out_17_port, A(16) => 
                           RB_out_16_port, A(15) => RB_out_15_port, A(14) => 
                           RB_out_14_port, A(13) => RB_out_13_port, A(12) => 
                           RB_out_12_port, A(11) => RB_out_11_port, A(10) => 
                           RB_out_10_port, A(9) => RB_out_9_port, A(8) => 
                           RB_out_8_port, A(7) => RB_out_7_port, A(6) => 
                           RB_out_6_port, A(5) => RB_out_5_port, A(4) => 
                           RB_out_4_port, A(3) => RB_out_3_port, A(2) => 
                           RB_out_2_port, A(1) => RB_out_1_port, A(0) => 
                           RB_out_0_port, B(31) => DATA_ADDR_31_port, B(30) => 
                           DATA_ADDR_30_port, B(29) => DATA_ADDR_29_port, B(28)
                           => DATA_ADDR_28_port, B(27) => DATA_ADDR_27_port, 
                           B(26) => DATA_ADDR_26_port, B(25) => 
                           DATA_ADDR_25_port, B(24) => DATA_ADDR_24_port, B(23)
                           => DATA_ADDR_23_port, B(22) => DATA_ADDR_22_port, 
                           B(21) => DATA_ADDR_21_port, B(20) => 
                           DATA_ADDR_20_port, B(19) => DATA_ADDR_19_port, B(18)
                           => DATA_ADDR_18_port, B(17) => DATA_ADDR_17_port, 
                           B(16) => DATA_ADDR_16_port, B(15) => 
                           DATA_ADDR_15_port, B(14) => DATA_ADDR_14_port, B(13)
                           => DATA_ADDR_13_port, B(12) => DATA_ADDR_12_port, 
                           B(11) => DATA_ADDR_11_port, B(10) => 
                           DATA_ADDR_10_port, B(9) => DATA_ADDR_9_port, B(8) =>
                           DATA_ADDR_8_port, B(7) => DATA_ADDR_7_port, B(6) => 
                           DATA_ADDR_6_port, B(5) => DATA_ADDR_5_port, B(4) => 
                           DATA_ADDR_4_port, B(3) => DATA_ADDR_3_port, B(2) => 
                           DATA_ADDR_2_port, B(1) => DATA_ADDR_1_port, B(0) => 
                           DATA_ADDR_0_port, C(31) => WB_in_31_port, C(30) => 
                           WB_in_30_port, C(29) => WB_in_29_port, C(28) => 
                           WB_in_28_port, C(27) => WB_in_27_port, C(26) => 
                           WB_in_26_port, C(25) => WB_in_25_port, C(24) => 
                           WB_in_24_port, C(23) => WB_in_23_port, C(22) => 
                           WB_in_22_port, C(21) => WB_in_21_port, C(20) => 
                           WB_in_20_port, C(19) => WB_in_19_port, C(18) => 
                           WB_in_18_port, C(17) => WB_in_17_port, C(16) => 
                           WB_in_16_port, C(15) => WB_in_15_port, C(14) => 
                           WB_in_14_port, C(13) => WB_in_13_port, C(12) => 
                           WB_in_12_port, C(11) => WB_in_11_port, C(10) => 
                           WB_in_10_port, C(9) => WB_in_9_port, C(8) => 
                           WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => FWDB_SEL_1_port, SEL(0) => 
                           FWDB_SEL_0_port, Y(31) => FWDB_OUT_31_port, Y(30) =>
                           FWDB_OUT_30_port, Y(29) => FWDB_OUT_29_port, Y(28) 
                           => FWDB_OUT_28_port, Y(27) => FWDB_OUT_27_port, 
                           Y(26) => FWDB_OUT_26_port, Y(25) => FWDB_OUT_25_port
                           , Y(24) => FWDB_OUT_24_port, Y(23) => 
                           FWDB_OUT_23_port, Y(22) => FWDB_OUT_22_port, Y(21) 
                           => FWDB_OUT_21_port, Y(20) => FWDB_OUT_20_port, 
                           Y(19) => FWDB_OUT_19_port, Y(18) => FWDB_OUT_18_port
                           , Y(17) => FWDB_OUT_17_port, Y(16) => 
                           FWDB_OUT_16_port, Y(15) => FWDB_OUT_15_port, Y(14) 
                           => FWDB_OUT_14_port, Y(13) => FWDB_OUT_13_port, 
                           Y(12) => FWDB_OUT_12_port, Y(11) => FWDB_OUT_11_port
                           , Y(10) => FWDB_OUT_10_port, Y(9) => FWDB_OUT_9_port
                           , Y(8) => FWDB_OUT_8_port, Y(7) => FWDB_OUT_7_port, 
                           Y(6) => FWDB_OUT_6_port, Y(5) => FWDB_OUT_5_port, 
                           Y(4) => FWDB_OUT_4_port, Y(3) => FWDB_OUT_3_port, 
                           Y(2) => FWDB_OUT_2_port, Y(1) => FWDB_OUT_1_port, 
                           Y(0) => FWDB_OUT_0_port);
   ZDU_MUX : MUX3to1_NBIT32_1 port map( A(31) => RA_out_31_port, A(30) => 
                           RA_out_30_port, A(29) => RA_out_29_port, A(28) => 
                           RA_out_28_port, A(27) => RA_out_27_port, A(26) => 
                           RA_out_26_port, A(25) => RA_out_25_port, A(24) => 
                           RA_out_24_port, A(23) => RA_out_23_port, A(22) => 
                           RA_out_22_port, A(21) => RA_out_21_port, A(20) => 
                           RA_out_20_port, A(19) => RA_out_19_port, A(18) => 
                           RA_out_18_port, A(17) => RA_out_17_port, A(16) => 
                           RA_out_16_port, A(15) => RA_out_15_port, A(14) => 
                           RA_out_14_port, A(13) => RA_out_13_port, A(12) => 
                           RA_out_12_port, A(11) => RA_out_11_port, A(10) => 
                           RA_out_10_port, A(9) => RA_out_9_port, A(8) => 
                           RA_out_8_port, A(7) => RA_out_7_port, A(6) => 
                           RA_out_6_port, A(5) => RA_out_5_port, A(4) => 
                           RA_out_4_port, A(3) => RA_out_3_port, A(2) => 
                           RA_out_2_port, A(1) => RA_out_1_port, A(0) => 
                           RA_out_0_port, B(31) => CWB_MUX2_out_31_port, B(30) 
                           => CWB_MUX2_out_30_port, B(29) => 
                           CWB_MUX2_out_29_port, B(28) => CWB_MUX2_out_28_port,
                           B(27) => CWB_MUX2_out_27_port, B(26) => 
                           CWB_MUX2_out_26_port, B(25) => CWB_MUX2_out_25_port,
                           B(24) => CWB_MUX2_out_24_port, B(23) => 
                           CWB_MUX2_out_23_port, B(22) => CWB_MUX2_out_22_port,
                           B(21) => CWB_MUX2_out_21_port, B(20) => 
                           CWB_MUX2_out_20_port, B(19) => CWB_MUX2_out_19_port,
                           B(18) => CWB_MUX2_out_18_port, B(17) => 
                           CWB_MUX2_out_17_port, B(16) => CWB_MUX2_out_16_port,
                           B(15) => CWB_MUX2_out_15_port, B(14) => 
                           CWB_MUX2_out_14_port, B(13) => CWB_MUX2_out_13_port,
                           B(12) => CWB_MUX2_out_12_port, B(11) => 
                           CWB_MUX2_out_11_port, B(10) => CWB_MUX2_out_10_port,
                           B(9) => CWB_MUX2_out_9_port, B(8) => 
                           CWB_MUX2_out_8_port, B(7) => CWB_MUX2_out_7_port, 
                           B(6) => CWB_MUX2_out_6_port, B(5) => 
                           CWB_MUX2_out_5_port, B(4) => CWB_MUX2_out_4_port, 
                           B(3) => CWB_MUX2_out_3_port, B(2) => 
                           CWB_MUX2_out_2_port, B(1) => CWB_MUX2_out_1_port, 
                           B(0) => CWB_MUX2_out_0_port, C(31) => WB_in_31_port,
                           C(30) => WB_in_30_port, C(29) => WB_in_29_port, 
                           C(28) => WB_in_28_port, C(27) => WB_in_27_port, 
                           C(26) => WB_in_26_port, C(25) => WB_in_25_port, 
                           C(24) => WB_in_24_port, C(23) => WB_in_23_port, 
                           C(22) => WB_in_22_port, C(21) => WB_in_21_port, 
                           C(20) => WB_in_20_port, C(19) => WB_in_19_port, 
                           C(18) => WB_in_18_port, C(17) => WB_in_17_port, 
                           C(16) => WB_in_16_port, C(15) => WB_in_15_port, 
                           C(14) => WB_in_14_port, C(13) => WB_in_13_port, 
                           C(12) => WB_in_12_port, C(11) => WB_in_11_port, 
                           C(10) => WB_in_10_port, C(9) => WB_in_9_port, C(8) 
                           => WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => ZDU_SEL_1_port, SEL(0) => 
                           ZDU_SEL_0_port, Y(31) => n_1791, Y(30) => 
                           ZDU_MUX_out_30_port, Y(29) => ZDU_MUX_out_29_port, 
                           Y(28) => ZDU_MUX_out_28_port, Y(27) => 
                           ZDU_MUX_out_27_port, Y(26) => ZDU_MUX_out_26_port, 
                           Y(25) => ZDU_MUX_out_25_port, Y(24) => 
                           ZDU_MUX_out_24_port, Y(23) => ZDU_MUX_out_23_port, 
                           Y(22) => ZDU_MUX_out_22_port, Y(21) => 
                           ZDU_MUX_out_21_port, Y(20) => ZDU_MUX_out_20_port, 
                           Y(19) => ZDU_MUX_out_19_port, Y(18) => 
                           ZDU_MUX_out_18_port, Y(17) => ZDU_MUX_out_17_port, 
                           Y(16) => ZDU_MUX_out_16_port, Y(15) => 
                           ZDU_MUX_out_15_port, Y(14) => ZDU_MUX_out_14_port, 
                           Y(13) => ZDU_MUX_out_13_port, Y(12) => 
                           ZDU_MUX_out_12_port, Y(11) => ZDU_MUX_out_11_port, 
                           Y(10) => ZDU_MUX_out_10_port, Y(9) => 
                           ZDU_MUX_out_9_port, Y(8) => ZDU_MUX_out_8_port, Y(7)
                           => ZDU_MUX_out_7_port, Y(6) => ZDU_MUX_out_6_port, 
                           Y(5) => ZDU_MUX_out_5_port, Y(4) => 
                           ZDU_MUX_out_4_port, Y(3) => ZDU_MUX_out_3_port, Y(2)
                           => ZDU_MUX_out_2_port, Y(1) => ZDU_MUX_out_1_port, 
                           Y(0) => ZDU_MUX_out_0_port);
   MEMDATAMUX : MUX2to1_NBIT32_4 port map( A(31) => ALR2_out_31_port, A(30) => 
                           ALR2_out_30_port, A(29) => ALR2_out_29_port, A(28) 
                           => ALR2_out_28_port, A(27) => ALR2_out_27_port, 
                           A(26) => ALR2_out_26_port, A(25) => ALR2_out_25_port
                           , A(24) => ALR2_out_24_port, A(23) => 
                           ALR2_out_23_port, A(22) => ALR2_out_22_port, A(21) 
                           => ALR2_out_21_port, A(20) => ALR2_out_20_port, 
                           A(19) => ALR2_out_19_port, A(18) => ALR2_out_18_port
                           , A(17) => ALR2_out_17_port, A(16) => 
                           ALR2_out_16_port, A(15) => ALR2_out_15_port, A(14) 
                           => ALR2_out_14_port, A(13) => ALR2_out_13_port, 
                           A(12) => ALR2_out_12_port, A(11) => ALR2_out_11_port
                           , A(10) => ALR2_out_10_port, A(9) => ALR2_out_9_port
                           , A(8) => ALR2_out_8_port, A(7) => ALR2_out_7_port, 
                           A(6) => ALR2_out_6_port, A(5) => ALR2_out_5_port, 
                           A(4) => ALR2_out_4_port, A(3) => ALR2_out_3_port, 
                           A(2) => ALR2_out_2_port, A(1) => ALR2_out_1_port, 
                           A(0) => ALR2_out_0_port, B(31) => B2_MUX_out_31_port
                           , B(30) => B2_MUX_out_30_port, B(29) => 
                           B2_MUX_out_29_port, B(28) => B2_MUX_out_28_port, 
                           B(27) => B2_MUX_out_27_port, B(26) => 
                           B2_MUX_out_26_port, B(25) => B2_MUX_out_25_port, 
                           B(24) => B2_MUX_out_24_port, B(23) => 
                           B2_MUX_out_23_port, B(22) => B2_MUX_out_22_port, 
                           B(21) => B2_MUX_out_21_port, B(20) => 
                           B2_MUX_out_20_port, B(19) => B2_MUX_out_19_port, 
                           B(18) => B2_MUX_out_18_port, B(17) => 
                           B2_MUX_out_17_port, B(16) => B2_MUX_out_16_port, 
                           B(15) => B2_MUX_out_15_port, B(14) => 
                           B2_MUX_out_14_port, B(13) => B2_MUX_out_13_port, 
                           B(12) => B2_MUX_out_12_port, B(11) => 
                           B2_MUX_out_11_port, B(10) => B2_MUX_out_10_port, 
                           B(9) => B2_MUX_out_9_port, B(8) => B2_MUX_out_8_port
                           , B(7) => B2_MUX_out_7_port, B(6) => 
                           B2_MUX_out_6_port, B(5) => B2_MUX_out_5_port, B(4) 
                           => B2_MUX_out_4_port, B(3) => B2_MUX_out_3_port, 
                           B(2) => B2_MUX_out_2_port, B(1) => B2_MUX_out_1_port
                           , B(0) => B2_MUX_out_0_port, SEL => MEM_DATA_SEL, 
                           Y(31) => DATA_OUT(31), Y(30) => DATA_OUT(30), Y(29) 
                           => DATA_OUT(29), Y(28) => DATA_OUT(28), Y(27) => 
                           DATA_OUT(27), Y(26) => DATA_OUT(26), Y(25) => 
                           DATA_OUT(25), Y(24) => DATA_OUT(24), Y(23) => 
                           DATA_OUT(23), Y(22) => DATA_OUT(22), Y(21) => 
                           DATA_OUT(21), Y(20) => DATA_OUT(20), Y(19) => 
                           DATA_OUT(19), Y(18) => DATA_OUT(18), Y(17) => 
                           DATA_OUT(17), Y(16) => DATA_OUT(16), Y(15) => 
                           DATA_OUT(15), Y(14) => DATA_OUT(14), Y(13) => 
                           DATA_OUT(13), Y(12) => DATA_OUT(12), Y(11) => 
                           DATA_OUT(11), Y(10) => DATA_OUT(10), Y(9) => 
                           DATA_OUT(9), Y(8) => DATA_OUT(8), Y(7) => 
                           DATA_OUT(7), Y(6) => DATA_OUT(6), Y(5) => 
                           DATA_OUT(5), Y(4) => DATA_OUT(4), Y(3) => 
                           DATA_OUT(3), Y(2) => DATA_OUT(2), Y(1) => 
                           DATA_OUT(1), Y(0) => DATA_OUT(0));
   LMDMUX : MUX5to1_NBIT32_0 port map( A(31) => n12, A(30) => DATA_IN(6), A(29)
                           => DATA_IN(5), A(28) => DATA_IN(4), A(27) => 
                           DATA_IN(3), A(26) => DATA_IN(2), A(25) => DATA_IN(1)
                           , A(24) => DATA_IN(0), A(23) => DATA_IN(15), A(22) 
                           => DATA_IN(14), A(21) => DATA_IN(13), A(20) => 
                           DATA_IN(12), A(19) => DATA_IN(11), A(18) => 
                           DATA_IN(10), A(17) => DATA_IN(9), A(16) => 
                           DATA_IN(8), A(15) => DATA_IN(23), A(14) => 
                           DATA_IN(22), A(13) => DATA_IN(21), A(12) => 
                           DATA_IN(20), A(11) => DATA_IN(19), A(10) => 
                           DATA_IN(18), A(9) => DATA_IN(17), A(8) => 
                           DATA_IN(16), A(7) => DATA_IN(31), A(6) => 
                           DATA_IN(30), A(5) => DATA_IN(29), A(4) => 
                           DATA_IN(28), A(3) => DATA_IN(27), A(2) => 
                           DATA_IN(26), A(1) => DATA_IN(25), A(0) => 
                           DATA_IN(24), B(31) => n10, B(30) => n10, B(29) => 
                           n10, B(28) => n10, B(27) => n10, B(26) => n10, B(25)
                           => n10, B(24) => n10, B(23) => n10, B(22) => n10, 
                           B(21) => n10, B(20) => n11, B(19) => n11, B(18) => 
                           n11, B(17) => n11, B(16) => n11, B(15) => n11, B(14)
                           => n11, B(13) => n11, B(12) => n11, B(11) => n11, 
                           B(10) => n11, B(9) => n11, B(8) => n12, B(7) => n12,
                           B(6) => DATA_IN(6), B(5) => DATA_IN(5), B(4) => 
                           DATA_IN(4), B(3) => DATA_IN(3), B(2) => DATA_IN(2), 
                           B(1) => DATA_IN(1), B(0) => DATA_IN(0), C(31) => 
                           X_Logic0_port, C(30) => X_Logic0_port, C(29) => 
                           X_Logic0_port, C(28) => X_Logic0_port, C(27) => 
                           X_Logic0_port, C(26) => X_Logic0_port, C(25) => 
                           X_Logic0_port, C(24) => X_Logic0_port, C(23) => 
                           X_Logic0_port, C(22) => X_Logic0_port, C(21) => 
                           X_Logic0_port, C(20) => X_Logic0_port, C(19) => 
                           X_Logic0_port, C(18) => X_Logic0_port, C(17) => 
                           X_Logic0_port, C(16) => X_Logic0_port, C(15) => 
                           X_Logic0_port, C(14) => X_Logic0_port, C(13) => 
                           X_Logic0_port, C(12) => X_Logic0_port, C(11) => 
                           X_Logic0_port, C(10) => X_Logic0_port, C(9) => 
                           X_Logic0_port, C(8) => X_Logic0_port, C(7) => n10, 
                           C(6) => DATA_IN(6), C(5) => DATA_IN(5), C(4) => 
                           DATA_IN(4), C(3) => DATA_IN(3), C(2) => DATA_IN(2), 
                           C(1) => DATA_IN(1), C(0) => DATA_IN(0), D(31) => n12
                           , D(30) => n12, D(29) => n12, D(28) => n12, D(27) =>
                           n12, D(26) => n12, D(25) => n12, D(24) => n19, D(23)
                           => n12, D(22) => n19, D(21) => n19, D(20) => n19, 
                           D(19) => n19, D(18) => n19, D(17) => n19, D(16) => 
                           n19, D(15) => n19, D(14) => DATA_IN(6), D(13) => 
                           DATA_IN(5), D(12) => DATA_IN(4), D(11) => DATA_IN(3)
                           , D(10) => DATA_IN(2), D(9) => DATA_IN(1), D(8) => 
                           DATA_IN(0), D(7) => DATA_IN(15), D(6) => DATA_IN(14)
                           , D(5) => DATA_IN(13), D(4) => DATA_IN(12), D(3) => 
                           DATA_IN(11), D(2) => DATA_IN(10), D(1) => DATA_IN(9)
                           , D(0) => DATA_IN(8), E(31) => X_Logic0_port, E(30) 
                           => X_Logic0_port, E(29) => X_Logic0_port, E(28) => 
                           X_Logic0_port, E(27) => X_Logic0_port, E(26) => 
                           X_Logic0_port, E(25) => X_Logic0_port, E(24) => 
                           X_Logic0_port, E(23) => X_Logic0_port, E(22) => 
                           X_Logic0_port, E(21) => X_Logic0_port, E(20) => 
                           X_Logic0_port, E(19) => X_Logic0_port, E(18) => 
                           X_Logic0_port, E(17) => X_Logic0_port, E(16) => 
                           X_Logic0_port, E(15) => n12, E(14) => DATA_IN(6), 
                           E(13) => DATA_IN(5), E(12) => DATA_IN(4), E(11) => 
                           DATA_IN(3), E(10) => DATA_IN(2), E(9) => DATA_IN(1),
                           E(8) => DATA_IN(0), E(7) => DATA_IN(15), E(6) => 
                           DATA_IN(14), E(5) => DATA_IN(13), E(4) => 
                           DATA_IN(12), E(3) => DATA_IN(11), E(2) => 
                           DATA_IN(10), E(1) => DATA_IN(9), E(0) => DATA_IN(8),
                           SEL(2) => LD_SEL(2), SEL(1) => LD_SEL(1), SEL(0) => 
                           LD_SEL(0), Y(31) => LMD_out_31_port, Y(30) => 
                           LMD_out_30_port, Y(29) => LMD_out_29_port, Y(28) => 
                           LMD_out_28_port, Y(27) => LMD_out_27_port, Y(26) => 
                           LMD_out_26_port, Y(25) => LMD_out_25_port, Y(24) => 
                           LMD_out_24_port, Y(23) => LMD_out_23_port, Y(22) => 
                           LMD_out_22_port, Y(21) => LMD_out_21_port, Y(20) => 
                           LMD_out_20_port, Y(19) => LMD_out_19_port, Y(18) => 
                           LMD_out_18_port, Y(17) => LMD_out_17_port, Y(16) => 
                           LMD_out_16_port, Y(15) => LMD_out_15_port, Y(14) => 
                           LMD_out_14_port, Y(13) => LMD_out_13_port, Y(12) => 
                           LMD_out_12_port, Y(11) => LMD_out_11_port, Y(10) => 
                           LMD_out_10_port, Y(9) => LMD_out_9_port, Y(8) => 
                           LMD_out_8_port, Y(7) => LMD_out_7_port, Y(6) => 
                           LMD_out_6_port, Y(5) => LMD_out_5_port, Y(4) => 
                           LMD_out_4_port, Y(3) => LMD_out_3_port, Y(2) => 
                           LMD_out_2_port, Y(1) => LMD_out_1_port, Y(0) => 
                           LMD_out_0_port);
   ALR2_MUX : MUX2to1_NBIT32_3 port map( A(31) => CWB_MUX2_out_31_port, A(30) 
                           => CWB_MUX2_out_30_port, A(29) => 
                           CWB_MUX2_out_29_port, A(28) => CWB_MUX2_out_28_port,
                           A(27) => CWB_MUX2_out_27_port, A(26) => 
                           CWB_MUX2_out_26_port, A(25) => CWB_MUX2_out_25_port,
                           A(24) => CWB_MUX2_out_24_port, A(23) => 
                           CWB_MUX2_out_23_port, A(22) => CWB_MUX2_out_22_port,
                           A(21) => CWB_MUX2_out_21_port, A(20) => 
                           CWB_MUX2_out_20_port, A(19) => CWB_MUX2_out_19_port,
                           A(18) => CWB_MUX2_out_18_port, A(17) => 
                           CWB_MUX2_out_17_port, A(16) => CWB_MUX2_out_16_port,
                           A(15) => CWB_MUX2_out_15_port, A(14) => 
                           CWB_MUX2_out_14_port, A(13) => CWB_MUX2_out_13_port,
                           A(12) => CWB_MUX2_out_12_port, A(11) => 
                           CWB_MUX2_out_11_port, A(10) => CWB_MUX2_out_10_port,
                           A(9) => CWB_MUX2_out_9_port, A(8) => 
                           CWB_MUX2_out_8_port, A(7) => CWB_MUX2_out_7_port, 
                           A(6) => CWB_MUX2_out_6_port, A(5) => 
                           CWB_MUX2_out_5_port, A(4) => CWB_MUX2_out_4_port, 
                           A(3) => CWB_MUX2_out_3_port, A(2) => 
                           CWB_MUX2_out_2_port, A(1) => CWB_MUX2_out_1_port, 
                           A(0) => CWB_MUX2_out_0_port, B(31) => 
                           NPC3_out_31_port, B(30) => NPC3_out_30_port, B(29) 
                           => NPC3_out_29_port, B(28) => NPC3_out_28_port, 
                           B(27) => NPC3_out_27_port, B(26) => NPC3_out_26_port
                           , B(25) => NPC3_out_25_port, B(24) => 
                           NPC3_out_24_port, B(23) => NPC3_out_23_port, B(22) 
                           => NPC3_out_22_port, B(21) => NPC3_out_21_port, 
                           B(20) => NPC3_out_20_port, B(19) => NPC3_out_19_port
                           , B(18) => NPC3_out_18_port, B(17) => 
                           NPC3_out_17_port, B(16) => NPC3_out_16_port, B(15) 
                           => NPC3_out_15_port, B(14) => NPC3_out_14_port, 
                           B(13) => NPC3_out_13_port, B(12) => NPC3_out_12_port
                           , B(11) => NPC3_out_11_port, B(10) => 
                           NPC3_out_10_port, B(9) => NPC3_out_9_port, B(8) => 
                           NPC3_out_8_port, B(7) => NPC3_out_7_port, B(6) => 
                           NPC3_out_6_port, B(5) => NPC3_out_5_port, B(4) => 
                           NPC3_out_4_port, B(3) => NPC3_out_3_port, B(2) => 
                           NPC3_out_2_port, B(1) => NPC3_out_1_port, B(0) => 
                           NPC3_out_0_port, SEL => ALR2_SEL, Y(31) => 
                           ALR2_in_31_port, Y(30) => ALR2_in_30_port, Y(29) => 
                           ALR2_in_29_port, Y(28) => ALR2_in_28_port, Y(27) => 
                           ALR2_in_27_port, Y(26) => ALR2_in_26_port, Y(25) => 
                           ALR2_in_25_port, Y(24) => ALR2_in_24_port, Y(23) => 
                           ALR2_in_23_port, Y(22) => ALR2_in_22_port, Y(21) => 
                           ALR2_in_21_port, Y(20) => ALR2_in_20_port, Y(19) => 
                           ALR2_in_19_port, Y(18) => ALR2_in_18_port, Y(17) => 
                           ALR2_in_17_port, Y(16) => ALR2_in_16_port, Y(15) => 
                           ALR2_in_15_port, Y(14) => ALR2_in_14_port, Y(13) => 
                           ALR2_in_13_port, Y(12) => ALR2_in_12_port, Y(11) => 
                           ALR2_in_11_port, Y(10) => ALR2_in_10_port, Y(9) => 
                           ALR2_in_9_port, Y(8) => ALR2_in_8_port, Y(7) => 
                           ALR2_in_7_port, Y(6) => ALR2_in_6_port, Y(5) => 
                           ALR2_in_5_port, Y(4) => ALR2_in_4_port, Y(3) => 
                           ALR2_in_3_port, Y(2) => ALR2_in_2_port, Y(1) => 
                           ALR2_in_1_port, Y(0) => ALR2_in_0_port);
   CWB_MUX1 : MUX3to1_NBIT2 port map( A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, C(1) => CWB_out_1_port, C(0) => 
                           CWB_out_0_port, SEL(1) => CWB_MUX_SEL_1_port, SEL(0)
                           => CWB_MUX_SEL_0_port, Y(1) => CWB2_SEL_1_port, Y(0)
                           => CWB2_SEL_0_port);
   CWB_MUX2 : MUX4to1_NBIT32_0 port map( A(31) => DATA_ADDR_31_port, A(30) => 
                           DATA_ADDR_30_port, A(29) => DATA_ADDR_29_port, A(28)
                           => DATA_ADDR_28_port, A(27) => DATA_ADDR_27_port, 
                           A(26) => DATA_ADDR_26_port, A(25) => 
                           DATA_ADDR_25_port, A(24) => DATA_ADDR_24_port, A(23)
                           => DATA_ADDR_23_port, A(22) => DATA_ADDR_22_port, 
                           A(21) => DATA_ADDR_21_port, A(20) => 
                           DATA_ADDR_20_port, A(19) => DATA_ADDR_19_port, A(18)
                           => DATA_ADDR_18_port, A(17) => DATA_ADDR_17_port, 
                           A(16) => DATA_ADDR_16_port, A(15) => 
                           DATA_ADDR_15_port, A(14) => DATA_ADDR_14_port, A(13)
                           => DATA_ADDR_13_port, A(12) => DATA_ADDR_12_port, 
                           A(11) => DATA_ADDR_11_port, A(10) => 
                           DATA_ADDR_10_port, A(9) => DATA_ADDR_9_port, A(8) =>
                           DATA_ADDR_8_port, A(7) => DATA_ADDR_7_port, A(6) => 
                           DATA_ADDR_6_port, A(5) => DATA_ADDR_5_port, A(4) => 
                           DATA_ADDR_4_port, A(3) => DATA_ADDR_3_port, A(2) => 
                           DATA_ADDR_2_port, A(1) => DATA_ADDR_1_port, A(0) => 
                           DATA_ADDR_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, C(31) => X_Logic0_port, C(30) => 
                           X_Logic0_port, C(29) => X_Logic0_port, C(28) => 
                           X_Logic0_port, C(27) => X_Logic0_port, C(26) => 
                           X_Logic0_port, C(25) => X_Logic0_port, C(24) => 
                           X_Logic0_port, C(23) => X_Logic0_port, C(22) => 
                           X_Logic0_port, C(21) => X_Logic0_port, C(20) => 
                           X_Logic0_port, C(19) => X_Logic0_port, C(18) => 
                           X_Logic0_port, C(17) => X_Logic0_port, C(16) => 
                           X_Logic0_port, C(15) => X_Logic0_port, C(14) => 
                           X_Logic0_port, C(13) => X_Logic0_port, C(12) => 
                           X_Logic0_port, C(11) => X_Logic0_port, C(10) => 
                           X_Logic0_port, C(9) => X_Logic0_port, C(8) => 
                           X_Logic0_port, C(7) => X_Logic0_port, C(6) => 
                           X_Logic0_port, C(5) => X_Logic0_port, C(4) => 
                           X_Logic0_port, C(3) => X_Logic0_port, C(2) => 
                           X_Logic0_port, C(1) => X_Logic0_port, C(0) => 
                           X_Logic0_port, D(31) => DATA_ADDR_15_port, D(30) => 
                           DATA_ADDR_14_port, D(29) => DATA_ADDR_13_port, D(28)
                           => DATA_ADDR_12_port, D(27) => DATA_ADDR_11_port, 
                           D(26) => DATA_ADDR_10_port, D(25) => 
                           DATA_ADDR_9_port, D(24) => DATA_ADDR_8_port, D(23) 
                           => DATA_ADDR_7_port, D(22) => DATA_ADDR_6_port, 
                           D(21) => DATA_ADDR_5_port, D(20) => DATA_ADDR_4_port
                           , D(19) => DATA_ADDR_3_port, D(18) => 
                           DATA_ADDR_2_port, D(17) => DATA_ADDR_1_port, D(16) 
                           => DATA_ADDR_0_port, D(15) => X_Logic0_port, D(14) 
                           => X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, SEL(1) => CWB2_SEL_1_port, SEL(0) => 
                           CWB2_SEL_0_port, Y(31) => CWB_MUX2_out_31_port, 
                           Y(30) => CWB_MUX2_out_30_port, Y(29) => 
                           CWB_MUX2_out_29_port, Y(28) => CWB_MUX2_out_28_port,
                           Y(27) => CWB_MUX2_out_27_port, Y(26) => 
                           CWB_MUX2_out_26_port, Y(25) => CWB_MUX2_out_25_port,
                           Y(24) => CWB_MUX2_out_24_port, Y(23) => 
                           CWB_MUX2_out_23_port, Y(22) => CWB_MUX2_out_22_port,
                           Y(21) => CWB_MUX2_out_21_port, Y(20) => 
                           CWB_MUX2_out_20_port, Y(19) => CWB_MUX2_out_19_port,
                           Y(18) => CWB_MUX2_out_18_port, Y(17) => 
                           CWB_MUX2_out_17_port, Y(16) => CWB_MUX2_out_16_port,
                           Y(15) => CWB_MUX2_out_15_port, Y(14) => 
                           CWB_MUX2_out_14_port, Y(13) => CWB_MUX2_out_13_port,
                           Y(12) => CWB_MUX2_out_12_port, Y(11) => 
                           CWB_MUX2_out_11_port, Y(10) => CWB_MUX2_out_10_port,
                           Y(9) => CWB_MUX2_out_9_port, Y(8) => 
                           CWB_MUX2_out_8_port, Y(7) => CWB_MUX2_out_7_port, 
                           Y(6) => CWB_MUX2_out_6_port, Y(5) => 
                           CWB_MUX2_out_5_port, Y(4) => CWB_MUX2_out_4_port, 
                           Y(3) => CWB_MUX2_out_3_port, Y(2) => 
                           CWB_MUX2_out_2_port, Y(1) => CWB_MUX2_out_1_port, 
                           Y(0) => CWB_MUX2_out_0_port);
   B2_MUX : MUX2to1_NBIT32_2 port map( A(31) => B2_out_31_port, A(30) => 
                           B2_out_30_port, A(29) => B2_out_29_port, A(28) => 
                           B2_out_28_port, A(27) => B2_out_27_port, A(26) => 
                           B2_out_26_port, A(25) => B2_out_25_port, A(24) => 
                           B2_out_24_port, A(23) => B2_out_23_port, A(22) => 
                           B2_out_22_port, A(21) => B2_out_21_port, A(20) => 
                           B2_out_20_port, A(19) => B2_out_19_port, A(18) => 
                           B2_out_18_port, A(17) => B2_out_17_port, A(16) => 
                           B2_out_16_port, A(15) => B2_out_15_port, A(14) => 
                           B2_out_14_port, A(13) => B2_out_13_port, A(12) => 
                           B2_out_12_port, A(11) => B2_out_11_port, A(10) => 
                           B2_out_10_port, A(9) => B2_out_9_port, A(8) => 
                           B2_out_8_port, A(7) => B2_out_7_port, A(6) => 
                           B2_out_6_port, A(5) => B2_out_5_port, A(4) => 
                           B2_out_4_port, A(3) => B2_out_3_port, A(2) => 
                           B2_out_2_port, A(1) => B2_out_1_port, A(0) => 
                           B2_out_0_port, B(31) => WB_in_31_port, B(30) => 
                           WB_in_30_port, B(29) => WB_in_29_port, B(28) => 
                           WB_in_28_port, B(27) => WB_in_27_port, B(26) => 
                           WB_in_26_port, B(25) => WB_in_25_port, B(24) => 
                           WB_in_24_port, B(23) => WB_in_23_port, B(22) => 
                           WB_in_22_port, B(21) => WB_in_21_port, B(20) => 
                           WB_in_20_port, B(19) => WB_in_19_port, B(18) => 
                           WB_in_18_port, B(17) => WB_in_17_port, B(16) => 
                           WB_in_16_port, B(15) => WB_in_15_port, B(14) => 
                           WB_in_14_port, B(13) => WB_in_13_port, B(12) => 
                           WB_in_12_port, B(11) => WB_in_11_port, B(10) => 
                           WB_in_10_port, B(9) => WB_in_9_port, B(8) => 
                           WB_in_8_port, B(7) => WB_in_7_port, B(6) => 
                           WB_in_6_port, B(5) => WB_in_5_port, B(4) => 
                           WB_in_4_port, B(3) => WB_in_3_port, B(2) => 
                           WB_in_2_port, B(1) => WB_in_1_port, B(0) => 
                           WB_in_0_port, SEL => FWDB2_SEL, Y(31) => 
                           B2_MUX_out_31_port, Y(30) => B2_MUX_out_30_port, 
                           Y(29) => B2_MUX_out_29_port, Y(28) => 
                           B2_MUX_out_28_port, Y(27) => B2_MUX_out_27_port, 
                           Y(26) => B2_MUX_out_26_port, Y(25) => 
                           B2_MUX_out_25_port, Y(24) => B2_MUX_out_24_port, 
                           Y(23) => B2_MUX_out_23_port, Y(22) => 
                           B2_MUX_out_22_port, Y(21) => B2_MUX_out_21_port, 
                           Y(20) => B2_MUX_out_20_port, Y(19) => 
                           B2_MUX_out_19_port, Y(18) => B2_MUX_out_18_port, 
                           Y(17) => B2_MUX_out_17_port, Y(16) => 
                           B2_MUX_out_16_port, Y(15) => B2_MUX_out_15_port, 
                           Y(14) => B2_MUX_out_14_port, Y(13) => 
                           B2_MUX_out_13_port, Y(12) => B2_MUX_out_12_port, 
                           Y(11) => B2_MUX_out_11_port, Y(10) => 
                           B2_MUX_out_10_port, Y(9) => B2_MUX_out_9_port, Y(8) 
                           => B2_MUX_out_8_port, Y(7) => B2_MUX_out_7_port, 
                           Y(6) => B2_MUX_out_6_port, Y(5) => B2_MUX_out_5_port
                           , Y(4) => B2_MUX_out_4_port, Y(3) => 
                           B2_MUX_out_3_port, Y(2) => B2_MUX_out_2_port, Y(1) 
                           => B2_MUX_out_1_port, Y(0) => B2_MUX_out_0_port);
   WBMUX : MUX2to1_NBIT32_1 port map( A(31) => ALR2_out_31_port, A(30) => 
                           ALR2_out_30_port, A(29) => ALR2_out_29_port, A(28) 
                           => ALR2_out_28_port, A(27) => ALR2_out_27_port, 
                           A(26) => ALR2_out_26_port, A(25) => ALR2_out_25_port
                           , A(24) => ALR2_out_24_port, A(23) => 
                           ALR2_out_23_port, A(22) => ALR2_out_22_port, A(21) 
                           => ALR2_out_21_port, A(20) => ALR2_out_20_port, 
                           A(19) => ALR2_out_19_port, A(18) => ALR2_out_18_port
                           , A(17) => ALR2_out_17_port, A(16) => 
                           ALR2_out_16_port, A(15) => ALR2_out_15_port, A(14) 
                           => ALR2_out_14_port, A(13) => ALR2_out_13_port, 
                           A(12) => ALR2_out_12_port, A(11) => ALR2_out_11_port
                           , A(10) => ALR2_out_10_port, A(9) => ALR2_out_9_port
                           , A(8) => ALR2_out_8_port, A(7) => ALR2_out_7_port, 
                           A(6) => ALR2_out_6_port, A(5) => ALR2_out_5_port, 
                           A(4) => ALR2_out_4_port, A(3) => ALR2_out_3_port, 
                           A(2) => ALR2_out_2_port, A(1) => ALR2_out_1_port, 
                           A(0) => ALR2_out_0_port, B(31) => LMD_out_31_port, 
                           B(30) => LMD_out_30_port, B(29) => LMD_out_29_port, 
                           B(28) => LMD_out_28_port, B(27) => LMD_out_27_port, 
                           B(26) => LMD_out_26_port, B(25) => LMD_out_25_port, 
                           B(24) => LMD_out_24_port, B(23) => LMD_out_23_port, 
                           B(22) => LMD_out_22_port, B(21) => LMD_out_21_port, 
                           B(20) => LMD_out_20_port, B(19) => LMD_out_19_port, 
                           B(18) => LMD_out_18_port, B(17) => LMD_out_17_port, 
                           B(16) => LMD_out_16_port, B(15) => LMD_out_15_port, 
                           B(14) => LMD_out_14_port, B(13) => LMD_out_13_port, 
                           B(12) => LMD_out_12_port, B(11) => LMD_out_11_port, 
                           B(10) => LMD_out_10_port, B(9) => LMD_out_9_port, 
                           B(8) => LMD_out_8_port, B(7) => LMD_out_7_port, B(6)
                           => LMD_out_6_port, B(5) => LMD_out_5_port, B(4) => 
                           LMD_out_4_port, B(3) => LMD_out_3_port, B(2) => 
                           LMD_out_2_port, B(1) => LMD_out_1_port, B(0) => 
                           LMD_out_0_port, SEL => WB_SEL, Y(31) => 
                           WB_in_31_port, Y(30) => WB_in_30_port, Y(29) => 
                           WB_in_29_port, Y(28) => WB_in_28_port, Y(27) => 
                           WB_in_27_port, Y(26) => WB_in_26_port, Y(25) => 
                           WB_in_25_port, Y(24) => WB_in_24_port, Y(23) => 
                           WB_in_23_port, Y(22) => WB_in_22_port, Y(21) => 
                           WB_in_21_port, Y(20) => WB_in_20_port, Y(19) => 
                           WB_in_19_port, Y(18) => WB_in_18_port, Y(17) => 
                           WB_in_17_port, Y(16) => WB_in_16_port, Y(15) => 
                           WB_in_15_port, Y(14) => WB_in_14_port, Y(13) => 
                           WB_in_13_port, Y(12) => WB_in_12_port, Y(11) => 
                           WB_in_11_port, Y(10) => WB_in_10_port, Y(9) => 
                           WB_in_9_port, Y(8) => WB_in_8_port, Y(7) => 
                           WB_in_7_port, Y(6) => WB_in_6_port, Y(5) => 
                           WB_in_5_port, Y(4) => WB_in_4_port, Y(3) => 
                           WB_in_3_port, Y(2) => WB_in_2_port, Y(1) => 
                           WB_in_1_port, Y(0) => WB_in_0_port);
   RF_MUX_ADDR : MUX3to1_NBIT5 port map( A(4) => RWB3_out_15_port, A(3) => 
                           RWB3_out_14_port, A(2) => RWB3_out_13_port, A(1) => 
                           RWB3_out_12_port, A(0) => RWB3_out_11_port, B(4) => 
                           RWB3_out_20_port, B(3) => RWB3_out_19_port, B(2) => 
                           RWB3_out_18_port, B(1) => RWB3_out_17_port, B(0) => 
                           RWB3_out_16_port, C(4) => X_Logic1_port, C(3) => 
                           X_Logic1_port, C(2) => X_Logic1_port, C(1) => 
                           X_Logic1_port, C(0) => X_Logic1_port, SEL(1) => 
                           RF_MUX_SEL(1), SEL(0) => RF_MUX_SEL(0), Y(4) => 
                           RF_MUX_out_4_port, Y(3) => RF_MUX_out_3_port, Y(2) 
                           => RF_MUX_out_2_port, Y(1) => RF_MUX_out_1_port, 
                           Y(0) => RF_MUX_out_0_port);
   ALU1 : ALU_NBIT32 port map( CLOCK => CLK, AluOpcode(0) => ALU_OPCODE(0), 
                           AluOpcode(1) => ALU_OPCODE(1), AluOpcode(2) => 
                           ALU_OPCODE(2), AluOpcode(3) => ALU_OPCODE(3), 
                           AluOpcode(4) => ALU_OPCODE(4), A(31) => A_in_31_port
                           , A(30) => A_in_30_port, A(29) => A_in_29_port, 
                           A(28) => A_in_28_port, A(27) => A_in_27_port, A(26) 
                           => A_in_26_port, A(25) => A_in_25_port, A(24) => 
                           A_in_24_port, A(23) => A_in_23_port, A(22) => 
                           A_in_22_port, A(21) => A_in_21_port, A(20) => 
                           A_in_20_port, A(19) => A_in_19_port, A(18) => 
                           A_in_18_port, A(17) => A_in_17_port, A(16) => 
                           A_in_16_port, A(15) => A_in_15_port, A(14) => 
                           A_in_14_port, A(13) => A_in_13_port, A(12) => 
                           A_in_12_port, A(11) => A_in_11_port, A(10) => 
                           A_in_10_port, A(9) => A_in_9_port, A(8) => 
                           A_in_8_port, A(7) => A_in_7_port, A(6) => 
                           A_in_6_port, A(5) => A_in_5_port, A(4) => 
                           A_in_4_port, A(3) => A_in_3_port, A(2) => 
                           A_in_2_port, A(1) => A_in_1_port, A(0) => 
                           A_in_0_port, B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Cin => PSW_out_6_port, ALU_out(31) => 
                           ALR_in_31_port, ALU_out(30) => ALR_in_30_port, 
                           ALU_out(29) => ALR_in_29_port, ALU_out(28) => 
                           ALR_in_28_port, ALU_out(27) => ALR_in_27_port, 
                           ALU_out(26) => ALR_in_26_port, ALU_out(25) => 
                           ALR_in_25_port, ALU_out(24) => ALR_in_24_port, 
                           ALU_out(23) => ALR_in_23_port, ALU_out(22) => 
                           ALR_in_22_port, ALU_out(21) => ALR_in_21_port, 
                           ALU_out(20) => ALR_in_20_port, ALU_out(19) => 
                           ALR_in_19_port, ALU_out(18) => ALR_in_18_port, 
                           ALU_out(17) => ALR_in_17_port, ALU_out(16) => 
                           ALR_in_16_port, ALU_out(15) => ALR_in_15_port, 
                           ALU_out(14) => ALR_in_14_port, ALU_out(13) => 
                           ALR_in_13_port, ALU_out(12) => ALR_in_12_port, 
                           ALU_out(11) => ALR_in_11_port, ALU_out(10) => 
                           ALR_in_10_port, ALU_out(9) => ALR_in_9_port, 
                           ALU_out(8) => ALR_in_8_port, ALU_out(7) => 
                           ALR_in_7_port, ALU_out(6) => ALR_in_6_port, 
                           ALU_out(5) => ALR_in_5_port, ALU_out(4) => 
                           ALR_in_4_port, ALU_out(3) => ALR_in_3_port, 
                           ALU_out(2) => ALR_in_2_port, ALU_out(1) => 
                           ALR_in_1_port, ALU_out(0) => ALR_in_0_port, Cout => 
                           PSW_in_6_port, COND(5) => PSW_in_5_port, COND(4) => 
                           PSW_in_4_port, COND(3) => PSW_in_3_port, COND(2) => 
                           PSW_in_2_port, COND(1) => PSW_in_1_port, COND(0) => 
                           PSW_in_0_port);
   FWD1 : FWDU_IR_SIZE32 port map( CLOCK => CLK, RESET => n23, EN => n35, 
                           IR(31) => IR_out_31_port, IR(30) => IR_out_30_port, 
                           IR(29) => IR_out_29_port, IR(28) => IR_out_28_port, 
                           IR(27) => IR_out_27_port, IR(26) => IR_out_26_port, 
                           IR(25) => IR_out_25_port, IR(24) => IR_out_24_port, 
                           IR(23) => IR_out_23_port, IR(22) => IR_out_22_port, 
                           IR(21) => IR_out_21_port, IR(20) => IR_out_20_port, 
                           IR(19) => IR_out_19_port, IR(18) => IR_out_18_port, 
                           IR(17) => IR_out_17_port, IR(16) => IR_out_16_port, 
                           IR(15) => IR_out_15_port, IR(14) => IR_out_14_port, 
                           IR(13) => IR_out_13_port, IR(12) => IR_out_12_port, 
                           IR(11) => IR_out_11_port, IR(10) => IR_out_10_port, 
                           IR(9) => IR_out_9_port, IR(8) => IR_out_8_port, 
                           IR(7) => IR_out_7_port, IR(6) => IR_out_6_port, 
                           IR(5) => IR_out_5_port, IR(4) => IR_out_4_port, 
                           IR(3) => IR_out_3_port, IR(2) => IR_out_2_port, 
                           IR(1) => IR_out_1_port, IR(0) => IR_out_0_port, 
                           FWD_A(1) => FWDA_SEL_1_port, FWD_A(0) => 
                           FWDA_SEL_0_port, FWD_B(1) => FWDB_SEL_1_port, 
                           FWD_B(0) => FWDB_SEL_0_port, FWD_B2 => FWDB2_SEL, 
                           ZDU_SEL(1) => ZDU_SEL_1_port, ZDU_SEL(0) => 
                           ZDU_SEL_0_port);
   HDU1 : HDU_IR_SIZE32 port map( clk => CLK, rst => n23, IR(31) => 
                           IR_out_31_port, IR(30) => IR_out_30_port, IR(29) => 
                           IR_out_29_port, IR(28) => IR_out_28_port, IR(27) => 
                           IR_out_27_port, IR(26) => IR_out_26_port, IR(25) => 
                           IR_out_25_port, IR(24) => IR_out_24_port, IR(23) => 
                           IR_out_23_port, IR(22) => IR_out_22_port, IR(21) => 
                           IR_out_21_port, IR(20) => IR_out_20_port, IR(19) => 
                           IR_out_19_port, IR(18) => IR_out_18_port, IR(17) => 
                           IR_out_17_port, IR(16) => IR_out_16_port, IR(15) => 
                           IR_out_15_port, IR(14) => IR_out_14_port, IR(13) => 
                           IR_out_13_port, IR(12) => IR_out_12_port, IR(11) => 
                           IR_out_11_port, IR(10) => IR_out_10_port, IR(9) => 
                           IR_out_9_port, IR(8) => IR_out_8_port, IR(7) => 
                           IR_out_7_port, IR(6) => IR_out_6_port, IR(5) => 
                           IR_out_5_port, IR(4) => IR_out_4_port, IR(3) => 
                           IR_out_3_port, IR(2) => IR_out_2_port, IR(1) => 
                           IR_out_1_port, IR(0) => IR_out_0_port, STALL_CODE(1)
                           => STALL(1), STALL_CODE(0) => STALL(0), IF_STALL => 
                           IF_STALL, ID_STALL => ID_STALL, EX_STALL => EX_STALL
                           , MEM_STALL => MEM_STALL, WB_STALL => n_1792);
   BHT1 : BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 port map( clock => CLK, rst => n24
                           , address(31) => BHT_in_31_port, address(30) => 
                           BHT_in_30_port, address(29) => BHT_in_29_port, 
                           address(28) => BHT_in_28_port, address(27) => 
                           BHT_in_27_port, address(26) => BHT_in_26_port, 
                           address(25) => BHT_in_25_port, address(24) => 
                           BHT_in_24_port, address(23) => BHT_in_23_port, 
                           address(22) => BHT_in_22_port, address(21) => 
                           BHT_in_21_port, address(20) => BHT_in_20_port, 
                           address(19) => BHT_in_19_port, address(18) => 
                           BHT_in_18_port, address(17) => BHT_in_17_port, 
                           address(16) => BHT_in_16_port, address(15) => 
                           BHT_in_15_port, address(14) => BHT_in_14_port, 
                           address(13) => BHT_in_13_port, address(12) => 
                           BHT_in_12_port, address(11) => BHT_in_11_port, 
                           address(10) => BHT_in_10_port, address(9) => 
                           BHT_in_9_port, address(8) => BHT_in_8_port, 
                           address(7) => BHT_in_7_port, address(6) => 
                           BHT_in_6_port, address(5) => BHT_in_5_port, 
                           address(4) => BHT_in_4_port, address(3) => 
                           BHT_in_3_port, address(2) => BHT_in_2_port, 
                           address(1) => BHT_in_1_port, address(0) => 
                           BHT_in_0_port, d_in => ZDU_out, w_en => n7, d_out =>
                           BHT_out);
   CWBU1 : CWBU port map( CLOCK => CLK, ALU_OP(0) => ALU_OPCODE(0), ALU_OP(1) 
                           => ALU_OPCODE(1), ALU_OP(2) => ALU_OPCODE(2), 
                           ALU_OP(3) => ALU_OPCODE(3), ALU_OP(4) => 
                           ALU_OPCODE(4), PSW(6) => PSW_out_6_port, PSW(5) => 
                           PSW_out_5_port, PSW(4) => PSW_out_4_port, PSW(3) => 
                           PSW_out_3_port, PSW(2) => PSW_out_2_port, PSW(1) => 
                           PSW_out_1_port, PSW(0) => PSW_out_0_port, 
                           COND_SEL(1) => CWB_out_1_port, COND_SEL(0) => 
                           CWB_out_0_port, CWB_SEL(1) => CWB_SEL(1), CWB_SEL(0)
                           => CWB_SEL(0), CWB_MUW_SEL(1) => CWB_MUX_SEL_1_port,
                           CWB_MUW_SEL(0) => CWB_MUX_SEL_0_port);
   RF1 : RF_NBIT32_NREG32 port map( CLK => CLK, RESET => n23, ENABLE => 
                           X_Logic1_port, RD1 => n4, RD2 => n4, WR => RF_WR, 
                           ADD_WR(4) => RF_MUX_out_4_port, ADD_WR(3) => 
                           RF_MUX_out_3_port, ADD_WR(2) => RF_MUX_out_2_port, 
                           ADD_WR(1) => RF_MUX_out_1_port, ADD_WR(0) => 
                           RF_MUX_out_0_port, ADD_RD1(4) => IR_out_25_port, 
                           ADD_RD1(3) => IR_out_24_port, ADD_RD1(2) => 
                           IR_out_23_port, ADD_RD1(1) => IR_out_22_port, 
                           ADD_RD1(0) => IR_out_21_port, ADD_RD2(4) => 
                           IR_out_20_port, ADD_RD2(3) => IR_out_19_port, 
                           ADD_RD2(2) => IR_out_18_port, ADD_RD2(1) => 
                           IR_out_17_port, ADD_RD2(0) => IR_out_16_port, 
                           DATAIN(31) => WB_in_31_port, DATAIN(30) => 
                           WB_in_30_port, DATAIN(29) => WB_in_29_port, 
                           DATAIN(28) => WB_in_28_port, DATAIN(27) => 
                           WB_in_27_port, DATAIN(26) => WB_in_26_port, 
                           DATAIN(25) => WB_in_25_port, DATAIN(24) => 
                           WB_in_24_port, DATAIN(23) => WB_in_23_port, 
                           DATAIN(22) => WB_in_22_port, DATAIN(21) => 
                           WB_in_21_port, DATAIN(20) => WB_in_20_port, 
                           DATAIN(19) => WB_in_19_port, DATAIN(18) => 
                           WB_in_18_port, DATAIN(17) => WB_in_17_port, 
                           DATAIN(16) => WB_in_16_port, DATAIN(15) => 
                           WB_in_15_port, DATAIN(14) => WB_in_14_port, 
                           DATAIN(13) => WB_in_13_port, DATAIN(12) => 
                           WB_in_12_port, DATAIN(11) => WB_in_11_port, 
                           DATAIN(10) => WB_in_10_port, DATAIN(9) => 
                           WB_in_9_port, DATAIN(8) => WB_in_8_port, DATAIN(7) 
                           => WB_in_7_port, DATAIN(6) => WB_in_6_port, 
                           DATAIN(5) => WB_in_5_port, DATAIN(4) => WB_in_4_port
                           , DATAIN(3) => WB_in_3_port, DATAIN(2) => 
                           WB_in_2_port, DATAIN(1) => WB_in_1_port, DATAIN(0) 
                           => WB_in_0_port, OUT1(31) => RA_out_31_port, 
                           OUT1(30) => RA_out_30_port, OUT1(29) => 
                           RA_out_29_port, OUT1(28) => RA_out_28_port, OUT1(27)
                           => RA_out_27_port, OUT1(26) => RA_out_26_port, 
                           OUT1(25) => RA_out_25_port, OUT1(24) => 
                           RA_out_24_port, OUT1(23) => RA_out_23_port, OUT1(22)
                           => RA_out_22_port, OUT1(21) => RA_out_21_port, 
                           OUT1(20) => RA_out_20_port, OUT1(19) => 
                           RA_out_19_port, OUT1(18) => RA_out_18_port, OUT1(17)
                           => RA_out_17_port, OUT1(16) => RA_out_16_port, 
                           OUT1(15) => RA_out_15_port, OUT1(14) => 
                           RA_out_14_port, OUT1(13) => RA_out_13_port, OUT1(12)
                           => RA_out_12_port, OUT1(11) => RA_out_11_port, 
                           OUT1(10) => RA_out_10_port, OUT1(9) => RA_out_9_port
                           , OUT1(8) => RA_out_8_port, OUT1(7) => RA_out_7_port
                           , OUT1(6) => RA_out_6_port, OUT1(5) => RA_out_5_port
                           , OUT1(4) => RA_out_4_port, OUT1(3) => RA_out_3_port
                           , OUT1(2) => RA_out_2_port, OUT1(1) => RA_out_1_port
                           , OUT1(0) => RA_out_0_port, OUT2(31) => 
                           RB_out_31_port, OUT2(30) => RB_out_30_port, OUT2(29)
                           => RB_out_29_port, OUT2(28) => RB_out_28_port, 
                           OUT2(27) => RB_out_27_port, OUT2(26) => 
                           RB_out_26_port, OUT2(25) => RB_out_25_port, OUT2(24)
                           => RB_out_24_port, OUT2(23) => RB_out_23_port, 
                           OUT2(22) => RB_out_22_port, OUT2(21) => 
                           RB_out_21_port, OUT2(20) => RB_out_20_port, OUT2(19)
                           => RB_out_19_port, OUT2(18) => RB_out_18_port, 
                           OUT2(17) => RB_out_17_port, OUT2(16) => 
                           RB_out_16_port, OUT2(15) => RB_out_15_port, OUT2(14)
                           => RB_out_14_port, OUT2(13) => RB_out_13_port, 
                           OUT2(12) => RB_out_12_port, OUT2(11) => 
                           RB_out_11_port, OUT2(10) => RB_out_10_port, OUT2(9) 
                           => RB_out_9_port, OUT2(8) => RB_out_8_port, OUT2(7) 
                           => RB_out_7_port, OUT2(6) => RB_out_6_port, OUT2(5) 
                           => RB_out_5_port, OUT2(4) => RB_out_4_port, OUT2(3) 
                           => RB_out_3_port, OUT2(2) => RB_out_2_port, OUT2(1) 
                           => RB_out_1_port, OUT2(0) => RB_out_0_port);
   U3 : NOR2_X2 port map( A1 => n30, A2 => n29, ZN => IRAMMUX_SEL);
   U4 : AND4_X1 port map( A1 => n15, A2 => n16, A3 => n13, A4 => n14_port, ZN 
                           => n28);
   U5 : AND2_X1 port map( A1 => ID_EN, A2 => n35, ZN => n1);
   U6 : CLKBUF_X1 port map( A => n31, Z => n2);
   U7 : BUF_X1 port map( A => n22, Z => n24);
   U8 : BUF_X1 port map( A => n22, Z => n23);
   U9 : BUF_X1 port map( A => n9, Z => n20);
   U10 : BUF_X1 port map( A => MEM_ENABLE, Z => n5);
   U11 : BUF_X1 port map( A => EX_ENABLE, Z => n6);
   U12 : BUF_X1 port map( A => n20, Z => n11);
   U13 : BUF_X1 port map( A => n20, Z => n12);
   U14 : BUF_X1 port map( A => n20, Z => n19);
   U15 : INV_X1 port map( A => n8, ZN => n7);
   U16 : BUF_X1 port map( A => n21, Z => n10);
   U17 : BUF_X1 port map( A => n9, Z => n21);
   U18 : INV_X1 port map( A => BPR_EN2, ZN => n8);
   U19 : XNOR2_X1 port map( A => n3, B => RWB1_out_26_port, ZN => n31);
   U20 : AND4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => n3
                           );
   U21 : NOR2_X1 port map( A1 => MEM_STALL, A2 => n37, ZN => MEM_ENABLE);
   U22 : INV_X1 port map( A => MEM_EN, ZN => n37);
   U23 : OR4_X1 port map( A1 => ZDU_MUX_out_13_port, A2 => ZDU_MUX_out_12_port,
                           A3 => ZDU_MUX_out_15_port, A4 => ZDU_MUX_out_14_port
                           , ZN => n17);
   U24 : NOR4_X1 port map( A1 => ZDU_MUX_out_2_port, A2 => ZDU_MUX_out_29_port,
                           A3 => ZDU_MUX_out_28_port, A4 => ZDU_MUX_out_27_port
                           , ZN => n14_port);
   U25 : NOR4_X1 port map( A1 => ZDU_MUX_out_26_port, A2 => ZDU_MUX_out_25_port
                           , A3 => ZDU_MUX_out_24_port, A4 => 
                           ZDU_MUX_out_23_port, ZN => n13);
   U26 : NOR4_X1 port map( A1 => ZDU_MUX_out_9_port, A2 => ZDU_MUX_out_8_port, 
                           A3 => ZDU_MUX_out_7_port, A4 => ZDU_MUX_out_6_port, 
                           ZN => n16);
   U27 : NOR4_X1 port map( A1 => ZDU_MUX_out_5_port, A2 => ZDU_MUX_out_4_port, 
                           A3 => ZDU_MUX_out_3_port, A4 => ZDU_MUX_out_30_port,
                           ZN => n15);
   U28 : AND2_X1 port map( A1 => SIGND, A2 => IR_out_15_port, ZN => N14);
   U29 : NOR2_X1 port map( A1 => EX_STALL, A2 => n36, ZN => EX_ENABLE);
   U30 : INV_X1 port map( A => EX_EN, ZN => n36);
   U31 : INV_X1 port map( A => n18, ZN => n34);
   U32 : AOI21_X1 port map( B1 => BPR_EN, B2 => BHT_out, A => UCB_EN, ZN => n18
                           );
   U33 : AND2_X1 port map( A1 => RF_RD, A2 => n35, ZN => n4);
   U34 : BUF_X1 port map( A => DATA_IN(7), Z => n9);
   U35 : BUF_X1 port map( A => RST, Z => n22);
   U36 : NOR4_X1 port map( A1 => ZDU_MUX_out_19_port, A2 => ZDU_MUX_out_20_port
                           , A3 => ZDU_MUX_out_21_port, A4 => 
                           ZDU_MUX_out_22_port, ZN => n27);
   U37 : NOR4_X1 port map( A1 => ZDU_MUX_out_11_port, A2 => ZDU_MUX_out_16_port
                           , A3 => ZDU_MUX_out_17_port, A4 => 
                           ZDU_MUX_out_18_port, ZN => n26);
   U38 : NOR4_X1 port map( A1 => n17, A2 => ZDU_MUX_out_0_port, A3 => 
                           ZDU_MUX_out_1_port, A4 => ZDU_MUX_out_10_port, ZN =>
                           n25);
   U39 : INV_X1 port map( A => n2, ZN => ZDU_out);
   U40 : INV_X1 port map( A => ID_STALL, ZN => n35);
   U41 : INV_X1 port map( A => BMP, ZN => n30);
   U42 : INV_X1 port map( A => PRD_OUT, ZN => n29);
   U43 : INV_X1 port map( A => IF_STALL, ZN => n33);
   U44 : NOR3_X1 port map( A1 => n34, A2 => PRD_OUT, A3 => n30, ZN => 
                           PC_SEL_1_port);
   U45 : XOR2_X1 port map( A => n31, B => PRD_OUT, Z => n32);
   U46 : NOR2_X1 port map( A1 => n32, A2 => n8, ZN => BMP);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26 is

   port( Clk, Rst : in std_logic;  STALL : in std_logic_vector (1 downto 0);  
         IR_IN : in std_logic_vector (31 downto 0);  BMP : in std_logic;  ID_EN
         , RF_RD, SIGND, IMM_SEL, BPR_EN, UCB_EN : out std_logic;  ALU_OPCODE :
         out std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, ALUB_SEL, MEM_EN, 
         MEM_DATA_SEL, MEM_RD, MEM_WR, CS, MEM_BLC0, MEM_BLC1, LD_SEL0, LD_SEL1
         , LD_SEL2, ALR2_SEL, CWB_SEL0, CWB_SEL1, WB_SEL, RF_WR, RF_MUX_SEL0, 
         RF_MUX_SEL1 : out std_logic);

end CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26;

architecture SYN_dlx_cu_hw of 
   CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal ALU_OPCODE_3_port, ALU_OPCODE_0_port, MEM_EN_port, MEM_DATA_SEL_port,
      MEM_RD_port, MEM_WR_port, CS_port, MEM_BLC0_port, MEM_BLC1_port, 
      LD_SEL0_port, LD_SEL1_port, LD_SEL2_port, ALR2_SEL_port, CWB_SEL0_port, 
      CWB_SEL1_port, WB_SEL_port, RF_WR_port, RF_MUX_SEL0_port, 
      RF_MUX_SEL1_port, cw3_16_port, cw3_15_port, cw3_14_port, cw3_13_port, 
      cw3_12_port, cw3_11_port, cw3_10_port, cw3_9_port, cw3_8_port, cw3_7_port
      , cw3_6_port, cw3_5_port, cw3_4_port, cw3_3_port, cw3_2_port, cw3_1_port,
      cw3_0_port, cw4_3_port, cw4_2_port, cw4_1_port, cw4_0_port, 
      aluOpcode1_4_port, aluOpcode1_3_port, aluOpcode1_2_port, 
      aluOpcode1_1_port, aluOpcode1_0_port, n2, n3, n4, n5, n6, n10, n12, n14, 
      n16, n18, n20, n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44
      , n45, n46, n47, n48, n49, n51, n52, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n108, n109, n110, n115, n116,
      n117, n121, n123, n124, n125, n126, n127, n135, n136, n137, n138, n139, 
      n140, n141, n143, n146, n189, n190, n192, n1, n7, n8, ALU_OPCODE_4_port, 
      ALU_OPCODE_2_port, ALU_OPCODE_1_port, n15, n19, n21, n23, n25, n27, n29, 
      n31, n33, n35, n37, n39, n41, n43, n50, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n104, n105, n106, n107, n111, n112, n113, n114, n118, n119, n120, n122,
      n128, n129, n130, n131, n132, n133, n134, n142, n144, n145, n147, n148, 
      n149, n150, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, 
      n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, 
      n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, 
      n_1818 : std_logic;

begin
   ALU_OPCODE <= ( ALU_OPCODE_4_port, ALU_OPCODE_3_port, ALU_OPCODE_2_port, 
      ALU_OPCODE_1_port, ALU_OPCODE_0_port );
   MEM_EN <= MEM_EN_port;
   MEM_DATA_SEL <= MEM_DATA_SEL_port;
   MEM_RD <= MEM_RD_port;
   MEM_WR <= MEM_WR_port;
   CS <= CS_port;
   MEM_BLC0 <= MEM_BLC0_port;
   MEM_BLC1 <= MEM_BLC1_port;
   LD_SEL0 <= LD_SEL0_port;
   LD_SEL1 <= LD_SEL1_port;
   LD_SEL2 <= LD_SEL2_port;
   ALR2_SEL <= ALR2_SEL_port;
   CWB_SEL0 <= CWB_SEL0_port;
   CWB_SEL1 <= CWB_SEL1_port;
   WB_SEL <= WB_SEL_port;
   RF_WR <= RF_WR_port;
   RF_MUX_SEL0 <= RF_MUX_SEL0_port;
   RF_MUX_SEL1 <= RF_MUX_SEL1_port;
   
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => n192, CK => Clk, RN => n19, Q
                           => aluOpcode1_4_port, QN => n48);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => n190, CK => Clk, RN => n19, Q
                           => aluOpcode1_1_port, QN => n51);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => n189, CK => Clk, RN => n19, Q
                           => aluOpcode1_0_port, QN => n52);
   UCB_EN <= '0';
   BPR_EN <= '0';
   IMM_SEL <= '0';
   SIGND <= '0';
   RF_RD <= '0';
   ID_EN <= '0';
   cw4_reg_16_inst : DFFR_X1 port map( D => n10, CK => Clk, RN => n23, Q => 
                           MEM_EN_port, QN => n_1793);
   cw4_reg_15_inst : DFFR_X1 port map( D => n12, CK => Clk, RN => n23, Q => 
                           MEM_DATA_SEL_port, QN => n_1794);
   cw4_reg_14_inst : DFFR_X1 port map( D => n14, CK => Clk, RN => n23, Q => 
                           MEM_RD_port, QN => n_1795);
   cw4_reg_13_inst : DFFR_X1 port map( D => n16, CK => Clk, RN => n23, Q => 
                           MEM_WR_port, QN => n_1796);
   cw4_reg_12_inst : DFFR_X1 port map( D => n18, CK => Clk, RN => n23, Q => 
                           CS_port, QN => n_1797);
   cw4_reg_11_inst : DFFR_X1 port map( D => n20, CK => Clk, RN => n23, Q => 
                           MEM_BLC0_port, QN => n_1798);
   cw4_reg_10_inst : DFFR_X1 port map( D => n22, CK => Clk, RN => n23, Q => 
                           MEM_BLC1_port, QN => n_1799);
   cw4_reg_9_inst : DFFR_X1 port map( D => n24, CK => Clk, RN => n23, Q => 
                           LD_SEL0_port, QN => n_1800);
   cw4_reg_8_inst : DFFR_X1 port map( D => n26, CK => Clk, RN => n23, Q => 
                           LD_SEL1_port, QN => n_1801);
   cw4_reg_7_inst : DFFR_X1 port map( D => n28, CK => Clk, RN => n23, Q => 
                           LD_SEL2_port, QN => n_1802);
   cw4_reg_6_inst : DFFR_X1 port map( D => n30, CK => Clk, RN => n23, Q => 
                           ALR2_SEL_port, QN => n_1803);
   cw4_reg_5_inst : DFFR_X1 port map( D => n32, CK => Clk, RN => n23, Q => 
                           CWB_SEL0_port, QN => n_1804);
   cw4_reg_4_inst : DFFR_X1 port map( D => n34, CK => Clk, RN => n23, Q => 
                           CWB_SEL1_port, QN => n_1805);
   cw4_reg_3_inst : DFFR_X1 port map( D => n36, CK => Clk, RN => n23, Q => 
                           cw4_3_port, QN => n_1806);
   cw4_reg_2_inst : DFFR_X1 port map( D => n38, CK => Clk, RN => n23, Q => 
                           cw4_2_port, QN => n_1807);
   cw4_reg_1_inst : DFFR_X1 port map( D => n40, CK => Clk, RN => n23, Q => 
                           cw4_1_port, QN => n_1808);
   cw4_reg_0_inst : DFFR_X1 port map( D => n42, CK => Clk, RN => n23, Q => 
                           cw4_0_port, QN => n_1809);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => n49, CK => Clk, RN => n23, Q 
                           => aluOpcode1_3_port, QN => n113);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => n7, CK => Clk, RN => n23, Q 
                           => aluOpcode1_2_port, QN => n_1810);
   cw5_reg_3_inst : DFFR_X1 port map( D => n44, CK => Clk, RN => n23, Q => 
                           WB_SEL_port, QN => n_1811);
   cw5_reg_2_inst : DFFR_X1 port map( D => n45, CK => Clk, RN => n23, Q => 
                           RF_WR_port, QN => n_1812);
   cw5_reg_1_inst : DFFR_X1 port map( D => n46, CK => Clk, RN => n23, Q => 
                           RF_MUX_SEL0_port, QN => n_1813);
   cw5_reg_0_inst : DFFR_X1 port map( D => n47, CK => Clk, RN => n23, Q => 
                           RF_MUX_SEL1_port, QN => n_1814);
   aluOpcode2_reg_3_inst : DFFR_X2 port map( D => n3, CK => Clk, RN => n23, Q 
                           => ALU_OPCODE_3_port, QN => n112);
   aluOpcode2_reg_2_inst : DFFR_X2 port map( D => n4, CK => Clk, RN => n23, Q 
                           => ALU_OPCODE_2_port, QN => n_1815);
   aluOpcode2_reg_1_inst : DFFR_X2 port map( D => n5, CK => Clk, RN => n23, Q 
                           => ALU_OPCODE_1_port, QN => n_1816);
   aluOpcode2_reg_0_inst : DFFR_X2 port map( D => n6, CK => Clk, RN => n23, Q 
                           => ALU_OPCODE_0_port, QN => n_1817);
   aluOpcode2_reg_4_inst : DFFR_X2 port map( D => n2, CK => Clk, RN => n23, Q 
                           => ALU_OPCODE_4_port, QN => n_1818);
   U3 : MUX2_X1 port map( A => cw3_15_port, B => MEM_DATA_SEL_port, S => n1, Z 
                           => n12);
   U4 : MUX2_X1 port map( A => cw3_14_port, B => MEM_RD_port, S => n1, Z => n14
                           );
   U5 : MUX2_X1 port map( A => cw3_10_port, B => MEM_BLC1_port, S => n1, Z => 
                           n22);
   U6 : MUX2_X1 port map( A => cw3_9_port, B => LD_SEL0_port, S => n1, Z => n24
                           );
   U7 : MUX2_X1 port map( A => cw3_6_port, B => ALR2_SEL_port, S => n1, Z => 
                           n30);
   U8 : MUX2_X1 port map( A => cw3_5_port, B => CWB_SEL0_port, S => n1, Z => 
                           n32);
   U9 : MUX2_X1 port map( A => cw3_2_port, B => cw4_2_port, S => n1, Z => n38);
   U10 : MUX2_X1 port map( A => cw3_1_port, B => cw4_1_port, S => n1, Z => n40)
                           ;
   U11 : MUX2_X1 port map( A => cw3_12_port, B => CS_port, S => n1, Z => n18);
   U12 : MUX2_X1 port map( A => cw3_16_port, B => MEM_EN_port, S => n1, Z => 
                           n10);
   U13 : MUX2_X1 port map( A => cw3_13_port, B => MEM_WR_port, S => n1, Z => 
                           n16);
   U14 : MUX2_X1 port map( A => cw3_11_port, B => MEM_BLC0_port, S => n1, Z => 
                           n20);
   U15 : MUX2_X1 port map( A => cw3_8_port, B => LD_SEL1_port, S => n1, Z => 
                           n26);
   U16 : MUX2_X1 port map( A => cw3_7_port, B => LD_SEL2_port, S => n1, Z => 
                           n28);
   U17 : MUX2_X1 port map( A => cw3_4_port, B => CWB_SEL1_port, S => n1, Z => 
                           n34);
   U18 : MUX2_X1 port map( A => cw3_3_port, B => cw4_3_port, S => n1, Z => n36)
                           ;
   U19 : MUX2_X1 port map( A => cw3_0_port, B => cw4_0_port, S => n1, Z => n42)
                           ;
   U20 : INV_X2 port map( A => Rst, ZN => n23);
   U21 : BUF_X1 port map( A => n129, Z => n15);
   U22 : OAI22_X1 port map( A1 => n101, A2 => n136, B1 => n27, B2 => n100, ZN 
                           => n126);
   U23 : BUF_X1 port map( A => n21, Z => n19);
   U30 : AND2_X2 port map( A1 => STALL(1), A2 => n60, ZN => n1);
   U31 : NAND2_X1 port map( A1 => n149, A2 => n150, ZN => n101);
   U32 : NAND2_X1 port map( A1 => n133, A2 => n134, ZN => n110);
   U33 : NOR2_X1 port map( A1 => n97, A2 => n137, ZN => n116);
   U34 : NOR4_X1 port map( A1 => n101, A2 => n145, A3 => n147, A4 => n148, ZN 
                           => n137);
   U35 : NAND2_X1 port map( A1 => n140, A2 => n148, ZN => n100);
   U36 : NOR2_X1 port map( A1 => n124, A2 => n110, ZN => n93);
   U37 : NOR2_X1 port map( A1 => n132, A2 => n110, ZN => n92);
   U38 : INV_X1 port map( A => n103, ZN => n144);
   U39 : NAND2_X1 port map( A1 => n141, A2 => n147, ZN => n136);
   U40 : OR2_X1 port map( A1 => n90, A2 => n109, ZN => n123);
   U41 : BUF_X1 port map( A => n23, Z => n21);
   U42 : MUX2_X1 port map( A => n8, B => aluOpcode1_2_port, S => n122, Z => n7)
                           ;
   U43 : OR4_X1 port map( A1 => n84, A2 => n83, A3 => n82, A4 => n81, ZN => n8)
                           ;
   U44 : NOR4_X1 port map( A1 => n145, A2 => n147, A3 => IR_IN(2), A4 => 
                           IR_IN(4), ZN => n103);
   U45 : NOR4_X1 port map( A1 => n133, A2 => n134, A3 => IR_IN(29), A4 => 
                           IR_IN(31), ZN => n91);
   U46 : OAI222_X1 port map( A1 => IR_IN(1), A2 => n98, B1 => n99, B2 => n150, 
                           C1 => n100, C2 => n101, ZN => n96);
   U47 : AOI21_X1 port map( B1 => n102, B2 => IR_IN(1), A => n103, ZN => n99);
   U48 : NOR2_X1 port map( A1 => n149, A2 => IR_IN(0), ZN => n95);
   U49 : NOR3_X1 port map( A1 => n147, A2 => IR_IN(2), A3 => n145, ZN => n102);
   U50 : NOR3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(4), A3 => n145, ZN => 
                           n140);
   U51 : NOR3_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), A3 => n148, ZN => 
                           n141);
   U52 : AOI211_X1 port map( C1 => n130, C2 => IR_IN(1), A => n125, B => n126, 
                           ZN => n121);
   U53 : OAI22_X1 port map( A1 => IR_IN(1), A2 => n144, B1 => n127, B2 => n98, 
                           ZN => n125);
   U54 : AOI21_X1 port map( B1 => IR_IN(0), B2 => n149, A => n95, ZN => n127);
   U55 : NOR3_X1 port map( A1 => n132, A2 => IR_IN(30), A3 => IR_IN(29), ZN => 
                           n94);
   U56 : NOR3_X1 port map( A1 => n124, A2 => IR_IN(28), A3 => n133, ZN => n89);
   U57 : NOR2_X1 port map( A1 => n131, A2 => IR_IN(26), ZN => n90);
   U58 : INV_X1 port map( A => IR_IN(5), ZN => n145);
   U59 : OAI21_X1 port map( B1 => n27, B2 => n98, A => n138, ZN => n97);
   U60 : NAND4_X1 port map( A1 => IR_IN(2), A2 => n149, A3 => IR_IN(3), A4 => 
                           n139, ZN => n138);
   U61 : NOR2_X1 port map( A1 => n150, A2 => n145, ZN => n139);
   U62 : INV_X1 port map( A => IR_IN(1), ZN => n149);
   U63 : NAND2_X1 port map( A1 => n140, A2 => IR_IN(2), ZN => n98);
   U64 : NOR3_X1 port map( A1 => n110, A2 => IR_IN(31), A3 => IR_IN(29), ZN => 
                           n143);
   U65 : INV_X1 port map( A => IR_IN(3), ZN => n147);
   U66 : OAI211_X1 port map( C1 => n101, C2 => n98, A => n142, B => n116, ZN =>
                           n115);
   U67 : INV_X1 port map( A => n117, ZN => n142);
   U68 : OAI22_X1 port map( A1 => n149, A2 => n100, B1 => IR_IN(1), B2 => n144,
                           ZN => n117);
   U69 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n132, ZN => n124);
   U70 : INV_X1 port map( A => IR_IN(2), ZN => n148);
   U71 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n146);
   U72 : INV_X1 port map( A => IR_IN(31), ZN => n132);
   U73 : INV_X1 port map( A => IR_IN(30), ZN => n133);
   U74 : INV_X1 port map( A => IR_IN(0), ZN => n150);
   U75 : AOI22_X1 port map( A1 => n102, A2 => IR_IN(1), B1 => n130, B2 => n95, 
                           ZN => n135);
   U76 : AND3_X1 port map( A1 => IR_IN(29), A2 => n134, A3 => IR_IN(30), ZN => 
                           n108);
   U77 : AND2_X1 port map( A1 => IR_IN(27), A2 => IR_IN(26), ZN => n109);
   cw3_0_port <= '0';
   cw3_3_port <= '0';
   cw3_4_port <= '0';
   cw3_7_port <= '0';
   cw3_8_port <= '0';
   cw3_11_port <= '0';
   cw3_13_port <= '0';
   cw3_16_port <= '0';
   ALUB_SEL <= '0';
   ALUA_SEL <= '0';
   cw3_12_port <= '0';
   cw3_1_port <= '0';
   cw3_2_port <= '0';
   cw3_5_port <= '0';
   cw3_6_port <= '0';
   cw3_9_port <= '0';
   cw3_10_port <= '0';
   cw3_14_port <= '0';
   cw3_15_port <= '0';
   EX_EN <= '0';
   U98 : INV_X1 port map( A => BMP, ZN => n60);
   U99 : OAI21_X1 port map( B1 => STALL(1), B2 => STALL(0), A => n60, ZN => 
                           n129);
   U100 : MUX2_X1 port map( A => cw4_0_port, B => RF_MUX_SEL1_port, S => n1, Z 
                           => n47);
   U101 : MUX2_X1 port map( A => cw4_1_port, B => RF_MUX_SEL0_port, S => n1, Z 
                           => n46);
   U102 : MUX2_X1 port map( A => cw4_2_port, B => RF_WR_port, S => n1, Z => n45
                           );
   U103 : MUX2_X1 port map( A => cw4_3_port, B => WB_SEL_port, S => n1, Z => 
                           n44);
   U104 : INV_X1 port map( A => n124, ZN => n25);
   U105 : NAND3_X1 port map( A1 => IR_IN(28), A2 => n133, A3 => n25, ZN => n75)
                           ;
   U106 : INV_X1 port map( A => IR_IN(27), ZN => n131);
   U107 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n131, ZN => n76);
   U108 : INV_X1 port map( A => n141, ZN => n29);
   U109 : INV_X1 port map( A => n95, ZN => n27);
   U110 : NOR4_X1 port map( A1 => n76, A2 => n147, A3 => n29, A4 => n27, ZN => 
                           n33);
   U111 : OR3_X1 port map( A1 => IR_IN(10), A2 => n146, A3 => IR_IN(6), ZN => 
                           n50);
   U112 : NOR4_X1 port map( A1 => n110, A2 => IR_IN(31), A3 => IR_IN(29), A4 =>
                           n50, ZN => n31);
   U113 : NAND2_X1 port map( A1 => n33, A2 => n31, ZN => n118);
   U114 : NAND3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => IR_IN(28),
                           ZN => n65);
   U115 : INV_X1 port map( A => n65, ZN => n37);
   U116 : INV_X1 port map( A => n76, ZN => n35);
   U117 : OAI21_X1 port map( B1 => n89, B2 => n37, A => n35, ZN => n41);
   U118 : OAI21_X1 port map( B1 => n108, B2 => n92, A => n109, ZN => n39);
   U119 : NAND4_X1 port map( A1 => n75, A2 => n118, A3 => n41, A4 => n39, ZN =>
                           n57);
   U120 : INV_X1 port map( A => n136, ZN => n130);
   U121 : AOI211_X1 port map( C1 => n95, C2 => n130, A => n97, B => n96, ZN => 
                           n55);
   U122 : INV_X1 port map( A => IR_IN(26), ZN => n43);
   U123 : NAND2_X1 port map( A1 => n131, A2 => n43, ZN => n80);
   U124 : INV_X1 port map( A => n80, ZN => n86);
   U125 : INV_X1 port map( A => n50, ZN => n53);
   U126 : NAND3_X1 port map( A1 => n143, A2 => n86, A3 => n53, ZN => n74);
   U127 : NAND2_X1 port map( A1 => n80, A2 => n76, ZN => n68);
   U128 : INV_X1 port map( A => n68, ZN => n66);
   U129 : NOR3_X1 port map( A1 => n93, A2 => n94, A3 => n92, ZN => n54);
   U130 : OAI22_X1 port map( A1 => n55, A2 => n74, B1 => n66, B2 => n54, ZN => 
                           n56);
   U131 : AOI211_X1 port map( C1 => n91, C2 => n90, A => n57, B => n56, ZN => 
                           n58);
   U132 : INV_X1 port map( A => n129, ZN => n122);
   U133 : MUX2_X1 port map( A => n58, B => n52, S => n122, Z => n59);
   U134 : INV_X1 port map( A => n59, ZN => n189);
   U135 : NAND2_X1 port map( A1 => n15, A2 => n60, ZN => n114);
   U136 : INV_X1 port map( A => n114, ZN => n120);
   U137 : AOI22_X1 port map( A1 => ALU_OPCODE_0_port, A2 => n122, B1 => 
                           aluOpcode1_0_port, B2 => n120, ZN => n61);
   U138 : INV_X1 port map( A => n61, ZN => n6);
   U139 : INV_X1 port map( A => n74, ZN => n104);
   U140 : INV_X1 port map( A => n75, ZN => n70);
   U141 : INV_X1 port map( A => n93, ZN => n63);
   U142 : INV_X1 port map( A => n123, ZN => n79);
   U143 : INV_X1 port map( A => n90, ZN => n62);
   U144 : OAI22_X1 port map( A1 => n63, A2 => n79, B1 => n75, B2 => n62, ZN => 
                           n81);
   U145 : INV_X1 port map( A => n81, ZN => n64);
   U146 : OAI21_X1 port map( B1 => n66, B2 => n65, A => n64, ZN => n67);
   U147 : INV_X1 port map( A => n67, ZN => n107);
   U148 : NAND2_X1 port map( A1 => n89, A2 => n68, ZN => n77);
   U149 : NAND3_X1 port map( A1 => n107, A2 => n118, A3 => n77, ZN => n69);
   U150 : AOI221_X1 port map( B1 => n115, B2 => n104, C1 => n86, C2 => n70, A 
                           => n69, ZN => n71);
   U151 : MUX2_X1 port map( A => n71, B => n51, S => n122, Z => n72);
   U152 : INV_X1 port map( A => n72, ZN => n190);
   U153 : AOI22_X1 port map( A1 => ALU_OPCODE_1_port, A2 => n122, B1 => 
                           aluOpcode1_1_port, B2 => n120, ZN => n73);
   U154 : INV_X1 port map( A => n73, ZN => n5);
   U155 : OAI22_X1 port map( A1 => n76, A2 => n75, B1 => n121, B2 => n74, ZN =>
                           n84);
   U156 : INV_X1 port map( A => n77, ZN => n83);
   U157 : INV_X1 port map( A => n91, ZN => n78);
   U158 : AOI21_X1 port map( B1 => n80, B2 => n79, A => n78, ZN => n82);
   U159 : AOI22_X1 port map( A1 => ALU_OPCODE_2_port, A2 => n122, B1 => 
                           aluOpcode1_2_port, B2 => n120, ZN => n85);
   U160 : INV_X1 port map( A => n85, ZN => n4);
   U161 : OAI21_X1 port map( B1 => n90, B2 => n86, A => n91, ZN => n106);
   U162 : INV_X1 port map( A => n126, ZN => n87);
   U163 : NAND3_X1 port map( A1 => n116, A2 => n135, A3 => n87, ZN => n88);
   U164 : AOI22_X1 port map( A1 => n104, A2 => n88, B1 => n108, B2 => n123, ZN 
                           => n105);
   U165 : NAND3_X1 port map( A1 => n107, A2 => n106, A3 => n105, ZN => n111);
   U166 : MUX2_X1 port map( A => n111, B => aluOpcode1_3_port, S => n122, Z => 
                           n49);
   U167 : OAI22_X1 port map( A1 => n114, A2 => n113, B1 => n15, B2 => n112, ZN 
                           => n3);
   U168 : MUX2_X1 port map( A => n118, B => n48, S => n122, Z => n119);
   U169 : INV_X1 port map( A => n119, ZN => n192);
   U170 : AOI22_X1 port map( A1 => ALU_OPCODE_4_port, A2 => n122, B1 => 
                           aluOpcode1_4_port, B2 => n120, ZN => n128);
   U171 : INV_X1 port map( A => n128, ZN => n2);
   U172 : INV_X1 port map( A => IR_IN(28), ZN => n134);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector (31 
         downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out std_logic_vector (31 
         downto 0);  BLC : out std_logic_vector (1 downto 0);  MEM_WR, MEM_RD :
         out std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component Datapath
      port( CLK, RST : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector 
            (31 downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out 
            std_logic_vector (31 downto 0);  BMP : inout std_logic;  STALL : 
            out std_logic_vector (1 downto 0);  ID_EN, RF_RD, SIGND, IMM_SEL, 
            BPR_EN : in std_logic;  ALU_OPCODE : in std_logic_vector (0 to 4); 
            EX_EN, ALUA_SEL, ALUB_SEL, UCB_EN, MEM_EN, MEM_DATA_SEL : in 
            std_logic;  LD_SEL : in std_logic_vector (2 downto 0);  ALR2_SEL : 
            in std_logic;  CWB_SEL : in std_logic_vector (1 downto 0);  WB_SEL,
            RF_WR : in std_logic;  RF_MUX_SEL : in std_logic_vector (1 downto 
            0));
   end component;
   
   component 
      CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26
      port( Clk, Rst : in std_logic;  STALL : in std_logic_vector (1 downto 0);
            IR_IN : in std_logic_vector (31 downto 0);  BMP : in std_logic;  
            ID_EN, RF_RD, SIGND, IMM_SEL, BPR_EN, UCB_EN : out std_logic;  
            ALU_OPCODE : out std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, 
            ALUB_SEL, MEM_EN, MEM_DATA_SEL, MEM_RD, MEM_WR, CS, MEM_BLC0, 
            MEM_BLC1, LD_SEL0, LD_SEL1, LD_SEL2, ALR2_SEL, CWB_SEL0, CWB_SEL1, 
            WB_SEL, RF_WR, RF_MUX_SEL0, RF_MUX_SEL1 : out std_logic);
   end component;
   
   signal STALL_CODE_1_port, STALL_CODE_0_port, BMP_i, ID_EN_i, RF_RD_i, 
      SIGND_i, IMM_SEL_i, BPR_EN_i, UCB_EN_i, ALU_OPCODE_i_0_port, 
      ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_4_port, ALUA_SEL_i, MEM_EN_i, MEM_DATA_SEL_i, 
      LD_SEL_i_2_port, LD_SEL_i_1_port, LD_SEL_i_0_port, ALR2_SEL_i, 
      CWB_SEL_i_1_port, CWB_SEL_i_0_port, WB_SEL_i, RF_WR_i, 
      RF_MUX_SEL_i_1_port, RF_MUX_SEL_i_0_port, n1, n_1819, n_1820, n_1821, 
      n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828 : std_logic;
   
   signal ALU_OPCODE_pin : std_logic_vector (0 to 4);

begin
   
   ( ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port ) <= ALU_OPCODE_pin;
   CU_I : CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26
      port map( Clk => Clk, Rst => Rst, STALL(1) => STALL_CODE_1_port, STALL(0)
      => STALL_CODE_0_port, IR_IN(31) => IRAM_OUT(31), IR_IN(30) => 
      IRAM_OUT(30), IR_IN(29) => IRAM_OUT(29), IR_IN(28) => IRAM_OUT(28), 
      IR_IN(27) => IRAM_OUT(27), IR_IN(26) => IRAM_OUT(26), IR_IN(25) => 
      IRAM_OUT(25), IR_IN(24) => IRAM_OUT(24), IR_IN(23) => IRAM_OUT(23), 
      IR_IN(22) => IRAM_OUT(22), IR_IN(21) => IRAM_OUT(21), IR_IN(20) => 
      IRAM_OUT(20), IR_IN(19) => IRAM_OUT(19), IR_IN(18) => IRAM_OUT(18), 
      IR_IN(17) => IRAM_OUT(17), IR_IN(16) => IRAM_OUT(16), IR_IN(15) => 
      IRAM_OUT(15), IR_IN(14) => IRAM_OUT(14), IR_IN(13) => IRAM_OUT(13), 
      IR_IN(12) => IRAM_OUT(12), IR_IN(11) => IRAM_OUT(11), IR_IN(10) => 
      IRAM_OUT(10), IR_IN(9) => IRAM_OUT(9), IR_IN(8) => IRAM_OUT(8), IR_IN(7) 
      => IRAM_OUT(7), IR_IN(6) => IRAM_OUT(6), IR_IN(5) => IRAM_OUT(5), 
      IR_IN(4) => IRAM_OUT(4), IR_IN(3) => IRAM_OUT(3), IR_IN(2) => IRAM_OUT(2)
      , IR_IN(1) => IRAM_OUT(1), IR_IN(0) => IRAM_OUT(0), BMP => BMP_i, ID_EN 
      => n_1819, RF_RD => n_1820, SIGND => n_1821, IMM_SEL => n_1822, BPR_EN =>
      n_1823, UCB_EN => n_1824, ALU_OPCODE => ALU_OPCODE_pin, EX_EN => n_1825, 
      ALUA_SEL => n_1826, ALUB_SEL => n_1827, MEM_EN => MEM_EN_i, MEM_DATA_SEL 
      => MEM_DATA_SEL_i, MEM_RD => MEM_RD, MEM_WR => MEM_WR, CS => n_1828, 
      MEM_BLC0 => BLC(0), MEM_BLC1 => BLC(1), LD_SEL0 => LD_SEL_i_0_port, 
      LD_SEL1 => LD_SEL_i_1_port, LD_SEL2 => LD_SEL_i_2_port, ALR2_SEL => 
      ALR2_SEL_i, CWB_SEL0 => CWB_SEL_i_0_port, CWB_SEL1 => CWB_SEL_i_1_port, 
      WB_SEL => WB_SEL_i, RF_WR => RF_WR_i, RF_MUX_SEL0 => RF_MUX_SEL_i_0_port,
      RF_MUX_SEL1 => RF_MUX_SEL_i_1_port);
   DATAP : Datapath port map( CLK => Clk, RST => Rst, DATA_IN(31) => 
                           DATA_IN(31), DATA_IN(30) => DATA_IN(30), DATA_IN(29)
                           => DATA_IN(29), DATA_IN(28) => DATA_IN(28), 
                           DATA_IN(27) => DATA_IN(27), DATA_IN(26) => 
                           DATA_IN(26), DATA_IN(25) => DATA_IN(25), DATA_IN(24)
                           => DATA_IN(24), DATA_IN(23) => DATA_IN(23), 
                           DATA_IN(22) => DATA_IN(22), DATA_IN(21) => 
                           DATA_IN(21), DATA_IN(20) => DATA_IN(20), DATA_IN(19)
                           => DATA_IN(19), DATA_IN(18) => DATA_IN(18), 
                           DATA_IN(17) => DATA_IN(17), DATA_IN(16) => 
                           DATA_IN(16), DATA_IN(15) => DATA_IN(15), DATA_IN(14)
                           => DATA_IN(14), DATA_IN(13) => DATA_IN(13), 
                           DATA_IN(12) => DATA_IN(12), DATA_IN(11) => 
                           DATA_IN(11), DATA_IN(10) => DATA_IN(10), DATA_IN(9) 
                           => DATA_IN(9), DATA_IN(8) => DATA_IN(8), DATA_IN(7) 
                           => DATA_IN(7), DATA_IN(6) => DATA_IN(6), DATA_IN(5) 
                           => DATA_IN(5), DATA_IN(4) => DATA_IN(4), DATA_IN(3) 
                           => DATA_IN(3), DATA_IN(2) => DATA_IN(2), DATA_IN(1) 
                           => DATA_IN(1), DATA_IN(0) => DATA_IN(0), 
                           IRAM_OUT(31) => IRAM_OUT(31), IRAM_OUT(30) => 
                           IRAM_OUT(30), IRAM_OUT(29) => IRAM_OUT(29), 
                           IRAM_OUT(28) => IRAM_OUT(28), IRAM_OUT(27) => 
                           IRAM_OUT(27), IRAM_OUT(26) => IRAM_OUT(26), 
                           IRAM_OUT(25) => IRAM_OUT(25), IRAM_OUT(24) => 
                           IRAM_OUT(24), IRAM_OUT(23) => IRAM_OUT(23), 
                           IRAM_OUT(22) => IRAM_OUT(22), IRAM_OUT(21) => 
                           IRAM_OUT(21), IRAM_OUT(20) => IRAM_OUT(20), 
                           IRAM_OUT(19) => IRAM_OUT(19), IRAM_OUT(18) => 
                           IRAM_OUT(18), IRAM_OUT(17) => IRAM_OUT(17), 
                           IRAM_OUT(16) => IRAM_OUT(16), IRAM_OUT(15) => 
                           IRAM_OUT(15), IRAM_OUT(14) => IRAM_OUT(14), 
                           IRAM_OUT(13) => IRAM_OUT(13), IRAM_OUT(12) => 
                           IRAM_OUT(12), IRAM_OUT(11) => IRAM_OUT(11), 
                           IRAM_OUT(10) => IRAM_OUT(10), IRAM_OUT(9) => 
                           IRAM_OUT(9), IRAM_OUT(8) => IRAM_OUT(8), IRAM_OUT(7)
                           => IRAM_OUT(7), IRAM_OUT(6) => IRAM_OUT(6), 
                           IRAM_OUT(5) => IRAM_OUT(5), IRAM_OUT(4) => 
                           IRAM_OUT(4), IRAM_OUT(3) => IRAM_OUT(3), IRAM_OUT(2)
                           => IRAM_OUT(2), IRAM_OUT(1) => IRAM_OUT(1), 
                           IRAM_OUT(0) => IRAM_OUT(0), IRAM_ADDR(31) => 
                           IRAM_ADDR(31), IRAM_ADDR(30) => IRAM_ADDR(30), 
                           IRAM_ADDR(29) => IRAM_ADDR(29), IRAM_ADDR(28) => 
                           IRAM_ADDR(28), IRAM_ADDR(27) => IRAM_ADDR(27), 
                           IRAM_ADDR(26) => IRAM_ADDR(26), IRAM_ADDR(25) => 
                           IRAM_ADDR(25), IRAM_ADDR(24) => IRAM_ADDR(24), 
                           IRAM_ADDR(23) => IRAM_ADDR(23), IRAM_ADDR(22) => 
                           IRAM_ADDR(22), IRAM_ADDR(21) => IRAM_ADDR(21), 
                           IRAM_ADDR(20) => IRAM_ADDR(20), IRAM_ADDR(19) => 
                           IRAM_ADDR(19), IRAM_ADDR(18) => IRAM_ADDR(18), 
                           IRAM_ADDR(17) => IRAM_ADDR(17), IRAM_ADDR(16) => 
                           IRAM_ADDR(16), IRAM_ADDR(15) => IRAM_ADDR(15), 
                           IRAM_ADDR(14) => IRAM_ADDR(14), IRAM_ADDR(13) => 
                           IRAM_ADDR(13), IRAM_ADDR(12) => IRAM_ADDR(12), 
                           IRAM_ADDR(11) => IRAM_ADDR(11), IRAM_ADDR(10) => 
                           IRAM_ADDR(10), IRAM_ADDR(9) => IRAM_ADDR(9), 
                           IRAM_ADDR(8) => IRAM_ADDR(8), IRAM_ADDR(7) => 
                           IRAM_ADDR(7), IRAM_ADDR(6) => IRAM_ADDR(6), 
                           IRAM_ADDR(5) => IRAM_ADDR(5), IRAM_ADDR(4) => 
                           IRAM_ADDR(4), IRAM_ADDR(3) => IRAM_ADDR(3), 
                           IRAM_ADDR(2) => IRAM_ADDR(2), IRAM_ADDR(1) => 
                           IRAM_ADDR(1), IRAM_ADDR(0) => IRAM_ADDR(0), 
                           DATA_OUT(31) => DATA_OUT(31), DATA_OUT(30) => 
                           DATA_OUT(30), DATA_OUT(29) => DATA_OUT(29), 
                           DATA_OUT(28) => DATA_OUT(28), DATA_OUT(27) => 
                           DATA_OUT(27), DATA_OUT(26) => DATA_OUT(26), 
                           DATA_OUT(25) => DATA_OUT(25), DATA_OUT(24) => 
                           DATA_OUT(24), DATA_OUT(23) => DATA_OUT(23), 
                           DATA_OUT(22) => DATA_OUT(22), DATA_OUT(21) => 
                           DATA_OUT(21), DATA_OUT(20) => DATA_OUT(20), 
                           DATA_OUT(19) => DATA_OUT(19), DATA_OUT(18) => 
                           DATA_OUT(18), DATA_OUT(17) => DATA_OUT(17), 
                           DATA_OUT(16) => DATA_OUT(16), DATA_OUT(15) => 
                           DATA_OUT(15), DATA_OUT(14) => DATA_OUT(14), 
                           DATA_OUT(13) => DATA_OUT(13), DATA_OUT(12) => 
                           DATA_OUT(12), DATA_OUT(11) => DATA_OUT(11), 
                           DATA_OUT(10) => DATA_OUT(10), DATA_OUT(9) => 
                           DATA_OUT(9), DATA_OUT(8) => DATA_OUT(8), DATA_OUT(7)
                           => DATA_OUT(7), DATA_OUT(6) => DATA_OUT(6), 
                           DATA_OUT(5) => DATA_OUT(5), DATA_OUT(4) => 
                           DATA_OUT(4), DATA_OUT(3) => DATA_OUT(3), DATA_OUT(2)
                           => DATA_OUT(2), DATA_OUT(1) => DATA_OUT(1), 
                           DATA_OUT(0) => DATA_OUT(0), DATA_ADDR(31) => 
                           DATA_ADDR(31), DATA_ADDR(30) => DATA_ADDR(30), 
                           DATA_ADDR(29) => DATA_ADDR(29), DATA_ADDR(28) => 
                           DATA_ADDR(28), DATA_ADDR(27) => DATA_ADDR(27), 
                           DATA_ADDR(26) => DATA_ADDR(26), DATA_ADDR(25) => 
                           DATA_ADDR(25), DATA_ADDR(24) => DATA_ADDR(24), 
                           DATA_ADDR(23) => DATA_ADDR(23), DATA_ADDR(22) => 
                           DATA_ADDR(22), DATA_ADDR(21) => DATA_ADDR(21), 
                           DATA_ADDR(20) => DATA_ADDR(20), DATA_ADDR(19) => 
                           DATA_ADDR(19), DATA_ADDR(18) => DATA_ADDR(18), 
                           DATA_ADDR(17) => DATA_ADDR(17), DATA_ADDR(16) => 
                           DATA_ADDR(16), DATA_ADDR(15) => DATA_ADDR(15), 
                           DATA_ADDR(14) => DATA_ADDR(14), DATA_ADDR(13) => 
                           DATA_ADDR(13), DATA_ADDR(12) => DATA_ADDR(12), 
                           DATA_ADDR(11) => DATA_ADDR(11), DATA_ADDR(10) => 
                           DATA_ADDR(10), DATA_ADDR(9) => DATA_ADDR(9), 
                           DATA_ADDR(8) => DATA_ADDR(8), DATA_ADDR(7) => 
                           DATA_ADDR(7), DATA_ADDR(6) => DATA_ADDR(6), 
                           DATA_ADDR(5) => DATA_ADDR(5), DATA_ADDR(4) => 
                           DATA_ADDR(4), DATA_ADDR(3) => DATA_ADDR(3), 
                           DATA_ADDR(2) => DATA_ADDR(2), DATA_ADDR(1) => 
                           DATA_ADDR(1), DATA_ADDR(0) => DATA_ADDR(0), BMP => 
                           BMP_i, STALL(1) => STALL_CODE_1_port, STALL(0) => 
                           STALL_CODE_0_port, ID_EN => ID_EN_i, RF_RD => 
                           RF_RD_i, SIGND => SIGND_i, IMM_SEL => IMM_SEL_i, 
                           BPR_EN => BPR_EN_i, ALU_OPCODE(0) => 
                           ALU_OPCODE_i_0_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, EX_EN => n1, ALUA_SEL => 
                           ALUA_SEL_i, ALUB_SEL => n1, UCB_EN => UCB_EN_i, 
                           MEM_EN => MEM_EN_i, MEM_DATA_SEL => MEM_DATA_SEL_i, 
                           LD_SEL(2) => LD_SEL_i_2_port, LD_SEL(1) => 
                           LD_SEL_i_1_port, LD_SEL(0) => LD_SEL_i_0_port, 
                           ALR2_SEL => ALR2_SEL_i, CWB_SEL(1) => 
                           CWB_SEL_i_1_port, CWB_SEL(0) => CWB_SEL_i_0_port, 
                           WB_SEL => WB_SEL_i, RF_WR => RF_WR_i, RF_MUX_SEL(1) 
                           => RF_MUX_SEL_i_1_port, RF_MUX_SEL(0) => 
                           RF_MUX_SEL_i_0_port);
   n1 <= '0';
   ALUA_SEL_i <= '0';
   UCB_EN_i <= '0';
   BPR_EN_i <= '0';
   IMM_SEL_i <= '0';
   SIGND_i <= '0';
   RF_RD_i <= '0';
   ID_EN_i <= '0';

end SYN_dlx_rtl;
