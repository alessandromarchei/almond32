
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_NOP, OP_ADD, OP_ADC, OP_AND, OP_SRA, OP_OR, OP_SEQ, OP_SNE, 
   OP_SLT, OP_SGT, OP_SLE, OP_SGE, OP_SLL, OP_SRL, OP_SUB, OP_XOR, OP_NOR, 
   OP_XNOR, OP_NAND, OP_MUL);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011";

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_0_DW01_add_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_adder_0_DW01_add_2;

architecture SYN_cla of PC_adder_0_DW01_add_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n123, B2 => n124, A => n125, ZN => n120);
   U3 : NAND2_X1 port map( A1 => n61, A2 => n59, ZN => n1);
   U4 : INV_X1 port map( A => n11, ZN => n66);
   U5 : AND2_X1 port map( A1 => n70, A2 => n4, ZN => n2);
   U6 : OR2_X1 port map( A1 => n2, A2 => n3, ZN => n7);
   U7 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => n3);
   U8 : AND2_X1 port map( A1 => n71, A2 => n1, ZN => n4);
   U9 : CLKBUF_X1 port map( A => n140, Z => n5);
   U10 : INV_X1 port map( A => n61, ZN => n6);
   U11 : OR2_X1 port map( A1 => n9, A2 => n6, ZN => n8);
   U12 : INV_X1 port map( A => n69, ZN => n9);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n60);
   U14 : AND2_X1 port map( A1 => n70, A2 => n71, ZN => n10);
   U15 : NOR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n11);
   U16 : XOR2_X1 port map( A => n12, B => n60, Z => SUM(29));
   U17 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => n12);
   U18 : AND2_X1 port map( A1 => n5, A2 => n214, ZN => SUM(0));
   U19 : AOI21_X1 port map( B1 => n156, B2 => n157, A => n158, ZN => n154);
   U20 : OAI21_X1 port map( B1 => n212, B2 => n176, A => n156, ZN => n23);
   U21 : NAND2_X1 port map( A1 => n189, A2 => n190, ZN => n187);
   U22 : NAND2_X1 port map( A1 => n173, A2 => n23, ZN => n190);
   U23 : INV_X1 port map( A => n212, ZN => n45);
   U24 : NOR2_X1 port map( A1 => n17, A2 => n76, ZN => n75);
   U25 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n76);
   U26 : NOR2_X1 port map( A1 => n16, A2 => n101, ZN => n100);
   U27 : AOI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n101);
   U28 : NOR2_X1 port map( A1 => n126, A2 => n127, ZN => n125);
   U29 : NAND4_X1 port map( A1 => n191, A2 => n192, A3 => n20, A4 => n25, ZN =>
                           n158);
   U30 : INV_X1 port map( A => n161, ZN => n152);
   U31 : OAI21_X1 port map( B1 => n162, B2 => n163, A => n164, ZN => n161);
   U32 : XNOR2_X1 port map( A => n7, B => n58, ZN => SUM(30));
   U33 : NAND2_X1 port map( A1 => n57, A2 => n55, ZN => n58);
   U34 : AND4_X1 port map( A1 => n174, A2 => n175, A3 => n166, A4 => n165, ZN 
                           => n14);
   U35 : XNOR2_X1 port map( A => n87, B => n88, ZN => SUM(27));
   U36 : NOR2_X1 port map( A1 => n79, A2 => n17, ZN => n88);
   U37 : AOI21_X1 port map( B1 => n80, B2 => n89, A => n90, ZN => n87);
   U38 : NAND2_X1 port map( A1 => n92, A2 => n84, ZN => n89);
   U39 : NAND2_X1 port map( A1 => n85, A2 => n93, ZN => n92);
   U40 : OAI21_X1 port map( B1 => n215, B2 => n213, A => n53, ZN => n160);
   U41 : AOI21_X1 port map( B1 => n68, B2 => n216, A => n217, ZN => n215);
   U42 : OAI21_X1 port map( B1 => n11, B2 => n140, A => n65, ZN => n216);
   U43 : OAI21_X1 port map( B1 => n182, B2 => n170, A => n172, ZN => n180);
   U44 : XNOR2_X1 port map( A => n177, B => n178, ZN => SUM(15));
   U45 : NAND2_X1 port map( A1 => n164, A2 => n165, ZN => n177);
   U46 : NAND2_X1 port map( A1 => n179, A2 => n169, ZN => n178);
   U47 : NAND2_X1 port map( A1 => n166, A2 => n180, ZN => n179);
   U48 : OAI21_X1 port map( B1 => n185, B2 => n186, A => n171, ZN => n183);
   U49 : XNOR2_X1 port map( A => n89, B => n91, ZN => SUM(26));
   U50 : NAND2_X1 port map( A1 => n78, A2 => n80, ZN => n91);
   U51 : NAND4_X1 port map( A1 => n42, A2 => n43, A3 => n30, A4 => n32, ZN => 
                           n176);
   U52 : XNOR2_X1 port map( A => n112, B => n113, ZN => SUM(23));
   U53 : NOR2_X1 port map( A1 => n104, A2 => n16, ZN => n113);
   U54 : AOI21_X1 port map( B1 => n105, B2 => n114, A => n115, ZN => n112);
   U55 : NAND2_X1 port map( A1 => n117, A2 => n109, ZN => n114);
   U56 : NAND2_X1 port map( A1 => n110, A2 => n118, ZN => n117);
   U57 : XNOR2_X1 port map( A => n70, B => n72, ZN => SUM(28));
   U58 : NAND2_X1 port map( A1 => n69, A2 => n71, ZN => n72);
   U59 : XNOR2_X1 port map( A => n181, B => n180, ZN => SUM(14));
   U60 : NAND2_X1 port map( A1 => n169, A2 => n166, ZN => n181);
   U61 : OAI21_X1 port map( B1 => n199, B2 => n205, A => n21, ZN => n203);
   U62 : XNOR2_X1 port map( A => n200, B => n201, ZN => SUM(11));
   U63 : NAND2_X1 port map( A1 => n195, A2 => n191, ZN => n201);
   U64 : NAND2_X1 port map( A1 => n198, A2 => n202, ZN => n200);
   U65 : NAND2_X1 port map( A1 => n203, A2 => n192, ZN => n202);
   U66 : NAND2_X1 port map( A1 => n206, A2 => n24, ZN => n19);
   U67 : NAND2_X1 port map( A1 => n23, A2 => n25, ZN => n206);
   U68 : XNOR2_X1 port map( A => n94, B => n93, ZN => SUM(25));
   U69 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => n94);
   U70 : XNOR2_X1 port map( A => n141, B => n142, ZN => SUM(19));
   U71 : NAND2_X1 port map( A1 => n138, A2 => n131, ZN => n142);
   U72 : NAND2_X1 port map( A1 => n129, A2 => n143, ZN => n141);
   U73 : NAND2_X1 port map( A1 => n144, A2 => n132, ZN => n143);
   U74 : NAND2_X1 port map( A1 => n123, A2 => n135, ZN => n147);
   U75 : NAND2_X1 port map( A1 => n146, A2 => n136, ZN => n144);
   U76 : NAND2_X1 port map( A1 => n137, A2 => n147, ZN => n146);
   U77 : XNOR2_X1 port map( A => n114, B => n116, ZN => SUM(22));
   U78 : NAND2_X1 port map( A1 => n103, A2 => n105, ZN => n116);
   U79 : XNOR2_X1 port map( A => n95, B => n97, ZN => SUM(24));
   U80 : NAND2_X1 port map( A1 => n83, A2 => n96, ZN => n97);
   U81 : XNOR2_X1 port map( A => n184, B => n183, ZN => SUM(13));
   U82 : NAND2_X1 port map( A1 => n172, A2 => n175, ZN => n184);
   U83 : XNOR2_X1 port map( A => n204, B => n203, ZN => SUM(10));
   U84 : NAND2_X1 port map( A1 => n198, A2 => n192, ZN => n204);
   U85 : XNOR2_X1 port map( A => n145, B => n144, ZN => SUM(18));
   U86 : NAND2_X1 port map( A1 => n129, A2 => n132, ZN => n145);
   U87 : OAI21_X1 port map( B1 => n35, B2 => n36, A => n37, ZN => n31);
   U88 : OAI21_X1 port map( B1 => n40, B2 => n212, A => n41, ZN => n38);
   U89 : XNOR2_X1 port map( A => n26, B => n27, ZN => SUM(7));
   U90 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => n26);
   U91 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n27);
   U92 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => n28);
   U93 : XNOR2_X1 port map( A => n119, B => n118, ZN => SUM(21));
   U94 : NAND2_X1 port map( A1 => n109, A2 => n110, ZN => n119);
   U95 : XNOR2_X1 port map( A => n188, B => n187, ZN => SUM(12));
   U96 : NAND2_X1 port map( A1 => n171, A2 => n174, ZN => n188);
   U97 : XNOR2_X1 port map( A => n18, B => n19, ZN => SUM(9));
   U98 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n18);
   U99 : XNOR2_X1 port map( A => n34, B => n31, ZN => SUM(6));
   U100 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => n34);
   U101 : XNOR2_X1 port map( A => n148, B => n147, ZN => SUM(17));
   U102 : NAND2_X1 port map( A1 => n136, A2 => n137, ZN => n148);
   U103 : NAND2_X1 port map( A1 => n108, A2 => n121, ZN => n122);
   U104 : XNOR2_X1 port map( A => n22, B => n23, ZN => SUM(8));
   U105 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => n22);
   U106 : XNOR2_X1 port map( A => n39, B => n38, ZN => SUM(5));
   U107 : NAND2_X1 port map( A1 => n43, A2 => n37, ZN => n39);
   U108 : NAND2_X1 port map( A1 => n135, A2 => n150, ZN => n151);
   U109 : XNOR2_X1 port map( A => n44, B => n45, ZN => SUM(4));
   U110 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => n44);
   U111 : XNOR2_X1 port map( A => n46, B => n47, ZN => SUM(3));
   U112 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n46);
   U113 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n50, ZN => n47);
   U114 : INV_X1 port map( A => n5, ZN => n67);
   U115 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n51);
   U116 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => n64);
   U117 : XNOR2_X1 port map( A => n63, B => n51, ZN => SUM(2));
   U118 : NAND2_X1 port map( A1 => n68, A2 => n50, ZN => n63);
   U119 : XNOR2_X1 port map( A => n139, B => n67, ZN => SUM(1));
   U120 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => n139);
   U121 : AOI21_X1 port map( B1 => n128, B2 => n129, A => n130, ZN => n127);
   U122 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => n128);
   U123 : OAI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n133);
   U124 : AOI21_X1 port map( B1 => n166, B2 => n167, A => n168, ZN => n162);
   U125 : OAI21_X1 port map( B1 => n170, B2 => n171, A => n172, ZN => n167);
   U126 : OAI21_X1 port map( B1 => n193, B2 => n194, A => n195, ZN => n155);
   U127 : AOI21_X1 port map( B1 => n192, B2 => n196, A => n197, ZN => n193);
   U128 : OAI21_X1 port map( B1 => n36, B2 => n41, A => n37, ZN => n210);
   U129 : OAI21_X1 port map( B1 => n199, B2 => n24, A => n21, ZN => n196);
   U130 : OAI21_X1 port map( B1 => n208, B2 => n209, A => n33, ZN => n207);
   U131 : AOI21_X1 port map( B1 => n30, B2 => n210, A => n211, ZN => n208);
   U132 : NAND2_X1 port map( A1 => n105, A2 => n106, ZN => n102);
   U133 : OAI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n106);
   U134 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n77);
   U135 : OAI21_X1 port map( B1 => n82, B2 => n83, A => n84, ZN => n81);
   U136 : INV_X1 port map( A => A(0), ZN => n219);
   U137 : XOR2_X1 port map( A => B(31), B => A(31), Z => n15);
   U138 : OR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n191);
   U139 : OR2_X1 port map( A1 => B(14), A2 => A(14), ZN => n166);
   U140 : OR2_X1 port map( A1 => B(15), A2 => A(15), ZN => n165);
   U141 : OR2_X1 port map( A1 => B(13), A2 => A(13), ZN => n175);
   U142 : OR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n174);
   U143 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n140);
   U144 : OR2_X1 port map( A1 => B(6), A2 => A(6), ZN => n30);
   U145 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n32);
   U146 : OR2_X1 port map( A1 => B(2), A2 => A(2), ZN => n68);
   U147 : OR2_X1 port map( A1 => B(5), A2 => A(5), ZN => n43);
   U148 : OR2_X1 port map( A1 => B(4), A2 => A(4), ZN => n42);
   U149 : OR2_X1 port map( A1 => B(3), A2 => A(3), ZN => n52);
   U150 : OR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n192);
   U151 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n25);
   U152 : OR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n20);
   U153 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n132);
   U154 : OR2_X1 port map( A1 => B(17), A2 => A(17), ZN => n137);
   U155 : OR2_X1 port map( A1 => B(19), A2 => A(19), ZN => n131);
   U156 : OR2_X1 port map( A1 => B(16), A2 => A(16), ZN => n150);
   U157 : OR2_X1 port map( A1 => B(21), A2 => A(21), ZN => n110);
   U158 : OR2_X1 port map( A1 => B(22), A2 => A(22), ZN => n105);
   U159 : OR2_X1 port map( A1 => B(23), A2 => A(23), ZN => n111);
   U160 : OR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n121);
   U161 : OR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n85);
   U162 : OR2_X1 port map( A1 => B(26), A2 => A(26), ZN => n80);
   U163 : OR2_X1 port map( A1 => B(27), A2 => A(27), ZN => n86);
   U164 : OR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n96);
   U165 : OR2_X1 port map( A1 => B(28), A2 => A(28), ZN => n71);
   U166 : OR2_X1 port map( A1 => B(29), A2 => A(29), ZN => n62);
   U167 : OR2_X1 port map( A1 => B(30), A2 => A(30), ZN => n55);
   U168 : NAND2_X1 port map( A1 => n218, A2 => n219, ZN => n214);
   U169 : INV_X1 port map( A => B(0), ZN => n218);
   U170 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n16);
   U171 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => n17);
   U172 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n65);
   U173 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n24);
   U174 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n135);
   U175 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n37);
   U176 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n21);
   U177 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n136);
   U178 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n109);
   U179 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n84);
   U180 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n129);
   U181 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n41);
   U182 : NAND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n171);
   U183 : NAND2_X1 port map( A1 => B(13), A2 => A(13), ZN => n172);
   U184 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n29);
   U185 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n50);
   U186 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n103);
   U187 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => n78);
   U188 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n169);
   U189 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n108);
   U190 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n83);
   U191 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n198);
   U192 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n53);
   U193 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n33);
   U194 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n195);
   U195 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n164);
   U196 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n61);
   U197 : NAND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n69);
   U198 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n138);
   U199 : NAND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n57);
   U200 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U201 : NAND2_X1 port map( A1 => n98, A2 => n108, ZN => n118);
   U202 : XNOR2_X1 port map( A => n149, B => n151, ZN => SUM(16));
   U203 : NAND2_X1 port map( A1 => n73, A2 => n83, ZN => n93);
   U204 : OAI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n70);
   U205 : NAND2_X1 port map( A1 => n149, A2 => n150, ZN => n123);
   U206 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => n149);
   U207 : OAI21_X1 port map( B1 => n154, B2 => n155, A => n14, ZN => n153);
   U208 : NAND2_X1 port map( A1 => n159, A2 => n160, ZN => n157);
   U209 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => n73);
   U210 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => n98);
   U211 : XNOR2_X1 port map( A => n54, B => n15, ZN => SUM(31));
   U212 : INV_X1 port map( A => n38, ZN => n35);
   U213 : INV_X1 port map( A => n42, ZN => n40);
   U214 : INV_X1 port map( A => n51, ZN => n48);
   U215 : AOI21_X1 port map( B1 => n7, B2 => n55, A => n56, ZN => n54);
   U216 : INV_X1 port map( A => n57, ZN => n56);
   U217 : INV_X1 port map( A => n62, ZN => n59);
   U218 : INV_X1 port map( A => n85, ZN => n82);
   U219 : NAND3_X1 port map( A1 => n80, A2 => n86, A3 => n85, ZN => n74);
   U220 : INV_X1 port map( A => n86, ZN => n79);
   U221 : INV_X1 port map( A => n78, ZN => n90);
   U222 : INV_X1 port map( A => n110, ZN => n107);
   U223 : NAND3_X1 port map( A1 => n105, A2 => n111, A3 => n110, ZN => n99);
   U224 : INV_X1 port map( A => n111, ZN => n104);
   U225 : INV_X1 port map( A => n103, ZN => n115);
   U226 : XNOR2_X1 port map( A => n122, B => n120, ZN => SUM(20));
   U227 : INV_X1 port map( A => n131, ZN => n130);
   U228 : INV_X1 port map( A => n137, ZN => n134);
   U229 : INV_X1 port map( A => n138, ZN => n126);
   U230 : NAND3_X1 port map( A1 => n132, A2 => n131, A3 => n137, ZN => n124);
   U231 : INV_X1 port map( A => n165, ZN => n163);
   U232 : INV_X1 port map( A => n169, ZN => n168);
   U233 : INV_X1 port map( A => n176, ZN => n159);
   U234 : INV_X1 port map( A => n175, ZN => n170);
   U235 : INV_X1 port map( A => n183, ZN => n182);
   U236 : INV_X1 port map( A => n187, ZN => n186);
   U237 : INV_X1 port map( A => n174, ZN => n185);
   U238 : INV_X1 port map( A => n158, ZN => n173);
   U239 : INV_X1 port map( A => n155, ZN => n189);
   U240 : INV_X1 port map( A => n191, ZN => n194);
   U241 : INV_X1 port map( A => n198, ZN => n197);
   U242 : INV_X1 port map( A => n19, ZN => n205);
   U243 : INV_X1 port map( A => n207, ZN => n156);
   U244 : INV_X1 port map( A => n32, ZN => n209);
   U245 : INV_X1 port map( A => n29, ZN => n211);
   U246 : INV_X1 port map( A => n43, ZN => n36);
   U247 : INV_X1 port map( A => n68, ZN => n49);
   U248 : INV_X1 port map( A => n160, ZN => n212);
   U249 : INV_X1 port map( A => n52, ZN => n213);
   U250 : INV_X1 port map( A => n50, ZN => n217);
   U251 : INV_X1 port map( A => n20, ZN => n199);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_1_DW01_add_0_DW01_add_128 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_adder_1_DW01_add_0_DW01_add_128;

architecture SYN_rpl of PC_adder_1_DW01_add_0_DW01_add_128 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1004 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1004, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1;

architecture SYN_rpl of HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n46, n47, n48
      , n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
      n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n53, A2 => A(18), ZN => n103);
   U2 : INV_X1 port map( A => n11, ZN => n102);
   U3 : NOR2_X1 port map( A1 => n11, A2 => A(20), ZN => n101);
   U4 : INV_X1 port map( A => n1, ZN => n100);
   U5 : NOR2_X1 port map( A1 => n1, A2 => A(22), ZN => n99);
   U6 : INV_X1 port map( A => n8, ZN => n96);
   U7 : INV_X1 port map( A => A(31), ZN => n5);
   U8 : INV_X1 port map( A => A(19), ZN => n12);
   U9 : INV_X1 port map( A => A(25), ZN => n9);
   U10 : INV_X1 port map( A => A(21), ZN => n2);
   U11 : INV_X1 port map( A => A(23), ZN => n7);
   U12 : INV_X1 port map( A => A(27), ZN => n10);
   U13 : NAND2_X1 port map( A1 => n101, A2 => n2, ZN => n1);
   U14 : AND2_X2 port map( A1 => n99, A2 => n7, ZN => n98);
   U15 : NAND2_X1 port map( A1 => n98, A2 => n3, ZN => n8);
   U16 : NOR2_X1 port map( A1 => A(24), A2 => A(25), ZN => n3);
   U17 : INV_X1 port map( A => n4, ZN => n107);
   U18 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => n4);
   U19 : XNOR2_X1 port map( A => n5, B => n6, ZN => SUM(31));
   U20 : NOR2_X1 port map( A1 => A(30), A2 => n90, ZN => n6);
   U21 : AND2_X2 port map( A1 => n95, A2 => n42, ZN => n92);
   U22 : AND2_X1 port map( A1 => n94, A2 => n10, ZN => n95);
   U23 : NAND2_X1 port map( A1 => n103, A2 => n12, ZN => n11);
   U24 : INV_X1 port map( A => A(17), ZN => n15);
   U25 : OR2_X1 port map( A1 => n4, A2 => A(15), ZN => n13);
   U26 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => n104);
   U27 : OR2_X1 port map( A1 => A(17), A2 => A(16), ZN => n14);
   U28 : OR2_X1 port map( A1 => n4, A2 => A(15), ZN => n16);
   U29 : AND2_X1 port map( A1 => n114, A2 => n41, ZN => n84);
   U30 : INV_X1 port map( A => A(28), ZN => n42);
   U31 : INV_X1 port map( A => n93, ZN => SUM(28));
   U32 : INV_X1 port map( A => n112, ZN => SUM(11));
   U33 : INV_X1 port map( A => n109, ZN => SUM(13));
   U34 : INV_X1 port map( A => A(26), ZN => n66);
   U35 : INV_X1 port map( A => n81, ZN => SUM(9));
   U36 : INV_X1 port map( A => A(15), ZN => n72);
   U37 : INV_X1 port map( A => A(16), ZN => n71);
   U38 : INV_X1 port map( A => A(18), ZN => n70);
   U39 : INV_X1 port map( A => A(20), ZN => n69);
   U40 : INV_X1 port map( A => A(22), ZN => n68);
   U41 : INV_X1 port map( A => A(24), ZN => n67);
   U42 : INV_X1 port map( A => n85, ZN => SUM(7));
   U43 : INV_X1 port map( A => A(2), ZN => n80);
   U44 : INV_X1 port map( A => A(3), ZN => n79);
   U45 : INV_X1 port map( A => A(4), ZN => n78);
   U46 : INV_X1 port map( A => A(6), ZN => n76);
   U47 : INV_X1 port map( A => A(10), ZN => n74);
   U48 : INV_X1 port map( A => A(12), ZN => n73);
   U49 : INV_X1 port map( A => A(29), ZN => n65);
   U50 : INV_X1 port map( A => n94, ZN => n47);
   U51 : NOR2_X1 port map( A1 => n60, A2 => A(4), ZN => n17);
   U52 : AND2_X1 port map( A1 => n17, A2 => n18, ZN => n20);
   U53 : AND2_X1 port map( A1 => n21, A2 => n77, ZN => n18);
   U54 : NOR2_X1 port map( A1 => n22, A2 => A(6), ZN => n19);
   U55 : INV_X1 port map( A => A(14), ZN => n21);
   U56 : AND2_X1 port map( A1 => n87, A2 => n77, ZN => n86);
   U57 : INV_X1 port map( A => A(5), ZN => n77);
   U58 : INV_X1 port map( A => A(8), ZN => n75);
   U59 : INV_X1 port map( A => n24, ZN => n22);
   U60 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n23);
   U61 : AND2_X1 port map( A1 => n23, A2 => n24, ZN => n108);
   U62 : AND2_X1 port map( A1 => n25, A2 => n27, ZN => n24);
   U63 : INV_X1 port map( A => A(13), ZN => n25);
   U64 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n26);
   U65 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n110);
   U66 : AND2_X1 port map( A1 => n73, A2 => n29, ZN => n27);
   U67 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n28);
   U68 : AND2_X1 port map( A1 => n28, A2 => n29, ZN => n111);
   U69 : AND2_X1 port map( A1 => n30, A2 => n32, ZN => n29);
   U70 : INV_X1 port map( A => A(11), ZN => n30);
   U71 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n31);
   U72 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => n113);
   U73 : AND2_X1 port map( A1 => n74, A2 => n34, ZN => n32);
   U74 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n33);
   U75 : AND2_X1 port map( A1 => n33, A2 => n34, ZN => n83);
   U76 : AND2_X1 port map( A1 => n35, A2 => n37, ZN => n34);
   U77 : INV_X1 port map( A => A(9), ZN => n35);
   U78 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n36);
   U79 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n82);
   U80 : AND2_X1 port map( A1 => n75, A2 => n41, ZN => n37);
   U81 : INV_X1 port map( A => A(7), ZN => n41);
   U82 : CLKBUF_X1 port map( A => n53, Z => n38);
   U83 : CLKBUF_X1 port map( A => n4, Z => n39);
   U84 : INV_X1 port map( A => A(1), ZN => n64);
   U85 : CLKBUF_X1 port map( A => n1, Z => n40);
   U86 : INV_X1 port map( A => n86, ZN => n58);
   U87 : INV_X1 port map( A => A(0), ZN => n63);
   U88 : INV_X1 port map( A => n91, ZN => n62);
   U89 : INV_X1 port map( A => n98, ZN => n49);
   U90 : INV_X1 port map( A => n101, ZN => n51);
   U91 : INV_X1 port map( A => n88, ZN => n60);
   U92 : INV_X1 port map( A => n89, ZN => n61);
   U93 : INV_X1 port map( A => n97, ZN => n48);
   U94 : INV_X1 port map( A => n103, ZN => n52);
   U95 : INV_X1 port map( A => n87, ZN => n59);
   U96 : INV_X1 port map( A => n99, ZN => n50);
   U97 : INV_X1 port map( A => n105, ZN => n54);
   U98 : INV_X1 port map( A => n104, ZN => n53);
   U99 : INV_X1 port map( A => n95, ZN => n46);
   U100 : INV_X1 port map( A => n114, ZN => n57);
   U101 : AOI21_X1 port map( B1 => n82, B2 => A(9), A => n83, ZN => n81);
   U102 : OAI21_X1 port map( B1 => n84, B2 => n75, A => n82, ZN => SUM(8));
   U103 : AOI21_X1 port map( B1 => n57, B2 => A(7), A => n84, ZN => n85);
   U104 : OAI21_X1 port map( B1 => n86, B2 => n76, A => n57, ZN => SUM(6));
   U105 : OAI21_X1 port map( B1 => n87, B2 => n77, A => n58, ZN => SUM(5));
   U106 : OAI21_X1 port map( B1 => n88, B2 => n78, A => n59, ZN => SUM(4));
   U107 : OAI21_X1 port map( B1 => n89, B2 => n79, A => n60, ZN => SUM(3));
   U108 : XNOR2_X1 port map( A => A(30), B => n90, ZN => SUM(30));
   U109 : OAI21_X1 port map( B1 => n91, B2 => n80, A => n61, ZN => SUM(2));
   U110 : OAI21_X1 port map( B1 => n92, B2 => n65, A => n90, ZN => SUM(29));
   U111 : NAND2_X1 port map( A1 => n92, A2 => n65, ZN => n90);
   U112 : AOI21_X1 port map( B1 => n46, B2 => A(28), A => n92, ZN => n93);
   U113 : OAI21_X1 port map( B1 => n94, B2 => n10, A => n46, ZN => SUM(27));
   U114 : OAI21_X1 port map( B1 => n96, B2 => n66, A => n47, ZN => SUM(26));
   U115 : NOR2_X1 port map( A1 => n8, A2 => A(26), ZN => n94);
   U116 : OAI21_X1 port map( B1 => n97, B2 => n9, A => n8, ZN => SUM(25));
   U117 : OAI21_X1 port map( B1 => n98, B2 => n67, A => n48, ZN => SUM(24));
   U118 : NOR2_X1 port map( A1 => n49, A2 => A(24), ZN => n97);
   U119 : OAI21_X1 port map( B1 => n99, B2 => n7, A => n49, ZN => SUM(23));
   U120 : OAI21_X1 port map( B1 => n100, B2 => n68, A => n50, ZN => SUM(22));
   U121 : OAI21_X1 port map( B1 => n101, B2 => n2, A => n40, ZN => SUM(21));
   U122 : OAI21_X1 port map( B1 => n102, B2 => n69, A => n51, ZN => SUM(20));
   U123 : OAI21_X1 port map( B1 => n63, B2 => n64, A => n62, ZN => SUM(1));
   U124 : OAI21_X1 port map( B1 => n103, B2 => n12, A => n11, ZN => SUM(19));
   U125 : OAI21_X1 port map( B1 => n104, B2 => n70, A => n52, ZN => SUM(18));
   U126 : OAI21_X1 port map( B1 => n105, B2 => n15, A => n38, ZN => SUM(17));
   U127 : OAI21_X1 port map( B1 => n106, B2 => n71, A => n54, ZN => SUM(16));
   U128 : NOR2_X1 port map( A1 => n16, A2 => A(16), ZN => n105);
   U129 : OAI21_X1 port map( B1 => n107, B2 => n72, A => n16, ZN => SUM(15));
   U130 : NOR2_X1 port map( A1 => n4, A2 => A(15), ZN => n106);
   U131 : OAI21_X1 port map( B1 => n108, B2 => n21, A => n39, ZN => SUM(14));
   U132 : AOI21_X1 port map( B1 => n110, B2 => A(13), A => n108, ZN => n109);
   U133 : OAI21_X1 port map( B1 => n111, B2 => n73, A => n110, ZN => SUM(12));
   U134 : AOI21_X1 port map( B1 => n113, B2 => A(11), A => n111, ZN => n112);
   U135 : OAI21_X1 port map( B1 => n83, B2 => n74, A => n113, ZN => SUM(10));
   U136 : NOR2_X1 port map( A1 => n58, A2 => A(6), ZN => n114);
   U137 : NOR2_X1 port map( A1 => n60, A2 => A(4), ZN => n87);
   U138 : NOR2_X1 port map( A1 => n61, A2 => A(3), ZN => n88);
   U139 : NOR2_X1 port map( A1 => n62, A2 => A(2), ZN => n89);
   U140 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n91);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_63;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_62;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_61;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U4 : INV_X1 port map( A => n13, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_60;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : INV_X1 port map( A => n13, ZN => Y(3));
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_59;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : INV_X1 port map( A => n10, ZN => Y(0));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n1, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n1, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U9 : INV_X1 port map( A => n13, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_58;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n10, n11, n12, n13, n14 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(2));
   U2 : INV_X1 port map( A => n12, ZN => Y(1));
   U3 : BUF_X1 port map( A => SEL, Z => n1);
   U4 : INV_X1 port map( A => n11, ZN => Y(0));
   U5 : INV_X1 port map( A => SEL, ZN => n10);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n10, B1 => B(2), B2 => n1, ZN => 
                           n13);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n10, B1 => B(1), B2 => SEL, ZN => 
                           n12);
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n10, B1 => B(0), B2 => n1, ZN => 
                           n11);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n10, B1 => n1, B2 => B(3), ZN => 
                           n14);
   U10 : INV_X1 port map( A => n14, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_57;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(3));
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : INV_X1 port map( A => n10, ZN => Y(0));
   U4 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U5 : INV_X1 port map( A => n12, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_56;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n13, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_55;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_54;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_53;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_52;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_51;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_50;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_49;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_48;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U5 : INV_X1 port map( A => n10, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U7 : INV_X1 port map( A => SEL, ZN => n5);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_47;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_46;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n11, ZN => Y(1));
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : INV_X1 port map( A => n10, ZN => Y(0));
   U4 : INV_X1 port map( A => n13, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_45;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_44;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n11, ZN => Y(1));
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : INV_X1 port map( A => n10, ZN => Y(0));
   U4 : INV_X1 port map( A => n13, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_43;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6, n8 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : INV_X1 port map( A => n8, ZN => Y(2));
   U4 : INV_X1 port map( A => n6, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n6);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n8);
   U7 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_42;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_41;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_40;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_39;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_38;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_37;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_36;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_35;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_34;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => SEL, B2 => B(2), ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_33;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n10, n11, n12, n13, n14 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : INV_X1 port map( A => n12, ZN => Y(1));
   U3 : INV_X1 port map( A => n13, ZN => Y(2));
   U4 : INV_X1 port map( A => n14, ZN => Y(3));
   U5 : INV_X1 port map( A => n11, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n10, B1 => B(0), B2 => SEL, ZN => 
                           n11);
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n10, B1 => B(2), B2 => SEL, ZN => 
                           n13);
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n10, B1 => B(1), B2 => SEL, ZN => 
                           n12);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n10, B1 => B(3), B2 => n1, ZN => 
                           n14);
   U10 : INV_X1 port map( A => SEL, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_32;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U5 : INV_X1 port map( A => n10, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U7 : INV_X1 port map( A => SEL, ZN => n5);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_31;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_30;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_29;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => SEL, B2 => B(2), ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_28;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_27;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n8, n9, n10 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U2 : INV_X1 port map( A => n9, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n9);
   U4 : INV_X1 port map( A => n8, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n8);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A(3), B1 => B(3), B2 => SEL, ZN => 
                           n10);
   U7 : INV_X1 port map( A => SEL, ZN => n5);
   U8 : INV_X1 port map( A => n10, ZN => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_26;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_25;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_24;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_23;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_22;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_21;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_20;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_19;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_18;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_17;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n11, n12, n13, n14, n15 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : INV_X1 port map( A => n12, ZN => Y(0));
   U4 : AOI22_X1 port map( A1 => A(0), A2 => n11, B1 => B(0), B2 => SEL, ZN => 
                           n12);
   U5 : INV_X1 port map( A => n13, ZN => Y(1));
   U6 : AOI22_X1 port map( A1 => A(1), A2 => n11, B1 => B(1), B2 => SEL, ZN => 
                           n13);
   U7 : INV_X1 port map( A => n14, ZN => Y(2));
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n11, B1 => n1, B2 => B(2), ZN => 
                           n14);
   U9 : INV_X1 port map( A => n15, ZN => Y(3));
   U10 : INV_X1 port map( A => SEL, ZN => n11);
   U11 : AOI22_X1 port map( A1 => A(3), A2 => n11, B1 => n2, B2 => B(3), ZN => 
                           n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_16;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U5 : INV_X1 port map( A => n10, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U7 : INV_X1 port map( A => SEL, ZN => n5);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_15;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_14;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_13;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_12;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_11;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : INV_X1 port map( A => n13, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_10;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_9;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n13, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_8;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(3));
   U2 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U3 : INV_X1 port map( A => n12, ZN => Y(2));
   U4 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U5 : INV_X1 port map( A => n11, ZN => Y(1));
   U6 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U7 : INV_X1 port map( A => n10, ZN => Y(0));
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_7;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n13, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_6;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_5;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n13, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_4;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n13, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_3;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n11, ZN => Y(1));
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : INV_X1 port map( A => SEL, ZN => n5);
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U7 : INV_X1 port map( A => n13, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_2;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n11, ZN => Y(1));
   U3 : INV_X1 port map( A => n12, ZN => Y(2));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U5 : INV_X1 port map( A => n13, ZN => Y(3));
   U6 : INV_X1 port map( A => n10, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_1;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(2));
   U2 : INV_X1 port map( A => n10, ZN => Y(0));
   U3 : INV_X1 port map( A => n13, ZN => Y(3));
   U4 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n13);
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n10);
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n12);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n11);
   U8 : INV_X1 port map( A => SEL, ZN => n5);
   U9 : INV_X1 port map( A => n11, ZN => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_127 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_127;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_127 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_126 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_126;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_126 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_125 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_125;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_125 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_124 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_124;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_124 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_123 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_123;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_123 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_122 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_122;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_122 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_121 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_121;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_121 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_120 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_120;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_120 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_119 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_119;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_119 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_118 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_118;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_118 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_117 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_117;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_117 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_116 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_116;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_116 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_115 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_115;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_115 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_114 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_114;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_114 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_113 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_113;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_113 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_112 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_112;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_112 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_111 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_111;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_111 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_110 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_110;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_110 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_109 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_109;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_109 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_108 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_108;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_108 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_107 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_107;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_107 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_106 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_106;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_106 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_105 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_105;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_105 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_104 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_104;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_104 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_103 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_103;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_103 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_102 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_102;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_102 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_101 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_101;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_101 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_100 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_100;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_100 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_99 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_99;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_99 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_98 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_98;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_98 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_97 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_97;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_97 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_96 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_96;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_96 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_95 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_95;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_95 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_94 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_94;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_94 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_93 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_93;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_93 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_92 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_92;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_92 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_91 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_91;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_91 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_90 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_90;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_90 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_89 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_89;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_89 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_88 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_88;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_88 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_87 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_87;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_87 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_86 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_86;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_86 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_85 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_85;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_85 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_84 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_84;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_84 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_83 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_83;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_83 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_82 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_82;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_82 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_81 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_81;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_81 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_80 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_80;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_80 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_79 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_79;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_79 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_78 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_78;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_78 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_77 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_77;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_77 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_76 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_76;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_76 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_75 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_75;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_75 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_74 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_74;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_74 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_73 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_73;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_73 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_72 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_72;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_72 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_71 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_71;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_71 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_70 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_70;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_70 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_69 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_69;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_69 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_68 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_68;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_68 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_67 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_67;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_67 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_66 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_66;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_66 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_65 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_65;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_65 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_64 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_64;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_64 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_63;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_63 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_62;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_62 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_61;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_61 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_60;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_60 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_59;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_59 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_58;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_58 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_57;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_57 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_56;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_56 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_55;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_55 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_54;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_54 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_53;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_53 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_52;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_52 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_51;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_51 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_50;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_50 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_49;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_49 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_48;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_48 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_47;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_47 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_46;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_46 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_45;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_45 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_44;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_44 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_43;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_43 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_42;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_42 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_41;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_41 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_40;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_40 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_39;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_39 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_38;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_38 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_37;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_37 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_36;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_36 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_35;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_35 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_34;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_34 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_33;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_33 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_32;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_32 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_31;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_31 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_30;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_30 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_29;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_29 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_28;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_28 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_27;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_27 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_26;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_26 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_25;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_25 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_24;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_24 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_23;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_23 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_22;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_22 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_21;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_21 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_20;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_20 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_19;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_19 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_18;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_18 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_17;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_17 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_16;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_16 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_15;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_15 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_14;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_14 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_13;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_13 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_12;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_12 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_11;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_10;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_10 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_9;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_9 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_8;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_8 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_7;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_7 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_6;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_6 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_5;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_5 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_4;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_4 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_3;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_3 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_2;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_2 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_1;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_1 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_63;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_63 is

   component MUX2to1_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_125
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_126
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_126 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1006);
   RCA0 : RCAN_NBIT4_125 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1007);
   MUX21 : MUX2to1_NBIT4_63 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_62;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_62 is

   component MUX2to1_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_123
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_124
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_124 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1008);
   RCA0 : RCAN_NBIT4_123 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1009);
   MUX21 : MUX2to1_NBIT4_62 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_61;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_61 is

   component MUX2to1_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_121
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_122
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_122 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1010);
   RCA0 : RCAN_NBIT4_121 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1011);
   MUX21 : MUX2to1_NBIT4_61 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_60;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_60 is

   component MUX2to1_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_119
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_120
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_120 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1012);
   RCA0 : RCAN_NBIT4_119 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1013);
   MUX21 : MUX2to1_NBIT4_60 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_59;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_59 is

   component MUX2to1_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_117
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_118
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_118 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1014);
   RCA0 : RCAN_NBIT4_117 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1015);
   MUX21 : MUX2to1_NBIT4_59 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_58;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_58 is

   component MUX2to1_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_115
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_116
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1016, n_1017 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_116 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1016);
   RCA0 : RCAN_NBIT4_115 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1017);
   MUX21 : MUX2to1_NBIT4_58 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_57;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_57 is

   component MUX2to1_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_113
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_114
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1018, n_1019 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_114 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1018);
   RCA0 : RCAN_NBIT4_113 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1019);
   MUX21 : MUX2to1_NBIT4_57 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_56;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_56 is

   component MUX2to1_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_111
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_112
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1020, n_1021 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_112 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1020);
   RCA0 : RCAN_NBIT4_111 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1021);
   MUX21 : MUX2to1_NBIT4_56 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_55;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_55 is

   component MUX2to1_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_109
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_110
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1022, n_1023 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_110 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1022);
   RCA0 : RCAN_NBIT4_109 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1023);
   MUX21 : MUX2to1_NBIT4_55 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_54;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_54 is

   component MUX2to1_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_107
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_108
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1024, n_1025 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_108 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1024);
   RCA0 : RCAN_NBIT4_107 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1025);
   MUX21 : MUX2to1_NBIT4_54 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_53;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_53 is

   component MUX2to1_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_105
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_106
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1026, n_1027 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_106 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1026);
   RCA0 : RCAN_NBIT4_105 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1027);
   MUX21 : MUX2to1_NBIT4_53 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_52;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_52 is

   component MUX2to1_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_103
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_104
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1028, n_1029 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_104 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1028);
   RCA0 : RCAN_NBIT4_103 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1029);
   MUX21 : MUX2to1_NBIT4_52 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_51;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_51 is

   component MUX2to1_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_101
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_102
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1030, n_1031 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_102 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1030);
   RCA0 : RCAN_NBIT4_101 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1031);
   MUX21 : MUX2to1_NBIT4_51 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_50;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_50 is

   component MUX2to1_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_99
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_100
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1032, n_1033 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_100 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1032);
   RCA0 : RCAN_NBIT4_99 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1033);
   MUX21 : MUX2to1_NBIT4_50 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_49;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_49 is

   component MUX2to1_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_97
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_98
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1034, n_1035 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_98 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1034);
   RCA0 : RCAN_NBIT4_97 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1035);
   MUX21 : MUX2to1_NBIT4_49 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_48;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_48 is

   component MUX2to1_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_95
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_96
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1036, n_1037 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_96 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1036);
   RCA0 : RCAN_NBIT4_95 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1037);
   MUX21 : MUX2to1_NBIT4_48 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_47;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_47 is

   component MUX2to1_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_93
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_94
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1038, n_1039 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_94 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1038);
   RCA0 : RCAN_NBIT4_93 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1039);
   MUX21 : MUX2to1_NBIT4_47 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_46;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_46 is

   component MUX2to1_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_91
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_92
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1040, n_1041 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_92 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1040);
   RCA0 : RCAN_NBIT4_91 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1041);
   MUX21 : MUX2to1_NBIT4_46 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_45;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_45 is

   component MUX2to1_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_89
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_90
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1042, n_1043 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_90 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1042);
   RCA0 : RCAN_NBIT4_89 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1043);
   MUX21 : MUX2to1_NBIT4_45 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_44;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_44 is

   component MUX2to1_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_87
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_88
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1044, n_1045 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_88 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1044);
   RCA0 : RCAN_NBIT4_87 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1045);
   MUX21 : MUX2to1_NBIT4_44 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_43;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_43 is

   component MUX2to1_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_85
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_86
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1046, n_1047 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_86 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1046);
   RCA0 : RCAN_NBIT4_85 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1047);
   MUX21 : MUX2to1_NBIT4_43 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_42;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_42 is

   component MUX2to1_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_83
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_84
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1048, n_1049 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_84 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1048);
   RCA0 : RCAN_NBIT4_83 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1049);
   MUX21 : MUX2to1_NBIT4_42 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_41;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_41 is

   component MUX2to1_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_81
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_82
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1050, n_1051 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_82 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1050);
   RCA0 : RCAN_NBIT4_81 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1051);
   MUX21 : MUX2to1_NBIT4_41 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_40;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_40 is

   component MUX2to1_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_79
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_80
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1052, n_1053 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_80 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1052);
   RCA0 : RCAN_NBIT4_79 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1053);
   MUX21 : MUX2to1_NBIT4_40 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_39;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_39 is

   component MUX2to1_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_77
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_78
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1054, n_1055 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_78 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1054);
   RCA0 : RCAN_NBIT4_77 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1055);
   MUX21 : MUX2to1_NBIT4_39 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_38;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_38 is

   component MUX2to1_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_75
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_76
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1056, n_1057 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_76 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1056);
   RCA0 : RCAN_NBIT4_75 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1057);
   MUX21 : MUX2to1_NBIT4_38 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_37;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_37 is

   component MUX2to1_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_73
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_74
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1058, n_1059 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_74 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1058);
   RCA0 : RCAN_NBIT4_73 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1059);
   MUX21 : MUX2to1_NBIT4_37 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_36;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_36 is

   component MUX2to1_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_71
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_72
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1060, n_1061 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_72 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1060);
   RCA0 : RCAN_NBIT4_71 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1061);
   MUX21 : MUX2to1_NBIT4_36 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_35;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_35 is

   component MUX2to1_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_69
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_70
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1062, n_1063 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_70 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1062);
   RCA0 : RCAN_NBIT4_69 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1063);
   MUX21 : MUX2to1_NBIT4_35 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_34;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_34 is

   component MUX2to1_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_67
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_68
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1064, n_1065 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_68 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1064);
   RCA0 : RCAN_NBIT4_67 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1065);
   MUX21 : MUX2to1_NBIT4_34 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_33;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_33 is

   component MUX2to1_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_65
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_66
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1066, n_1067 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_66 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1066);
   RCA0 : RCAN_NBIT4_65 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1067);
   MUX21 : MUX2to1_NBIT4_33 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_32;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_32 is

   component MUX2to1_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_64
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1068, n_1069 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_64 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1068);
   RCA0 : RCAN_NBIT4_63 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1069);
   MUX21 : MUX2to1_NBIT4_32 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_31;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_31 is

   component MUX2to1_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1070, n_1071 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_62 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1070);
   RCA0 : RCAN_NBIT4_61 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1071);
   MUX21 : MUX2to1_NBIT4_31 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_30;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_30 is

   component MUX2to1_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1072, n_1073 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_60 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1072);
   RCA0 : RCAN_NBIT4_59 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1073);
   MUX21 : MUX2to1_NBIT4_30 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_29;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_29 is

   component MUX2to1_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1074, n_1075 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_58 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1074);
   RCA0 : RCAN_NBIT4_57 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1075);
   MUX21 : MUX2to1_NBIT4_29 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_28;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_28 is

   component MUX2to1_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1076, n_1077 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1076);
   RCA0 : RCAN_NBIT4_55 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1077);
   MUX21 : MUX2to1_NBIT4_28 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_27;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_27 is

   component MUX2to1_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1078, n_1079 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_54 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1078);
   RCA0 : RCAN_NBIT4_53 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1079);
   MUX21 : MUX2to1_NBIT4_27 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_26;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_26 is

   component MUX2to1_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1080, n_1081 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_52 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1080);
   RCA0 : RCAN_NBIT4_51 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1081);
   MUX21 : MUX2to1_NBIT4_26 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_25;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_25 is

   component MUX2to1_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1082, n_1083 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_50 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1082);
   RCA0 : RCAN_NBIT4_49 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1083);
   MUX21 : MUX2to1_NBIT4_25 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_24;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_24 is

   component MUX2to1_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1084, n_1085 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1084);
   RCA0 : RCAN_NBIT4_47 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1085);
   MUX21 : MUX2to1_NBIT4_24 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_23;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_23 is

   component MUX2to1_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1086, n_1087 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_46 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1086);
   RCA0 : RCAN_NBIT4_45 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1087);
   MUX21 : MUX2to1_NBIT4_23 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_22;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_22 is

   component MUX2to1_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1088, n_1089 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_44 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1088);
   RCA0 : RCAN_NBIT4_43 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1089);
   MUX21 : MUX2to1_NBIT4_22 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_21;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_21 is

   component MUX2to1_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1090, n_1091 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_42 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1090);
   RCA0 : RCAN_NBIT4_41 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1091);
   MUX21 : MUX2to1_NBIT4_21 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_20;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_20 is

   component MUX2to1_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1092, n_1093 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1092);
   RCA0 : RCAN_NBIT4_39 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1093);
   MUX21 : MUX2to1_NBIT4_20 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_19;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_19 is

   component MUX2to1_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1094, n_1095 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_38 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1094);
   RCA0 : RCAN_NBIT4_37 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1095);
   MUX21 : MUX2to1_NBIT4_19 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_18;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_18 is

   component MUX2to1_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1096, n_1097 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_36 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1096);
   RCA0 : RCAN_NBIT4_35 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1097);
   MUX21 : MUX2to1_NBIT4_18 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_17;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_17 is

   component MUX2to1_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1098, n_1099 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_34 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1098);
   RCA0 : RCAN_NBIT4_33 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1099);
   MUX21 : MUX2to1_NBIT4_17 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_16;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_16 is

   component MUX2to1_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1100, n_1101 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1100);
   RCA0 : RCAN_NBIT4_31 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1101);
   MUX21 : MUX2to1_NBIT4_16 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_15;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_15 is

   component MUX2to1_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1102, n_1103 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1102);
   RCA0 : RCAN_NBIT4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1103);
   MUX21 : MUX2to1_NBIT4_15 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_14;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_14 is

   component MUX2to1_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1104, n_1105 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1104);
   RCA0 : RCAN_NBIT4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1105);
   MUX21 : MUX2to1_NBIT4_14 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_13;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_13 is

   component MUX2to1_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1106, n_1107 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1106);
   RCA0 : RCAN_NBIT4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1107);
   MUX21 : MUX2to1_NBIT4_13 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_12;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_12 is

   component MUX2to1_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1108, n_1109 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1108);
   RCA0 : RCAN_NBIT4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1109);
   MUX21 : MUX2to1_NBIT4_12 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_11;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_11 is

   component MUX2to1_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1110, n_1111 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1110);
   RCA0 : RCAN_NBIT4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1111);
   MUX21 : MUX2to1_NBIT4_11 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_10;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_10 is

   component MUX2to1_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1112, n_1113 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1112);
   RCA0 : RCAN_NBIT4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1113);
   MUX21 : MUX2to1_NBIT4_10 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_9;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_9 is

   component MUX2to1_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1114, n_1115 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1114);
   RCA0 : RCAN_NBIT4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1115);
   MUX21 : MUX2to1_NBIT4_9 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_8;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_8 is

   component MUX2to1_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1116, n_1117 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1116);
   RCA0 : RCAN_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1117);
   MUX21 : MUX2to1_NBIT4_8 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_7;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_7 is

   component MUX2to1_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1118, n_1119 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1118);
   RCA0 : RCAN_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1119);
   MUX21 : MUX2to1_NBIT4_7 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_6;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_6 is

   component MUX2to1_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1120, n_1121 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1120);
   RCA0 : RCAN_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1121);
   MUX21 : MUX2to1_NBIT4_6 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_5;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_5 is

   component MUX2to1_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1122, n_1123 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1122);
   RCA0 : RCAN_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1123);
   MUX21 : MUX2to1_NBIT4_5 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_4;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_4 is

   component MUX2to1_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1124, n_1125 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1124);
   RCA0 : RCAN_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1125);
   MUX21 : MUX2to1_NBIT4_4 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_3;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_3 is

   component MUX2to1_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1126, n_1127 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1126);
   RCA0 : RCAN_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1127);
   MUX21 : MUX2to1_NBIT4_3 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_2;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_2 is

   component MUX2to1_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1128, n_1129 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1128);
   RCA0 : RCAN_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1129);
   MUX21 : MUX2to1_NBIT4_2 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_1;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_1 is

   component MUX2to1_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1130, n_1131 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1130);
   RCA0 : RCAN_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S0_3_port
                           , S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1131);
   MUX21 : MUX2to1_NBIT4_1 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_215 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_215;

architecture SYN_BEHAVIORAL of PG_block_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_214 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_214;

architecture SYN_BEHAVIORAL of PG_block_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_213 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_213;

architecture SYN_BEHAVIORAL of PG_block_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_212 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_212;

architecture SYN_BEHAVIORAL of PG_block_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_211 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_211;

architecture SYN_BEHAVIORAL of PG_block_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_210 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_210;

architecture SYN_BEHAVIORAL of PG_block_210 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_209 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_209;

architecture SYN_BEHAVIORAL of PG_block_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_208 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_208;

architecture SYN_BEHAVIORAL of PG_block_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_207 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_207;

architecture SYN_BEHAVIORAL of PG_block_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_206 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_206;

architecture SYN_BEHAVIORAL of PG_block_206 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_205 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_205;

architecture SYN_BEHAVIORAL of PG_block_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_204 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_204;

architecture SYN_BEHAVIORAL of PG_block_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_203 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_203;

architecture SYN_BEHAVIORAL of PG_block_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_202 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_202;

architecture SYN_BEHAVIORAL of PG_block_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_201 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_201;

architecture SYN_BEHAVIORAL of PG_block_201 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_200 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_200;

architecture SYN_BEHAVIORAL of PG_block_200 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_199 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_199;

architecture SYN_BEHAVIORAL of PG_block_199 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_198 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_198;

architecture SYN_BEHAVIORAL of PG_block_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_197 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_197;

architecture SYN_BEHAVIORAL of PG_block_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_196 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_196;

architecture SYN_BEHAVIORAL of PG_block_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_195 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_195;

architecture SYN_BEHAVIORAL of PG_block_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_194 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_194;

architecture SYN_BEHAVIORAL of PG_block_194 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_193 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_193;

architecture SYN_BEHAVIORAL of PG_block_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_192 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_192;

architecture SYN_BEHAVIORAL of PG_block_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_191 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_191;

architecture SYN_BEHAVIORAL of PG_block_191 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_190 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_190;

architecture SYN_BEHAVIORAL of PG_block_190 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_189 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_189;

architecture SYN_BEHAVIORAL of PG_block_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_188 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_188;

architecture SYN_BEHAVIORAL of PG_block_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_187 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_187;

architecture SYN_BEHAVIORAL of PG_block_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_186 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_186;

architecture SYN_BEHAVIORAL of PG_block_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_185 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_185;

architecture SYN_BEHAVIORAL of PG_block_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_184 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_184;

architecture SYN_BEHAVIORAL of PG_block_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_183 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_183;

architecture SYN_BEHAVIORAL of PG_block_183 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_182 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_182;

architecture SYN_BEHAVIORAL of PG_block_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_181 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_181;

architecture SYN_BEHAVIORAL of PG_block_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_180 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_180;

architecture SYN_BEHAVIORAL of PG_block_180 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_179 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_179;

architecture SYN_BEHAVIORAL of PG_block_179 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_178 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_178;

architecture SYN_BEHAVIORAL of PG_block_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_177 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_177;

architecture SYN_BEHAVIORAL of PG_block_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_176 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_176;

architecture SYN_BEHAVIORAL of PG_block_176 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_175 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_175;

architecture SYN_BEHAVIORAL of PG_block_175 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_174 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_174;

architecture SYN_BEHAVIORAL of PG_block_174 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_173 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_173;

architecture SYN_BEHAVIORAL of PG_block_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_172 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_172;

architecture SYN_BEHAVIORAL of PG_block_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_171 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_171;

architecture SYN_BEHAVIORAL of PG_block_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_170 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_170;

architecture SYN_BEHAVIORAL of PG_block_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_169 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_169;

architecture SYN_BEHAVIORAL of PG_block_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_168 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_168;

architecture SYN_BEHAVIORAL of PG_block_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_167 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_167;

architecture SYN_BEHAVIORAL of PG_block_167 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_166 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_166;

architecture SYN_BEHAVIORAL of PG_block_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_165 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_165;

architecture SYN_BEHAVIORAL of PG_block_165 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_164 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_164;

architecture SYN_BEHAVIORAL of PG_block_164 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_163 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_163;

architecture SYN_BEHAVIORAL of PG_block_163 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_162 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_162;

architecture SYN_BEHAVIORAL of PG_block_162 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_161 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_161;

architecture SYN_BEHAVIORAL of PG_block_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_160 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_160;

architecture SYN_BEHAVIORAL of PG_block_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_159 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_159;

architecture SYN_BEHAVIORAL of PG_block_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_158 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_158;

architecture SYN_BEHAVIORAL of PG_block_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_157 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_157;

architecture SYN_BEHAVIORAL of PG_block_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_156 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_156;

architecture SYN_BEHAVIORAL of PG_block_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_155 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_155;

architecture SYN_BEHAVIORAL of PG_block_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_154 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_154;

architecture SYN_BEHAVIORAL of PG_block_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_153 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_153;

architecture SYN_BEHAVIORAL of PG_block_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_152 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_152;

architecture SYN_BEHAVIORAL of PG_block_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_151 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_151;

architecture SYN_BEHAVIORAL of PG_block_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_150 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_150;

architecture SYN_BEHAVIORAL of PG_block_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_149 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_149;

architecture SYN_BEHAVIORAL of PG_block_149 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_148 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_148;

architecture SYN_BEHAVIORAL of PG_block_148 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_147 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_147;

architecture SYN_BEHAVIORAL of PG_block_147 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_146 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_146;

architecture SYN_BEHAVIORAL of PG_block_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_145 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_145;

architecture SYN_BEHAVIORAL of PG_block_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_144 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_144;

architecture SYN_BEHAVIORAL of PG_block_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_143 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_143;

architecture SYN_BEHAVIORAL of PG_block_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_142 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_142;

architecture SYN_BEHAVIORAL of PG_block_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_141 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_141;

architecture SYN_BEHAVIORAL of PG_block_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_140 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_140;

architecture SYN_BEHAVIORAL of PG_block_140 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_139 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_139;

architecture SYN_BEHAVIORAL of PG_block_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_138 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_138;

architecture SYN_BEHAVIORAL of PG_block_138 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_137 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_137;

architecture SYN_BEHAVIORAL of PG_block_137 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_136 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_136;

architecture SYN_BEHAVIORAL of PG_block_136 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_135 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_135;

architecture SYN_BEHAVIORAL of PG_block_135 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_134 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_134;

architecture SYN_BEHAVIORAL of PG_block_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_133 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_133;

architecture SYN_BEHAVIORAL of PG_block_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_132 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_132;

architecture SYN_BEHAVIORAL of PG_block_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_131 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_131;

architecture SYN_BEHAVIORAL of PG_block_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_130 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_130;

architecture SYN_BEHAVIORAL of PG_block_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_129 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_129;

architecture SYN_BEHAVIORAL of PG_block_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_128 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_128;

architecture SYN_BEHAVIORAL of PG_block_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_127 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_127;

architecture SYN_BEHAVIORAL of PG_block_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_126 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_126;

architecture SYN_BEHAVIORAL of PG_block_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_125 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_125;

architecture SYN_BEHAVIORAL of PG_block_125 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_124 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_124;

architecture SYN_BEHAVIORAL of PG_block_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_123 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_123;

architecture SYN_BEHAVIORAL of PG_block_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_122 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_122;

architecture SYN_BEHAVIORAL of PG_block_122 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_121 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_121;

architecture SYN_BEHAVIORAL of PG_block_121 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_120 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_120;

architecture SYN_BEHAVIORAL of PG_block_120 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_119 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_119;

architecture SYN_BEHAVIORAL of PG_block_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_118 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_118;

architecture SYN_BEHAVIORAL of PG_block_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_117 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_117;

architecture SYN_BEHAVIORAL of PG_block_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_116 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_116;

architecture SYN_BEHAVIORAL of PG_block_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_115 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_115;

architecture SYN_BEHAVIORAL of PG_block_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_114 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_114;

architecture SYN_BEHAVIORAL of PG_block_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_113 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_113;

architecture SYN_BEHAVIORAL of PG_block_113 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_112 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_112;

architecture SYN_BEHAVIORAL of PG_block_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n2, A2 => A(0), ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(1), ZN => n2);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_111 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_111;

architecture SYN_BEHAVIORAL of PG_block_111 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_110 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_110;

architecture SYN_BEHAVIORAL of PG_block_110 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_109 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_109;

architecture SYN_BEHAVIORAL of PG_block_109 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_108 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_108;

architecture SYN_BEHAVIORAL of PG_block_108 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_107 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_107;

architecture SYN_BEHAVIORAL of PG_block_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_106 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_106;

architecture SYN_BEHAVIORAL of PG_block_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_105 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_105;

architecture SYN_BEHAVIORAL of PG_block_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_104 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_104;

architecture SYN_BEHAVIORAL of PG_block_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_103 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_103;

architecture SYN_BEHAVIORAL of PG_block_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_102 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_102;

architecture SYN_BEHAVIORAL of PG_block_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_101 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_101;

architecture SYN_BEHAVIORAL of PG_block_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_100 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_100;

architecture SYN_BEHAVIORAL of PG_block_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_99 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_99;

architecture SYN_BEHAVIORAL of PG_block_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_98 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_98;

architecture SYN_BEHAVIORAL of PG_block_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_97 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_97;

architecture SYN_BEHAVIORAL of PG_block_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_96 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_96;

architecture SYN_BEHAVIORAL of PG_block_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_95 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_95;

architecture SYN_BEHAVIORAL of PG_block_95 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_94 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_94;

architecture SYN_BEHAVIORAL of PG_block_94 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_93 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_93;

architecture SYN_BEHAVIORAL of PG_block_93 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_92 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_92;

architecture SYN_BEHAVIORAL of PG_block_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_91 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_91;

architecture SYN_BEHAVIORAL of PG_block_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_90 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_90;

architecture SYN_BEHAVIORAL of PG_block_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_89 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_89;

architecture SYN_BEHAVIORAL of PG_block_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_88 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_88;

architecture SYN_BEHAVIORAL of PG_block_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_87 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_87;

architecture SYN_BEHAVIORAL of PG_block_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_86 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_86;

architecture SYN_BEHAVIORAL of PG_block_86 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_85 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_85;

architecture SYN_BEHAVIORAL of PG_block_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_84 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_84;

architecture SYN_BEHAVIORAL of PG_block_84 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_83 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_83;

architecture SYN_BEHAVIORAL of PG_block_83 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_82 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_82;

architecture SYN_BEHAVIORAL of PG_block_82 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_81 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_81;

architecture SYN_BEHAVIORAL of PG_block_81 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_80 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_80;

architecture SYN_BEHAVIORAL of PG_block_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_79 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_79;

architecture SYN_BEHAVIORAL of PG_block_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_78 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_78;

architecture SYN_BEHAVIORAL of PG_block_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_77 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_77;

architecture SYN_BEHAVIORAL of PG_block_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_76 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_76;

architecture SYN_BEHAVIORAL of PG_block_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_75 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_75;

architecture SYN_BEHAVIORAL of PG_block_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_74 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_74;

architecture SYN_BEHAVIORAL of PG_block_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_73 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_73;

architecture SYN_BEHAVIORAL of PG_block_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_72 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_72;

architecture SYN_BEHAVIORAL of PG_block_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_71 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_71;

architecture SYN_BEHAVIORAL of PG_block_71 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => A(1), B2 => B(0), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_70 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_70;

architecture SYN_BEHAVIORAL of PG_block_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_69 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_69;

architecture SYN_BEHAVIORAL of PG_block_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_68 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_68;

architecture SYN_BEHAVIORAL of PG_block_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_67 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_67;

architecture SYN_BEHAVIORAL of PG_block_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_66 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_66;

architecture SYN_BEHAVIORAL of PG_block_66 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_65 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_65;

architecture SYN_BEHAVIORAL of PG_block_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_64 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_64;

architecture SYN_BEHAVIORAL of PG_block_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_63 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_63;

architecture SYN_BEHAVIORAL of PG_block_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_62 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_62;

architecture SYN_BEHAVIORAL of PG_block_62 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_61 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_61;

architecture SYN_BEHAVIORAL of PG_block_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_60 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_60;

architecture SYN_BEHAVIORAL of PG_block_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_59 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_59;

architecture SYN_BEHAVIORAL of PG_block_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_58 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_58;

architecture SYN_BEHAVIORAL of PG_block_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_57 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_57;

architecture SYN_BEHAVIORAL of PG_block_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_56 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_56;

architecture SYN_BEHAVIORAL of PG_block_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_55 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_55;

architecture SYN_BEHAVIORAL of PG_block_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_54 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_54;

architecture SYN_BEHAVIORAL of PG_block_54 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_53 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_53;

architecture SYN_BEHAVIORAL of PG_block_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_52 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_52;

architecture SYN_BEHAVIORAL of PG_block_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_51 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_51;

architecture SYN_BEHAVIORAL of PG_block_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_50 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_50;

architecture SYN_BEHAVIORAL of PG_block_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_49 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_49;

architecture SYN_BEHAVIORAL of PG_block_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_48 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_48;

architecture SYN_BEHAVIORAL of PG_block_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_47 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_47;

architecture SYN_BEHAVIORAL of PG_block_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_46 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_46;

architecture SYN_BEHAVIORAL of PG_block_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_45 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_45;

architecture SYN_BEHAVIORAL of PG_block_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_44 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_44;

architecture SYN_BEHAVIORAL of PG_block_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_43 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_43;

architecture SYN_BEHAVIORAL of PG_block_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_42 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_42;

architecture SYN_BEHAVIORAL of PG_block_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_41 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_41;

architecture SYN_BEHAVIORAL of PG_block_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_40 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_40;

architecture SYN_BEHAVIORAL of PG_block_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_39 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_39;

architecture SYN_BEHAVIORAL of PG_block_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_38 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_38;

architecture SYN_BEHAVIORAL of PG_block_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_37 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_37;

architecture SYN_BEHAVIORAL of PG_block_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_36 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_36;

architecture SYN_BEHAVIORAL of PG_block_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_35 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_35;

architecture SYN_BEHAVIORAL of PG_block_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_34 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_34;

architecture SYN_BEHAVIORAL of PG_block_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_33 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_33;

architecture SYN_BEHAVIORAL of PG_block_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_32 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_32;

architecture SYN_BEHAVIORAL of PG_block_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_31 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_31;

architecture SYN_BEHAVIORAL of PG_block_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_30 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_30;

architecture SYN_BEHAVIORAL of PG_block_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_29 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_29;

architecture SYN_BEHAVIORAL of PG_block_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_28 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_28;

architecture SYN_BEHAVIORAL of PG_block_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_27 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_27;

architecture SYN_BEHAVIORAL of PG_block_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_26 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_26;

architecture SYN_BEHAVIORAL of PG_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_25 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_25;

architecture SYN_BEHAVIORAL of PG_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_24 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_24;

architecture SYN_BEHAVIORAL of PG_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_23 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_23;

architecture SYN_BEHAVIORAL of PG_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_22 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_22;

architecture SYN_BEHAVIORAL of PG_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_21 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_21;

architecture SYN_BEHAVIORAL of PG_block_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_20 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_20;

architecture SYN_BEHAVIORAL of PG_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_19 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_19;

architecture SYN_BEHAVIORAL of PG_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_18 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_18;

architecture SYN_BEHAVIORAL of PG_block_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_17 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_17;

architecture SYN_BEHAVIORAL of PG_block_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_16 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_16;

architecture SYN_BEHAVIORAL of PG_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_15 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_15;

architecture SYN_BEHAVIORAL of PG_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_14 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_14;

architecture SYN_BEHAVIORAL of PG_block_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_13 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_13;

architecture SYN_BEHAVIORAL of PG_block_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_12 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_12;

architecture SYN_BEHAVIORAL of PG_block_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_11 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_11;

architecture SYN_BEHAVIORAL of PG_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_10 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_10;

architecture SYN_BEHAVIORAL of PG_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_9 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_9;

architecture SYN_BEHAVIORAL of PG_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_8 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_8;

architecture SYN_BEHAVIORAL of PG_block_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_7 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_7;

architecture SYN_BEHAVIORAL of PG_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_6 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_6;

architecture SYN_BEHAVIORAL of PG_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U3 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_5 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_5;

architecture SYN_BEHAVIORAL of PG_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_4 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_4;

architecture SYN_BEHAVIORAL of PG_block_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : INV_X1 port map( A => n3, ZN => PGout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_3 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_3;

architecture SYN_BEHAVIORAL of PG_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_2 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_2;

architecture SYN_BEHAVIORAL of PG_block_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n3, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_1 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_1;

architecture SYN_BEHAVIORAL of PG_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PGout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_71 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_71;

architecture SYN_BEHAVIORAL of G_block_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_70 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_70;

architecture SYN_BEHAVIORAL of G_block_70 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_69 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_69;

architecture SYN_BEHAVIORAL of G_block_69 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_68 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_68;

architecture SYN_BEHAVIORAL of G_block_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_67 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_67;

architecture SYN_BEHAVIORAL of G_block_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_66 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_66;

architecture SYN_BEHAVIORAL of G_block_66 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_65 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_65;

architecture SYN_BEHAVIORAL of G_block_65 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_64 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_64;

architecture SYN_BEHAVIORAL of G_block_64 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_63 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_63;

architecture SYN_BEHAVIORAL of G_block_63 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_62 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_62;

architecture SYN_BEHAVIORAL of G_block_62 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_61 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_61;

architecture SYN_BEHAVIORAL of G_block_61 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_60 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_60;

architecture SYN_BEHAVIORAL of G_block_60 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_59 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_59;

architecture SYN_BEHAVIORAL of G_block_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_58 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_58;

architecture SYN_BEHAVIORAL of G_block_58 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_57 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_57;

architecture SYN_BEHAVIORAL of G_block_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_56 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_56;

architecture SYN_BEHAVIORAL of G_block_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_55 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_55;

architecture SYN_BEHAVIORAL of G_block_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_54 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_54;

architecture SYN_BEHAVIORAL of G_block_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_53 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_53;

architecture SYN_BEHAVIORAL of G_block_53 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_52 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_52;

architecture SYN_BEHAVIORAL of G_block_52 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_51 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_51;

architecture SYN_BEHAVIORAL of G_block_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_50 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_50;

architecture SYN_BEHAVIORAL of G_block_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_49 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_49;

architecture SYN_BEHAVIORAL of G_block_49 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_48 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_48;

architecture SYN_BEHAVIORAL of G_block_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_47 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_47;

architecture SYN_BEHAVIORAL of G_block_47 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_46 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_46;

architecture SYN_BEHAVIORAL of G_block_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_45 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_45;

architecture SYN_BEHAVIORAL of G_block_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_44 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_44;

architecture SYN_BEHAVIORAL of G_block_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_43 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_43;

architecture SYN_BEHAVIORAL of G_block_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_42 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_42;

architecture SYN_BEHAVIORAL of G_block_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_41 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_41;

architecture SYN_BEHAVIORAL of G_block_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X2 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_40 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_40;

architecture SYN_BEHAVIORAL of G_block_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_39 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_39;

architecture SYN_BEHAVIORAL of G_block_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_38 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_38;

architecture SYN_BEHAVIORAL of G_block_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Gout);
   U2 : NAND2_X1 port map( A1 => B, A2 => A(1), ZN => n2);
   U3 : INV_X1 port map( A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_37 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_37;

architecture SYN_BEHAVIORAL of G_block_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_36 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_36;

architecture SYN_BEHAVIORAL of G_block_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_35 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_35;

architecture SYN_BEHAVIORAL of G_block_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_34 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_34;

architecture SYN_BEHAVIORAL of G_block_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_33 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_33;

architecture SYN_BEHAVIORAL of G_block_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_32 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_32;

architecture SYN_BEHAVIORAL of G_block_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_31 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_31;

architecture SYN_BEHAVIORAL of G_block_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_30 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_30;

architecture SYN_BEHAVIORAL of G_block_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_29 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_29;

architecture SYN_BEHAVIORAL of G_block_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_28 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_28;

architecture SYN_BEHAVIORAL of G_block_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_27 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_27;

architecture SYN_BEHAVIORAL of G_block_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_26 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_26;

architecture SYN_BEHAVIORAL of G_block_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_25 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_25;

architecture SYN_BEHAVIORAL of G_block_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_24 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_24;

architecture SYN_BEHAVIORAL of G_block_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_23 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_23;

architecture SYN_BEHAVIORAL of G_block_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_22 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_22;

architecture SYN_BEHAVIORAL of G_block_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_21 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_21;

architecture SYN_BEHAVIORAL of G_block_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_20 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_20;

architecture SYN_BEHAVIORAL of G_block_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => Gout);
   U2 : INV_X1 port map( A => B, ZN => n1);
   U3 : INV_X1 port map( A => A(1), ZN => n2);
   U4 : INV_X1 port map( A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_19 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_19;

architecture SYN_BEHAVIORAL of G_block_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_18 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_18;

architecture SYN_BEHAVIORAL of G_block_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_17 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_17;

architecture SYN_BEHAVIORAL of G_block_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_16 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_16;

architecture SYN_BEHAVIORAL of G_block_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_15 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_15;

architecture SYN_BEHAVIORAL of G_block_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_14 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_14;

architecture SYN_BEHAVIORAL of G_block_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_13 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_13;

architecture SYN_BEHAVIORAL of G_block_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_12 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_12;

architecture SYN_BEHAVIORAL of G_block_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_11 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_11;

architecture SYN_BEHAVIORAL of G_block_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_10 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_10;

architecture SYN_BEHAVIORAL of G_block_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_9 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_9;

architecture SYN_BEHAVIORAL of G_block_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_8 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_8;

architecture SYN_BEHAVIORAL of G_block_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_7 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_7;

architecture SYN_BEHAVIORAL of G_block_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_6 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_6;

architecture SYN_BEHAVIORAL of G_block_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_5 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_5;

architecture SYN_BEHAVIORAL of G_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_4 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_4;

architecture SYN_BEHAVIORAL of G_block_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_3 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_3;

architecture SYN_BEHAVIORAL of G_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_2 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_2;

architecture SYN_BEHAVIORAL of G_block_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => Gout);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_1 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_1;

architecture SYN_BEHAVIORAL of G_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_7;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U2 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U3 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U4 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U5 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U6 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U7 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U8 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U9 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U10 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U11 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U14 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U18 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U20 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U21 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U22 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U23 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U24 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U25 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U26 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U27 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U28 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U29 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U30 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_6;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U2 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U3 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U4 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U5 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U6 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U7 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U8 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U9 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U10 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U11 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U12 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U13 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U14 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U15 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U18 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U19 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U20 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U21 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U22 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U23 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U24 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U25 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U26 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U27 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U28 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U29 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U30 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U31 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_5;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : INV_X1 port map( A => B(21), ZN => n1);
   U2 : INV_X1 port map( A => B(23), ZN => n2);
   U3 : XNOR2_X1 port map( A => n1, B => A(21), ZN => Pout(21));
   U4 : XNOR2_X1 port map( A => n2, B => A(23), ZN => Pout(23));
   U5 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U6 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U7 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U8 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U9 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U10 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U11 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U12 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U13 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U14 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U15 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U16 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U17 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U18 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U19 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U20 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U21 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U22 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U23 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U24 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U25 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U26 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U27 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U28 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U29 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U30 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U31 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U49 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U51 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U65 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U66 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_4;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U3 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U4 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U5 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U6 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U7 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U8 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U9 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U10 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U11 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U12 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U13 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U14 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U15 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U16 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U17 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U18 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U19 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U20 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U21 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U22 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U23 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U24 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U25 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U26 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U27 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U28 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U29 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U30 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_3;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : INV_X1 port map( A => B(23), ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => A(23), ZN => Pout(23));
   U3 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U4 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U5 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U6 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U7 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U8 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U9 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U10 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U11 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U12 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U13 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U14 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U15 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U16 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U17 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U18 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U19 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U20 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U21 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U22 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U23 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U24 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U25 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U26 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U27 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U28 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U29 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U30 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U31 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U32 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U49 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U65 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_2;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U2 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U3 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U4 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U5 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U6 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U7 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U8 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U9 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U10 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U11 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U12 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U13 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U14 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U15 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U18 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U19 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U20 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U21 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U22 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U23 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U24 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U25 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U26 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U27 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U28 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U29 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U30 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U31 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U32 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_1;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U2 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U3 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U4 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U5 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U6 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U7 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U8 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U9 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U10 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U11 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U12 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U14 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U15 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U16 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U18 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U19 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U20 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U21 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U22 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U23 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U24 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U25 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U26 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U27 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U28 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));
   U29 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U30 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U31 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U32 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_7 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_7;

architecture SYN_BEHAVIORAL of ENCODER_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_6 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_6;

architecture SYN_BEHAVIORAL of ENCODER_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_5 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_5;

architecture SYN_BEHAVIORAL of ENCODER_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_4 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_4;

architecture SYN_BEHAVIORAL of ENCODER_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_3 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_3;

architecture SYN_BEHAVIORAL of ENCODER_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_2 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_2;

architecture SYN_BEHAVIORAL of ENCODER_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_1 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_1;

architecture SYN_BEHAVIORAL of ENCODER_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n7);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => OUTPUT(1));
   U3 : INV_X1 port map( A => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U5 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n6, ZN => OUTPUT(0));
   U6 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_31 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_31;

architecture SYN_ARCH1 of ND4_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_30 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_30;

architecture SYN_ARCH1 of ND4_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_29 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_29;

architecture SYN_ARCH1 of ND4_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_28 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_28;

architecture SYN_ARCH1 of ND4_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_27 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_27;

architecture SYN_ARCH1 of ND4_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_26 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_26;

architecture SYN_ARCH1 of ND4_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_25 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_25;

architecture SYN_ARCH1 of ND4_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_24 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_24;

architecture SYN_ARCH1 of ND4_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_23 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_23;

architecture SYN_ARCH1 of ND4_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_22 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_22;

architecture SYN_ARCH1 of ND4_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_21 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_21;

architecture SYN_ARCH1 of ND4_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_20 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_20;

architecture SYN_ARCH1 of ND4_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_19 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_19;

architecture SYN_ARCH1 of ND4_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_18 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_18;

architecture SYN_ARCH1 of ND4_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_17 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_17;

architecture SYN_ARCH1 of ND4_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_16 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_16;

architecture SYN_ARCH1 of ND4_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_15 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_15;

architecture SYN_ARCH1 of ND4_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_14 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_14;

architecture SYN_ARCH1 of ND4_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_13 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_13;

architecture SYN_ARCH1 of ND4_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_12 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_12;

architecture SYN_ARCH1 of ND4_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_11 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_11;

architecture SYN_ARCH1 of ND4_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_10 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_10;

architecture SYN_ARCH1 of ND4_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_9 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_9;

architecture SYN_ARCH1 of ND4_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_8 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_8;

architecture SYN_ARCH1 of ND4_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_7 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_7;

architecture SYN_ARCH1 of ND4_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_6 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_6;

architecture SYN_ARCH1 of ND4_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_5 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_5;

architecture SYN_ARCH1 of ND4_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_4 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_4;

architecture SYN_ARCH1 of ND4_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_3 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_3;

architecture SYN_ARCH1 of ND4_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_2 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_2;

architecture SYN_ARCH1 of ND4_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_1 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_1;

architecture SYN_ARCH1 of ND4_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_127 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_127;

architecture SYN_ARCH1 of ND3_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_126 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_126;

architecture SYN_ARCH1 of ND3_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_125 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_125;

architecture SYN_ARCH1 of ND3_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_124 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_124;

architecture SYN_ARCH1 of ND3_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_123 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_123;

architecture SYN_ARCH1 of ND3_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_122 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_122;

architecture SYN_ARCH1 of ND3_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_121 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_121;

architecture SYN_ARCH1 of ND3_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_120 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_120;

architecture SYN_ARCH1 of ND3_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_119 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_119;

architecture SYN_ARCH1 of ND3_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_118 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_118;

architecture SYN_ARCH1 of ND3_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_117 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_117;

architecture SYN_ARCH1 of ND3_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_116 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_116;

architecture SYN_ARCH1 of ND3_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_115 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_115;

architecture SYN_ARCH1 of ND3_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_114 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_114;

architecture SYN_ARCH1 of ND3_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_113 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_113;

architecture SYN_ARCH1 of ND3_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_112 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_112;

architecture SYN_ARCH1 of ND3_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_111 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_111;

architecture SYN_ARCH1 of ND3_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_110 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_110;

architecture SYN_ARCH1 of ND3_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_109 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_109;

architecture SYN_ARCH1 of ND3_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_108 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_108;

architecture SYN_ARCH1 of ND3_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_107 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_107;

architecture SYN_ARCH1 of ND3_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_106 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_106;

architecture SYN_ARCH1 of ND3_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_105 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_105;

architecture SYN_ARCH1 of ND3_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_104 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_104;

architecture SYN_ARCH1 of ND3_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_103 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_103;

architecture SYN_ARCH1 of ND3_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_102 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_102;

architecture SYN_ARCH1 of ND3_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_101 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_101;

architecture SYN_ARCH1 of ND3_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_100 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_100;

architecture SYN_ARCH1 of ND3_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_99 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_99;

architecture SYN_ARCH1 of ND3_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_98 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_98;

architecture SYN_ARCH1 of ND3_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_97 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_97;

architecture SYN_ARCH1 of ND3_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_96 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_96;

architecture SYN_ARCH1 of ND3_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_95 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_95;

architecture SYN_ARCH1 of ND3_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_94 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_94;

architecture SYN_ARCH1 of ND3_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_93 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_93;

architecture SYN_ARCH1 of ND3_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_92 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_92;

architecture SYN_ARCH1 of ND3_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_91 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_91;

architecture SYN_ARCH1 of ND3_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_90 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_90;

architecture SYN_ARCH1 of ND3_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_89 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_89;

architecture SYN_ARCH1 of ND3_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_88 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_88;

architecture SYN_ARCH1 of ND3_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_87 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_87;

architecture SYN_ARCH1 of ND3_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_86 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_86;

architecture SYN_ARCH1 of ND3_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_85 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_85;

architecture SYN_ARCH1 of ND3_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_84 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_84;

architecture SYN_ARCH1 of ND3_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_83 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_83;

architecture SYN_ARCH1 of ND3_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_82 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_82;

architecture SYN_ARCH1 of ND3_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_81 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_81;

architecture SYN_ARCH1 of ND3_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_80 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_80;

architecture SYN_ARCH1 of ND3_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_79 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_79;

architecture SYN_ARCH1 of ND3_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_78 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_78;

architecture SYN_ARCH1 of ND3_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_77 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_77;

architecture SYN_ARCH1 of ND3_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_76 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_76;

architecture SYN_ARCH1 of ND3_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_75 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_75;

architecture SYN_ARCH1 of ND3_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_74 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_74;

architecture SYN_ARCH1 of ND3_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_73 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_73;

architecture SYN_ARCH1 of ND3_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_72 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_72;

architecture SYN_ARCH1 of ND3_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_71 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_71;

architecture SYN_ARCH1 of ND3_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_70 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_70;

architecture SYN_ARCH1 of ND3_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_69 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_69;

architecture SYN_ARCH1 of ND3_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_68 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_68;

architecture SYN_ARCH1 of ND3_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_67 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_67;

architecture SYN_ARCH1 of ND3_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_66 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_66;

architecture SYN_ARCH1 of ND3_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_65 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_65;

architecture SYN_ARCH1 of ND3_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_64 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_64;

architecture SYN_ARCH1 of ND3_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_63 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_63;

architecture SYN_ARCH1 of ND3_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_62 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_62;

architecture SYN_ARCH1 of ND3_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_61 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_61;

architecture SYN_ARCH1 of ND3_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_60 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_60;

architecture SYN_ARCH1 of ND3_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_59 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_59;

architecture SYN_ARCH1 of ND3_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_58 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_58;

architecture SYN_ARCH1 of ND3_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_57 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_57;

architecture SYN_ARCH1 of ND3_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_56 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_56;

architecture SYN_ARCH1 of ND3_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_55 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_55;

architecture SYN_ARCH1 of ND3_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_54 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_54;

architecture SYN_ARCH1 of ND3_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_53 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_53;

architecture SYN_ARCH1 of ND3_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_52 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_52;

architecture SYN_ARCH1 of ND3_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_51 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_51;

architecture SYN_ARCH1 of ND3_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_50 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_50;

architecture SYN_ARCH1 of ND3_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_49 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_49;

architecture SYN_ARCH1 of ND3_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_48 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_48;

architecture SYN_ARCH1 of ND3_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_47 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_47;

architecture SYN_ARCH1 of ND3_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_46 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_46;

architecture SYN_ARCH1 of ND3_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_45 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_45;

architecture SYN_ARCH1 of ND3_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_44 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_44;

architecture SYN_ARCH1 of ND3_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_43 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_43;

architecture SYN_ARCH1 of ND3_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_42 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_42;

architecture SYN_ARCH1 of ND3_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_41 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_41;

architecture SYN_ARCH1 of ND3_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_40 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_40;

architecture SYN_ARCH1 of ND3_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_39 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_39;

architecture SYN_ARCH1 of ND3_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_38 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_38;

architecture SYN_ARCH1 of ND3_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_37 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_37;

architecture SYN_ARCH1 of ND3_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_36 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_36;

architecture SYN_ARCH1 of ND3_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_35 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_35;

architecture SYN_ARCH1 of ND3_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_34 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_34;

architecture SYN_ARCH1 of ND3_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_33 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_33;

architecture SYN_ARCH1 of ND3_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_32 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_32;

architecture SYN_ARCH1 of ND3_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_31 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_31;

architecture SYN_ARCH1 of ND3_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_30 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_30;

architecture SYN_ARCH1 of ND3_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_29 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_29;

architecture SYN_ARCH1 of ND3_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_28 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_28;

architecture SYN_ARCH1 of ND3_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_27 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_27;

architecture SYN_ARCH1 of ND3_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_26 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_26;

architecture SYN_ARCH1 of ND3_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_25 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_25;

architecture SYN_ARCH1 of ND3_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_24 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_24;

architecture SYN_ARCH1 of ND3_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_23 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_23;

architecture SYN_ARCH1 of ND3_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_22 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_22;

architecture SYN_ARCH1 of ND3_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_21 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_21;

architecture SYN_ARCH1 of ND3_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_20 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_20;

architecture SYN_ARCH1 of ND3_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_19 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_19;

architecture SYN_ARCH1 of ND3_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_18 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_18;

architecture SYN_ARCH1 of ND3_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_17 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_17;

architecture SYN_ARCH1 of ND3_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_16 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_16;

architecture SYN_ARCH1 of ND3_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_15 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_15;

architecture SYN_ARCH1 of ND3_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_14 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_14;

architecture SYN_ARCH1 of ND3_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_13 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_13;

architecture SYN_ARCH1 of ND3_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_12 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_12;

architecture SYN_ARCH1 of ND3_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_11 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_11;

architecture SYN_ARCH1 of ND3_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_10 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_10;

architecture SYN_ARCH1 of ND3_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_9 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_9;

architecture SYN_ARCH1 of ND3_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_8 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_8;

architecture SYN_ARCH1 of ND3_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_7 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_7;

architecture SYN_ARCH1 of ND3_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_6 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_6;

architecture SYN_ARCH1 of ND3_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_5 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_5;

architecture SYN_ARCH1 of ND3_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_4 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_4;

architecture SYN_ARCH1 of ND3_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_3 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_3;

architecture SYN_ARCH1 of ND3_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_2 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_2;

architecture SYN_ARCH1 of ND3_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_1 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_1;

architecture SYN_ARCH1 of ND3_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 is

   component CARRY_SEL_N_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_55 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_54 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_53 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_52 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_51 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_50 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_49 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 is

   component CARRY_SEL_N_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_47 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_46 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_45 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_44 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_43 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_42 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_41 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 is

   component CARRY_SEL_N_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_39 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_38 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_37 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_36 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_35 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_34 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_33 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 is

   component CARRY_SEL_N_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_31 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_30 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_29 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_28 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_27 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_26 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_25 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 is

   component CARRY_SEL_N_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_23 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_22 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_21 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_20 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_19 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_18 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_17 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 is

   component CARRY_SEL_N_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_15 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_14 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_13 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_12 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_11 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_10 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_9 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 is

   component CARRY_SEL_N_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_55
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_56
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_57
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_58
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_163
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_164
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_59
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_60
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_165
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_166
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_167
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_61
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_168
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_169
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_170
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_171
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_172
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_173
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_174
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_62
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_175
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_176
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_177
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_178
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_179
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_180
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_181
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_182
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_183
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_184
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_185
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_186
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_187
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_188
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_189
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_63
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n2, n3, n4, n5, n6, n_1132 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n6);
   pgnetwork_0 : PG_network_NBIT32_7 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1132, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_63 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_189 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_188 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_187 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_186 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_185 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_184 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_183 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_182 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_181 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_180 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_179 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_178 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_177 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_176 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_175 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_62 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_174 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_173 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_172 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_171 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_170 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_169 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_168 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_61 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_167 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_166 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_165 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_60 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_59 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_164 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_163 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_58 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_57 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_56 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_55 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Cin, A2 => n6, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => n4, A2 => n5, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_46
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_47
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_48
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_49
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_136
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_137
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_50
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_51
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_138
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_139
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_140
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_52
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_141
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_142
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_143
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_144
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_145
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_146
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_147
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_53
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_148
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_149
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_150
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_151
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_152
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_153
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_154
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_155
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_156
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_157
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_158
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_159
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_160
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_161
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_162
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_54
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, n9,
      n10, G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, G_16_9_port, 
      G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, G_12_12_port, 
      G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, G_10_9_port, 
      G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, G_6_6_port, 
      G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, G_2_2_port, 
      G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, G_32_25_port, 
      G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, G_29_29_port, 
      G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, G_27_27_port, 
      G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, G_24_23_port, 
      G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, G_22_21_port, 
      G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, G_19_19_port, 
      G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, P_32_32_port, P_32_31_port, P_32_29_port, 
      P_32_25_port, P_32_17_port, P_31_31_port, P_30_30_port, P_30_29_port, 
      P_29_29_port, P_28_28_port, P_28_27_port, P_28_25_port, P_28_17_port, 
      P_27_27_port, P_26_26_port, P_26_25_port, P_25_25_port, P_24_24_port, 
      P_24_23_port, P_24_21_port, P_24_17_port, P_23_23_port, P_22_22_port, 
      P_22_21_port, P_21_21_port, P_20_20_port, P_20_19_port, P_20_17_port, 
      P_19_19_port, P_18_18_port, P_18_17_port, P_17_17_port, Co_2_port, 
      Co_1_port, n4, n5, n6, n7, n8, n_1133 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n8);
   pgnetwork_0 : PG_network_NBIT32_6 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1133, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n7);
   gblock1_1_1 : G_block_54 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_162 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_161 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_160 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_159 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_158 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_157 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_156 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_155 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_154 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_153 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_152 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_151 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_150 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_149 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_148 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_53 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => n10);
   pgblock1_2_2 : PG_block_147 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_146 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_145 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_144 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_143 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_142 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_141 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_52 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => n10, Gout => n9);
   pgblock1_3_2 : PG_block_140 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_139 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_138 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_51 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => n9, Gout => Co_3_port);
   gblock2_4_4 : G_block_50 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => n9, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_137 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_136 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_49 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_48 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_47 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_46 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : CLKBUF_X1 port map( A => n9, Z => Co_2_port);
   U2 : CLKBUF_X1 port map( A => n10, Z => Co_1_port);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Cin, A2 => n8, ZN => n4);
   U6 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n5);
   U7 : AND2_X1 port map( A1 => n6, A2 => n7, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_37
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_38
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_39
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_40
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_109
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_110
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_41
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_42
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_111
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_112
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_113
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_43
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_114
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_115
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_116
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_117
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_118
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_119
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_120
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_44
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_121
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_122
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_123
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_124
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_125
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_126
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_127
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_128
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_129
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_130
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_131
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_132
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_133
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_134
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_135
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_45
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n2, n3, n4, n5, n6, n_1134 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n6);
   pgnetwork_0 : PG_network_NBIT32_5 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1134, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_45 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_135 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_134 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_133 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_132 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_131 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_130 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_129 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_128 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_127 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_126 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_125 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_124 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_123 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_122 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_121 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_44 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_120 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_119 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_118 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_117 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_116 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_115 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_114 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_43 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_113 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_112 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_111 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_42 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_41 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_110 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_109 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_40 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_39 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_38 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_37 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Cin, A2 => n6, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => n4, A2 => n5, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_28
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_29
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_30
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_31
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_82
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_83
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_32
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_33
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_84
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_85
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_86
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_34
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_87
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_88
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_89
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_90
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_91
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_92
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_93
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_35
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_94
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_95
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_96
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_97
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_98
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_99
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_100
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_101
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_102
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_103
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_104
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_105
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_106
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_107
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_108
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_36
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, n8,
      n9, G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, G_16_9_port, 
      G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, G_12_12_port, 
      G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, G_10_9_port, 
      G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, G_6_6_port, 
      G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, G_2_2_port, 
      G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, G_32_25_port, 
      G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, G_29_29_port, 
      G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, G_27_27_port, 
      G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, G_24_23_port, 
      G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, G_22_21_port, 
      G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, G_19_19_port, 
      G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, P_32_32_port, P_32_31_port, P_32_29_port, 
      P_32_25_port, P_32_17_port, P_31_31_port, P_30_30_port, P_30_29_port, 
      P_29_29_port, P_28_28_port, P_28_27_port, P_28_25_port, P_28_17_port, 
      P_27_27_port, P_26_26_port, P_26_25_port, P_25_25_port, P_24_24_port, 
      P_24_23_port, P_24_21_port, P_24_17_port, P_23_23_port, P_22_22_port, 
      P_22_21_port, P_21_21_port, P_20_20_port, P_20_19_port, P_20_17_port, 
      P_19_19_port, P_18_18_port, P_18_17_port, P_17_17_port, N1, N2, n2_port, 
      Co_2_port, Co_1_port, n5, n6, n7, n_1135 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n7);
   pgnetwork_0 : PG_network_NBIT32_4 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1135, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n6);
   gblock1_1_1 : G_block_36 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_108 port map( A(1) => P_4_4_port, A(0) => G_4_4_port
                           , B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) 
                           => P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_107 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_106 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_105 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_104 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_103 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_102 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_101 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_100 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_99 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_98 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_97 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_96 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_95 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_94 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_35 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => n9);
   pgblock1_2_2 : PG_block_93 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_92 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_91 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_90 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_89 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_88 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_87 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_34 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => n9, Gout => n8);
   pgblock1_3_2 : PG_block_86 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_85 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_84 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_33 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_32 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => n8, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_83 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_82 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_31 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_30 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_29 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_28 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => n2_port, Gout => Co_8_port);
   U1 : CLKBUF_X1 port map( A => Co_4_port, Z => n2_port);
   U2 : BUF_X2 port map( A => n8, Z => Co_2_port);
   U4 : CLKBUF_X1 port map( A => n9, Z => Co_1_port);
   U5 : OR2_X1 port map( A1 => N1, A2 => N2, ZN => n5);
   U6 : AND2_X1 port map( A1 => Cin, A2 => n7, ZN => N1);
   U7 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => N2);
   U8 : AND2_X1 port map( A1 => n5, A2 => n6, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_block_19
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_20
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_21
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_22
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_55
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_56
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_23
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_24
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_57
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_58
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_59
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_25
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_60
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_61
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_62
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_63
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_64
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_65
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_66
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_26
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_67
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_68
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_69
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_70
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_71
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_72
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_73
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_74
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_75
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_76
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_77
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_78
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_79
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_80
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_81
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_27
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, n8, Co_3_port, Co_2_port,
      Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_16_16_port, 
      P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, 
      P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, 
      P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, 
      P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, 
      P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, Co_4_port, n3, n4, n5, n6, n7, n_1136 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n7);
   pgnetwork_0 : PG_network_NBIT32_3 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1136, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n6);
   gblock1_1_1 : G_block_27 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_81 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_80 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_79 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_78 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_77 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_76 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_75 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_74 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_73 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_72 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_71 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_70 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_69 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_68 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_67 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_26 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_66 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_65 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_64 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_63 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_62 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_61 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_60 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_25 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_59 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_58 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_57 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_24 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_23 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => n8);
   pgblock2_4_28_2 : PG_block_56 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_55 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_22 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => n8, Gout => Co_5_port);
   gblock2_5_6 : G_block_21 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => n8, Gout => Co_6_port);
   gblock2_5_7 : G_block_20 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => n8, Gout => Co_7_port);
   gblock2_5_8 : G_block_19 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : BUF_X1 port map( A => n8, Z => Co_4_port);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Cin, A2 => n7, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n4);
   U6 : AND2_X1 port map( A1 => n5, A2 => n6, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_10
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_11
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_12
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_13
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_28
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_29
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_14
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_15
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_30
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_31
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_32
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_16
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_33
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_34
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_35
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_36
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_37
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_38
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_39
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_17
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_40
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_41
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_42
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_43
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_44
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_45
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_46
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_47
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_48
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_49
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_50
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_51
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_52
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_53
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_54
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_18
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n2, n3, n4, n5, n6, n_1137 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n6);
   pgnetwork_0 : PG_network_NBIT32_2 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1137, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_18 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_54 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_53 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_52 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_51 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_50 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_49 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_48 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_47 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_46 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_45 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_44 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_43 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_42 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_41 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_40 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_17 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_39 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_38 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_37 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_36 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_35 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_34 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_33 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_16 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_32 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_31 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_30 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_15 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_14 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_29 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_28 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_13 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_12 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_11 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_10 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Cin, A2 => n6, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => n4, A2 => n5, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_1
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_2
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_3
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_4
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_1
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_2
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_5
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_6
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_3
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_4
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_5
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_7
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_6
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_7
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_8
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_9
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_10
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_11
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_12
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_8
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_13
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_14
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_15
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_16
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_17
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_18
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_19
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_20
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_21
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_22
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_23
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_24
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_25
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_26
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_27
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_9
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n2, n3, n4, n5, n6, n_1138 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => n6);
   pgnetwork_0 : PG_network_NBIT32_1 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1138, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_9 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B 
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_27 port map( A(1) => P_4_4_port, A(0) => G_4_4_port,
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_26 port map( A(1) => P_6_6_port, A(0) => G_6_6_port,
                           B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) => 
                           P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_25 port map( A(1) => P_8_8_port, A(0) => G_8_8_port,
                           B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) => 
                           P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_24 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_23 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_22 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_21 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_20 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_19 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_18 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_17 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_16 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_15 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_14 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_13 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_8 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B 
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_12 port map( A(1) => P_8_7_port, A(0) => G_8_7_port,
                           B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) => 
                           P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_11 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_10 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_9 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_8 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_7 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_6 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_7 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B 
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_5 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_4 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_3 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_6 port map( A(1) => P_12_9_port, A(0) => G_12_9_port, 
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_5 port map( A(1) => P_16_9_port, A(0) => G_16_9_port, 
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_2 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_1 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_4 port map( A(1) => P_20_17_port, A(0) => G_20_17_port
                           , B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_3 port map( A(1) => P_24_17_port, A(0) => G_24_17_port
                           , B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_2 port map( A(1) => P_28_17_port, A(0) => G_28_17_port
                           , B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_1 port map( A(1) => P_32_17_port, A(0) => G_32_17_port
                           , B => Co_4_port, Gout => Co_8_port);
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Cin, A2 => n6, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n3);
   U5 : AND2_X1 port map( A1 => n4, A2 => n5, ZN => G_1_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_7 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_7;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_7 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_7 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_6 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_6;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_6 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2 : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_6 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_6 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : INV_X1 port map( A => ADD_SUB, ZN => n1);
   U11 : INV_X1 port map( A => ADD_SUB, ZN => n2);
   U36 : XNOR2_X2 port map( A => B(3), B => n1, ZN => B_in_3_port);
   U37 : XNOR2_X2 port map( A => B(0), B => n2, ZN => B_in_0_port);
   U38 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_5 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_5;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_5 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3 : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_5 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_5 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => n1, A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : INV_X1 port map( A => ADD_SUB, ZN => n3);
   U21 : INV_X1 port map( A => ADD_SUB, ZN => n2);
   U23 : CLKBUF_X1 port map( A => A(22), Z => n1);
   U37 : XNOR2_X1 port map( A => B(21), B => n2, ZN => B_in_21_port);
   U38 : XNOR2_X1 port map( A => B(23), B => n3, ZN => B_in_23_port);
   U39 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_4 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_4;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1 : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_4 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_4 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : INV_X1 port map( A => ADD_SUB, ZN => n1);
   U36 : XNOR2_X2 port map( A => B(0), B => n1, ZN => B_in_0_port);
   U37 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2, n3 : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_3 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => n3, A(22) => A(22), A(21) => n1, 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : INV_X1 port map( A => ADD_SUB, ZN => n2);
   U21 : CLKBUF_X1 port map( A => A(21), Z => n1);
   U37 : XNOR2_X1 port map( A => B(23), B => n2, ZN => B_in_23_port);
   U38 : CLKBUF_X1 port map( A => A(23), Z => n3);
   U39 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_2 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U11 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U36 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, 
      B_in_12_port, B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, 
      B_in_7_port, B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, 
      B_in_2_port, B_in_1_port, B_in_0_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_in_16_port);
   U30 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_in_15_port);
   U31 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_in_14_port);
   U32 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_in_13_port);
   U33 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_in_10_port);
   U36 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_in_0_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => 
                           B_in_15_port, B(14) => B_in_14_port, B(13) => 
                           B_in_13_port, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => B_in_0_port, Cin => C_internal,
                           Co(8) => Cout, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_1 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : OR2_X1 port map( A1 => ADD_SUB, A2 => Cin, ZN => C_internal);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_228;

architecture SYN_Behavioral of AND2_228 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_227;

architecture SYN_Behavioral of AND2_227 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_226;

architecture SYN_Behavioral of AND2_226 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_225;

architecture SYN_Behavioral of AND2_225 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_224;

architecture SYN_Behavioral of AND2_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_223;

architecture SYN_Behavioral of AND2_223 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_222;

architecture SYN_Behavioral of AND2_222 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_221;

architecture SYN_Behavioral of AND2_221 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_220;

architecture SYN_Behavioral of AND2_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_219;

architecture SYN_Behavioral of AND2_219 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_218;

architecture SYN_Behavioral of AND2_218 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_217;

architecture SYN_Behavioral of AND2_217 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_216;

architecture SYN_Behavioral of AND2_216 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_215;

architecture SYN_Behavioral of AND2_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_214;

architecture SYN_Behavioral of AND2_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_213;

architecture SYN_Behavioral of AND2_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_212;

architecture SYN_Behavioral of AND2_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_211;

architecture SYN_Behavioral of AND2_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_210;

architecture SYN_Behavioral of AND2_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_209;

architecture SYN_Behavioral of AND2_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_208;

architecture SYN_Behavioral of AND2_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_207;

architecture SYN_Behavioral of AND2_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_206;

architecture SYN_Behavioral of AND2_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_205;

architecture SYN_Behavioral of AND2_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_204;

architecture SYN_Behavioral of AND2_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_203;

architecture SYN_Behavioral of AND2_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_202;

architecture SYN_Behavioral of AND2_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_201;

architecture SYN_Behavioral of AND2_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_200;

architecture SYN_Behavioral of AND2_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_199;

architecture SYN_Behavioral of AND2_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_198;

architecture SYN_Behavioral of AND2_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_197;

architecture SYN_Behavioral of AND2_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_196;

architecture SYN_Behavioral of AND2_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_195;

architecture SYN_Behavioral of AND2_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_194;

architecture SYN_Behavioral of AND2_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_193;

architecture SYN_Behavioral of AND2_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_192;

architecture SYN_Behavioral of AND2_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_191;

architecture SYN_Behavioral of AND2_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_190;

architecture SYN_Behavioral of AND2_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_189;

architecture SYN_Behavioral of AND2_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_188;

architecture SYN_Behavioral of AND2_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_187;

architecture SYN_Behavioral of AND2_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_186;

architecture SYN_Behavioral of AND2_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_185;

architecture SYN_Behavioral of AND2_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_184;

architecture SYN_Behavioral of AND2_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_183;

architecture SYN_Behavioral of AND2_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_182;

architecture SYN_Behavioral of AND2_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_181;

architecture SYN_Behavioral of AND2_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_180;

architecture SYN_Behavioral of AND2_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_179;

architecture SYN_Behavioral of AND2_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_178;

architecture SYN_Behavioral of AND2_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_177;

architecture SYN_Behavioral of AND2_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_176;

architecture SYN_Behavioral of AND2_176 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_175;

architecture SYN_Behavioral of AND2_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_174;

architecture SYN_Behavioral of AND2_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_173;

architecture SYN_Behavioral of AND2_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_172;

architecture SYN_Behavioral of AND2_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_171;

architecture SYN_Behavioral of AND2_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_170;

architecture SYN_Behavioral of AND2_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_169;

architecture SYN_Behavioral of AND2_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_168;

architecture SYN_Behavioral of AND2_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_167;

architecture SYN_Behavioral of AND2_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_166;

architecture SYN_Behavioral of AND2_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_165;

architecture SYN_Behavioral of AND2_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_164;

architecture SYN_Behavioral of AND2_164 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_163;

architecture SYN_Behavioral of AND2_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_162;

architecture SYN_Behavioral of AND2_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_161;

architecture SYN_Behavioral of AND2_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_160;

architecture SYN_Behavioral of AND2_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_159;

architecture SYN_Behavioral of AND2_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_158;

architecture SYN_Behavioral of AND2_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_157;

architecture SYN_Behavioral of AND2_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_156;

architecture SYN_Behavioral of AND2_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_155;

architecture SYN_Behavioral of AND2_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_154;

architecture SYN_Behavioral of AND2_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_153;

architecture SYN_Behavioral of AND2_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_152;

architecture SYN_Behavioral of AND2_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_151;

architecture SYN_Behavioral of AND2_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_150;

architecture SYN_Behavioral of AND2_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_149;

architecture SYN_Behavioral of AND2_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_148;

architecture SYN_Behavioral of AND2_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_147;

architecture SYN_Behavioral of AND2_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_146;

architecture SYN_Behavioral of AND2_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_145;

architecture SYN_Behavioral of AND2_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_144;

architecture SYN_Behavioral of AND2_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_143;

architecture SYN_Behavioral of AND2_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_142;

architecture SYN_Behavioral of AND2_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_141;

architecture SYN_Behavioral of AND2_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_140;

architecture SYN_Behavioral of AND2_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_139;

architecture SYN_Behavioral of AND2_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_138;

architecture SYN_Behavioral of AND2_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_137;

architecture SYN_Behavioral of AND2_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_136;

architecture SYN_Behavioral of AND2_136 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_135;

architecture SYN_Behavioral of AND2_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_134;

architecture SYN_Behavioral of AND2_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_133;

architecture SYN_Behavioral of AND2_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_132;

architecture SYN_Behavioral of AND2_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_131;

architecture SYN_Behavioral of AND2_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_130;

architecture SYN_Behavioral of AND2_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_129;

architecture SYN_Behavioral of AND2_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_128;

architecture SYN_Behavioral of AND2_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_127;

architecture SYN_Behavioral of AND2_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_126;

architecture SYN_Behavioral of AND2_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_125;

architecture SYN_Behavioral of AND2_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_124;

architecture SYN_Behavioral of AND2_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_123;

architecture SYN_Behavioral of AND2_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_122;

architecture SYN_Behavioral of AND2_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_121;

architecture SYN_Behavioral of AND2_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_120;

architecture SYN_Behavioral of AND2_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_119;

architecture SYN_Behavioral of AND2_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_118;

architecture SYN_Behavioral of AND2_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_117;

architecture SYN_Behavioral of AND2_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_116;

architecture SYN_Behavioral of AND2_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_115;

architecture SYN_Behavioral of AND2_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_114;

architecture SYN_Behavioral of AND2_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_113;

architecture SYN_Behavioral of AND2_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_112;

architecture SYN_Behavioral of AND2_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_111;

architecture SYN_Behavioral of AND2_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_110;

architecture SYN_Behavioral of AND2_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_109;

architecture SYN_Behavioral of AND2_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_108;

architecture SYN_Behavioral of AND2_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_107;

architecture SYN_Behavioral of AND2_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_106;

architecture SYN_Behavioral of AND2_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_105;

architecture SYN_Behavioral of AND2_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_104;

architecture SYN_Behavioral of AND2_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_103;

architecture SYN_Behavioral of AND2_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_102;

architecture SYN_Behavioral of AND2_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_101;

architecture SYN_Behavioral of AND2_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_100;

architecture SYN_Behavioral of AND2_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_99;

architecture SYN_Behavioral of AND2_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_98;

architecture SYN_Behavioral of AND2_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_97;

architecture SYN_Behavioral of AND2_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_96;

architecture SYN_Behavioral of AND2_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_95;

architecture SYN_Behavioral of AND2_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_94;

architecture SYN_Behavioral of AND2_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_93;

architecture SYN_Behavioral of AND2_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_92;

architecture SYN_Behavioral of AND2_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_91;

architecture SYN_Behavioral of AND2_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_90;

architecture SYN_Behavioral of AND2_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_89;

architecture SYN_Behavioral of AND2_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_88;

architecture SYN_Behavioral of AND2_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_87;

architecture SYN_Behavioral of AND2_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_86;

architecture SYN_Behavioral of AND2_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_85;

architecture SYN_Behavioral of AND2_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_84;

architecture SYN_Behavioral of AND2_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_83;

architecture SYN_Behavioral of AND2_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_82;

architecture SYN_Behavioral of AND2_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_81;

architecture SYN_Behavioral of AND2_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_80;

architecture SYN_Behavioral of AND2_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_79;

architecture SYN_Behavioral of AND2_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_78;

architecture SYN_Behavioral of AND2_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_77;

architecture SYN_Behavioral of AND2_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_76;

architecture SYN_Behavioral of AND2_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_75;

architecture SYN_Behavioral of AND2_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_74;

architecture SYN_Behavioral of AND2_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_73;

architecture SYN_Behavioral of AND2_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_72;

architecture SYN_Behavioral of AND2_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_71;

architecture SYN_Behavioral of AND2_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_70;

architecture SYN_Behavioral of AND2_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_69;

architecture SYN_Behavioral of AND2_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_68;

architecture SYN_Behavioral of AND2_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_67;

architecture SYN_Behavioral of AND2_67 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_66;

architecture SYN_Behavioral of AND2_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_65;

architecture SYN_Behavioral of AND2_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_64;

architecture SYN_Behavioral of AND2_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_63;

architecture SYN_Behavioral of AND2_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_62;

architecture SYN_Behavioral of AND2_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_61;

architecture SYN_Behavioral of AND2_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_60;

architecture SYN_Behavioral of AND2_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_59;

architecture SYN_Behavioral of AND2_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_58;

architecture SYN_Behavioral of AND2_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_57;

architecture SYN_Behavioral of AND2_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_56;

architecture SYN_Behavioral of AND2_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_55;

architecture SYN_Behavioral of AND2_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_54;

architecture SYN_Behavioral of AND2_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_53;

architecture SYN_Behavioral of AND2_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_52;

architecture SYN_Behavioral of AND2_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_51;

architecture SYN_Behavioral of AND2_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_50;

architecture SYN_Behavioral of AND2_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_49;

architecture SYN_Behavioral of AND2_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_48;

architecture SYN_Behavioral of AND2_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_47;

architecture SYN_Behavioral of AND2_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_46;

architecture SYN_Behavioral of AND2_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_45;

architecture SYN_Behavioral of AND2_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_44;

architecture SYN_Behavioral of AND2_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_43;

architecture SYN_Behavioral of AND2_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_42;

architecture SYN_Behavioral of AND2_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_41;

architecture SYN_Behavioral of AND2_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_40;

architecture SYN_Behavioral of AND2_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_39;

architecture SYN_Behavioral of AND2_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_38;

architecture SYN_Behavioral of AND2_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_37;

architecture SYN_Behavioral of AND2_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_36;

architecture SYN_Behavioral of AND2_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_35;

architecture SYN_Behavioral of AND2_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_34;

architecture SYN_Behavioral of AND2_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_33;

architecture SYN_Behavioral of AND2_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_32;

architecture SYN_Behavioral of AND2_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_31;

architecture SYN_Behavioral of AND2_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_30;

architecture SYN_Behavioral of AND2_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_29;

architecture SYN_Behavioral of AND2_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_28;

architecture SYN_Behavioral of AND2_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_27;

architecture SYN_Behavioral of AND2_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_26;

architecture SYN_Behavioral of AND2_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_25;

architecture SYN_Behavioral of AND2_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_24;

architecture SYN_Behavioral of AND2_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_23;

architecture SYN_Behavioral of AND2_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_22;

architecture SYN_Behavioral of AND2_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_21;

architecture SYN_Behavioral of AND2_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_20;

architecture SYN_Behavioral of AND2_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_19;

architecture SYN_Behavioral of AND2_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_18;

architecture SYN_Behavioral of AND2_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_17;

architecture SYN_Behavioral of AND2_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_16;

architecture SYN_Behavioral of AND2_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_15;

architecture SYN_Behavioral of AND2_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_14;

architecture SYN_Behavioral of AND2_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_13;

architecture SYN_Behavioral of AND2_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_12;

architecture SYN_Behavioral of AND2_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_11;

architecture SYN_Behavioral of AND2_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_10;

architecture SYN_Behavioral of AND2_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_9;

architecture SYN_Behavioral of AND2_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_8;

architecture SYN_Behavioral of AND2_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_7;

architecture SYN_Behavioral of AND2_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_6;

architecture SYN_Behavioral of AND2_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_5;

architecture SYN_Behavioral of AND2_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_4;

architecture SYN_Behavioral of AND2_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_3;

architecture SYN_Behavioral of AND2_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_2;

architecture SYN_Behavioral of AND2_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_1;

architecture SYN_Behavioral of AND2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX4to1_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX4to1_NBIT32_1;

architecture SYN_Behavioral of MUX4to1_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n5, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n147, Z => n72);
   U2 : BUF_X1 port map( A => n148, Z => n76);
   U3 : AND2_X1 port map( A1 => SEL(1), A2 => n84, ZN => n1);
   U4 : BUF_X1 port map( A => n149, Z => n80);
   U5 : BUF_X1 port map( A => n76, Z => n73);
   U6 : BUF_X1 port map( A => n76, Z => n74);
   U7 : BUF_X1 port map( A => n76, Z => n75);
   U8 : BUF_X1 port map( A => n1, Z => n77);
   U9 : BUF_X1 port map( A => n1, Z => n78);
   U10 : BUF_X1 port map( A => n1, Z => n79);
   U11 : BUF_X1 port map( A => n80, Z => n81);
   U12 : BUF_X1 port map( A => n80, Z => n82);
   U13 : BUF_X1 port map( A => n80, Z => n83);
   U14 : BUF_X1 port map( A => n72, Z => n5);
   U15 : BUF_X1 port map( A => n72, Z => n70);
   U16 : BUF_X1 port map( A => n72, Z => n71);
   U17 : AOI22_X1 port map( A1 => D(21), A2 => n82, B1 => C(21), B2 => n78, ZN 
                           => n111);
   U18 : AOI22_X1 port map( A1 => D(22), A2 => n82, B1 => C(22), B2 => n78, ZN 
                           => n113);
   U19 : AOI22_X1 port map( A1 => D(25), A2 => n82, B1 => C(25), B2 => n78, ZN 
                           => n119);
   U20 : AOI22_X1 port map( A1 => D(20), A2 => n82, B1 => C(20), B2 => n78, ZN 
                           => n109);
   U21 : AOI22_X1 port map( A1 => D(27), A2 => n82, B1 => C(27), B2 => n78, ZN 
                           => n123);
   U22 : AOI22_X1 port map( A1 => B(18), A2 => n73, B1 => A(18), B2 => n5, ZN 
                           => n104);
   U23 : AOI22_X1 port map( A1 => B(4), A2 => n75, B1 => A(4), B2 => n71, ZN =>
                           n138);
   U24 : AOI22_X1 port map( A1 => B(6), A2 => n75, B1 => A(6), B2 => n71, ZN =>
                           n142);
   U25 : AOI22_X1 port map( A1 => B(3), A2 => n75, B1 => A(3), B2 => n71, ZN =>
                           n136);
   U26 : AOI22_X1 port map( A1 => B(12), A2 => n73, B1 => A(12), B2 => n5, ZN 
                           => n92);
   U27 : AOI22_X1 port map( A1 => B(17), A2 => n73, B1 => A(17), B2 => n5, ZN 
                           => n102);
   U28 : AOI22_X1 port map( A1 => B(15), A2 => n73, B1 => A(15), B2 => n5, ZN 
                           => n98);
   U29 : AOI22_X1 port map( A1 => B(1), A2 => n73, B1 => A(1), B2 => n5, ZN => 
                           n108);
   U30 : AOI22_X1 port map( A1 => B(14), A2 => n73, B1 => A(14), B2 => n5, ZN 
                           => n96);
   U31 : AOI22_X1 port map( A1 => B(7), A2 => n75, B1 => A(7), B2 => n71, ZN =>
                           n144);
   U32 : AOI22_X1 port map( A1 => B(5), A2 => n75, B1 => A(5), B2 => n71, ZN =>
                           n140);
   U33 : AOI22_X1 port map( A1 => B(16), A2 => n73, B1 => A(16), B2 => n5, ZN 
                           => n100);
   U34 : AOI22_X1 port map( A1 => B(2), A2 => n74, B1 => A(2), B2 => n70, ZN =>
                           n130);
   U35 : AOI22_X1 port map( A1 => B(0), A2 => n73, B1 => A(0), B2 => n5, ZN => 
                           n86);
   U36 : AOI22_X1 port map( A1 => B(10), A2 => n73, B1 => A(10), B2 => n5, ZN 
                           => n88);
   U37 : AOI22_X1 port map( A1 => B(19), A2 => n73, B1 => A(19), B2 => n5, ZN 
                           => n106);
   U38 : AOI22_X1 port map( A1 => B(13), A2 => n73, B1 => A(13), B2 => n5, ZN 
                           => n94);
   U39 : AOI22_X1 port map( A1 => B(8), A2 => n75, B1 => A(8), B2 => n71, ZN =>
                           n146);
   U40 : AOI22_X1 port map( A1 => B(9), A2 => n75, B1 => A(9), B2 => n71, ZN =>
                           n151);
   U41 : AOI22_X1 port map( A1 => D(11), A2 => n81, B1 => C(11), B2 => n77, ZN 
                           => n89);
   U42 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => Y(20));
   U43 : AOI22_X1 port map( A1 => B(20), A2 => n74, B1 => A(20), B2 => n70, ZN 
                           => n110);
   U44 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => B(21), A2 => n74, B1 => A(21), B2 => n70, ZN 
                           => n112);
   U46 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => Y(22));
   U47 : AOI22_X1 port map( A1 => B(22), A2 => n74, B1 => A(22), B2 => n70, ZN 
                           => n114);
   U48 : AOI22_X1 port map( A1 => B(25), A2 => n74, B1 => A(25), B2 => n70, ZN 
                           => n120);
   U49 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => Y(28));
   U50 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => Y(24));
   U51 : AOI22_X1 port map( A1 => B(24), A2 => n74, B1 => A(24), B2 => n70, ZN 
                           => n118);
   U52 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => Y(26));
   U53 : AOI22_X1 port map( A1 => B(26), A2 => n74, B1 => A(26), B2 => n70, ZN 
                           => n122);
   U54 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => Y(31));
   U55 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n71, ZN 
                           => n134);
   U56 : AOI22_X1 port map( A1 => B(30), A2 => n74, B1 => A(30), B2 => n70, ZN 
                           => n132);
   U57 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => Y(29));
   U58 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => Y(18));
   U59 : AOI22_X1 port map( A1 => D(18), A2 => n81, B1 => C(18), B2 => n77, ZN 
                           => n103);
   U60 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => Y(3));
   U61 : AOI22_X1 port map( A1 => D(3), A2 => n83, B1 => C(3), B2 => n79, ZN =>
                           n135);
   U62 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => Y(4));
   U63 : AOI22_X1 port map( A1 => D(4), A2 => n83, B1 => C(4), B2 => n79, ZN =>
                           n137);
   U64 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => Y(6));
   U65 : AOI22_X1 port map( A1 => D(6), A2 => n83, B1 => C(6), B2 => n79, ZN =>
                           n141);
   U66 : AOI22_X1 port map( A1 => D(15), A2 => n81, B1 => C(15), B2 => n77, ZN 
                           => n97);
   U67 : AOI22_X1 port map( A1 => D(17), A2 => n81, B1 => C(17), B2 => n77, ZN 
                           => n101);
   U68 : AOI22_X1 port map( A1 => D(1), A2 => n81, B1 => C(1), B2 => n77, ZN =>
                           n107);
   U69 : AOI22_X1 port map( A1 => D(14), A2 => n81, B1 => C(14), B2 => n77, ZN 
                           => n95);
   U70 : AOI22_X1 port map( A1 => D(7), A2 => n83, B1 => C(7), B2 => n79, ZN =>
                           n143);
   U71 : AOI22_X1 port map( A1 => D(5), A2 => n83, B1 => C(5), B2 => n79, ZN =>
                           n139);
   U72 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => Y(0));
   U73 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Y(10));
   U74 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Y(13));
   U75 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => Y(19));
   U76 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Y(9));
   U77 : AOI22_X1 port map( A1 => B(28), A2 => n74, B1 => A(28), B2 => n70, ZN 
                           => n126);
   U78 : AOI22_X1 port map( A1 => B(23), A2 => n74, B1 => A(23), B2 => n70, ZN 
                           => n116);
   U79 : AOI22_X1 port map( A1 => B(29), A2 => n74, B1 => A(29), B2 => n70, ZN 
                           => n128);
   U80 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => Y(17));
   U81 : AND2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n149);
   U82 : INV_X1 port map( A => SEL(0), ZN => n84);
   U83 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n147);
   U84 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => Y(14));
   U85 : AOI22_X1 port map( A1 => D(16), A2 => n81, B1 => C(16), B2 => n77, ZN 
                           => n99);
   U86 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => Y(16));
   U87 : AOI22_X1 port map( A1 => D(30), A2 => n82, B1 => C(30), B2 => n78, ZN 
                           => n131);
   U88 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Y(12));
   U89 : AOI22_X1 port map( A1 => D(12), A2 => n81, B1 => C(12), B2 => n77, ZN 
                           => n91);
   U90 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => Y(30));
   U91 : AOI22_X1 port map( A1 => D(29), A2 => n82, B1 => C(29), B2 => n78, ZN 
                           => n127);
   U92 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => Y(5));
   U93 : AOI22_X1 port map( A1 => D(26), A2 => n82, B1 => C(26), B2 => n78, ZN 
                           => n121);
   U94 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Y(11));
   U95 : AOI22_X1 port map( A1 => B(11), A2 => n73, B1 => A(11), B2 => n5, ZN 
                           => n90);
   U96 : NOR2_X1 port map( A1 => n84, A2 => SEL(1), ZN => n148);
   U97 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => Y(25));
   U98 : AOI22_X1 port map( A1 => B(27), A2 => n74, B1 => A(27), B2 => n70, ZN 
                           => n124);
   U99 : AOI22_X1 port map( A1 => D(31), A2 => n83, B1 => C(31), B2 => n79, ZN 
                           => n133);
   U100 : AOI22_X1 port map( A1 => D(24), A2 => n82, B1 => C(24), B2 => n78, ZN
                           => n117);
   U101 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => Y(23));
   U102 : AOI22_X1 port map( A1 => D(23), A2 => n82, B1 => C(23), B2 => n78, ZN
                           => n115);
   U103 : AOI22_X1 port map( A1 => D(10), A2 => n81, B1 => C(10), B2 => n77, ZN
                           => n87);
   U104 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => Y(2));
   U105 : AOI22_X1 port map( A1 => D(2), A2 => n82, B1 => C(2), B2 => n78, ZN 
                           => n129);
   U106 : AOI22_X1 port map( A1 => D(19), A2 => n81, B1 => C(19), B2 => n77, ZN
                           => n105);
   U107 : AOI22_X1 port map( A1 => D(13), A2 => n81, B1 => C(13), B2 => n77, ZN
                           => n93);
   U108 : AOI22_X1 port map( A1 => D(9), A2 => n83, B1 => C(9), B2 => n79, ZN 
                           => n150);
   U109 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Y(15));
   U110 : AOI22_X1 port map( A1 => D(28), A2 => n82, B1 => C(28), B2 => n78, ZN
                           => n125);
   U111 : NAND2_X1 port map( A1 => n144, A2 => n143, ZN => Y(7));
   U112 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => Y(27));
   U113 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => Y(1));
   U114 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => Y(8));
   U115 : AOI22_X1 port map( A1 => D(8), A2 => n83, B1 => C(8), B2 => n79, ZN 
                           => n145);
   U116 : AOI22_X1 port map( A1 => D(0), A2 => n81, B1 => C(0), B2 => n77, ZN 
                           => n85);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_8 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_8;

architecture SYN_Behavioral of MUX5to1_NBIT32_8 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n166, Z => n90);
   U6 : BUF_X1 port map( A => n163, Z => n78);
   U7 : BUF_X1 port map( A => n162, Z => n74);
   U8 : BUF_X1 port map( A => n165, Z => n83);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : INV_X1 port map( A => SEL(1), ZN => n97);
   U17 : INV_X1 port map( A => SEL(0), ZN => n98);
   U18 : BUF_X1 port map( A => n90, Z => n87);
   U19 : BUF_X1 port map( A => n90, Z => n88);
   U20 : BUF_X1 port map( A => n78, Z => n76);
   U21 : BUF_X1 port map( A => n78, Z => n75);
   U22 : BUF_X1 port map( A => n74, Z => n2);
   U23 : BUF_X1 port map( A => n74, Z => n1);
   U24 : BUF_X1 port map( A => n83, Z => n85);
   U25 : BUF_X1 port map( A => n83, Z => n84);
   U26 : BUF_X1 port map( A => n82, Z => n79);
   U27 : BUF_X1 port map( A => n82, Z => n80);
   U28 : BUF_X1 port map( A => n83, Z => n86);
   U29 : BUF_X1 port map( A => n82, Z => n81);
   U30 : BUF_X1 port map( A => n78, Z => n77);
   U31 : BUF_X1 port map( A => n74, Z => n73);
   U32 : BUF_X1 port map( A => n90, Z => n89);
   U33 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U36 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U37 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U38 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U39 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN =>
                           n103);
   U40 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U41 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U42 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN =>
                           n105);
   U43 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U44 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U45 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN =>
                           n107);
   U46 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U47 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U48 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN =>
                           n109);
   U49 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U50 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U51 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n111);
   U52 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U53 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U54 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n113);
   U55 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U56 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U57 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n115);
   U58 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U59 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U60 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n117);
   U61 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U62 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U63 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n119);
   U64 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U65 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U66 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U67 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n79, ZN => n120);
   U68 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U69 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U70 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n122);
   U71 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U72 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U73 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U74 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U75 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U76 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U77 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U78 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U79 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U80 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U81 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U82 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U83 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U84 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U85 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U86 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U87 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U88 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U89 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U90 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U91 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U92 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U93 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U94 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U95 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U96 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U97 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U98 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U99 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U100 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, 
                           C1 => D(21), C2 => n80, ZN => n142);
   U101 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U102 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U103 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, 
                           C1 => D(22), C2 => n80, ZN => n144);
   U104 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U105 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U106 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, 
                           C1 => D(23), C2 => n81, ZN => n146);
   U107 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U108 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U109 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, 
                           C1 => D(24), C2 => n81, ZN => n148);
   U110 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U111 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U112 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n81, ZN => n150);
   U113 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U114 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U115 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n81, ZN => n152);
   U116 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U117 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U118 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n81, ZN => n154);
   U119 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U120 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U121 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n81, ZN => n156);
   U122 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U123 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U124 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n81, ZN => n158);
   U125 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U126 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U127 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n81, ZN => n160);
   U128 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U129 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U130 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n167);
   U131 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U132 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n101);
   U133 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_7 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_7;

architecture SYN_Behavioral of MUX5to1_NBIT32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U39 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN =>
                           n107);
   U40 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U41 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U42 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN =>
                           n109);
   U43 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U44 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U45 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n111);
   U46 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U47 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U48 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n113);
   U49 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U50 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U51 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n115);
   U52 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U53 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U54 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n117);
   U55 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U56 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U57 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n119);
   U58 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U59 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U60 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U61 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n79, ZN => n120);
   U62 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U63 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U64 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n122);
   U65 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U66 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U67 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U68 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U69 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U70 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U71 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U72 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U73 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U74 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U75 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U76 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U77 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U78 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U79 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U80 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U81 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U82 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U83 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U84 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U85 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U86 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U87 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U88 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U89 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U90 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U91 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U92 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U93 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U94 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U95 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U96 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U97 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U98 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U99 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U100 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, 
                           C1 => D(23), C2 => n81, ZN => n146);
   U101 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U102 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U103 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, 
                           C1 => D(24), C2 => n81, ZN => n148);
   U104 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U105 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U106 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n81, ZN => n150);
   U107 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U108 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U109 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n81, ZN => n152);
   U110 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U111 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U112 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n81, ZN => n154);
   U113 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U114 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U115 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n81, ZN => n156);
   U116 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U117 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U118 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n81, ZN => n158);
   U119 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U120 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U121 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n81, ZN => n160);
   U122 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U123 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U124 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n167);
   U125 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U126 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n105);
   U127 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U128 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U129 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n101);
   U130 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U131 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U132 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n103);
   U133 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_6 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_6;

architecture SYN_Behavioral of MUX5to1_NBIT32_6 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U39 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U40 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U41 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U42 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n111);
   U43 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U44 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U45 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n113);
   U46 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U47 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U48 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n115);
   U49 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U50 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U51 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n117);
   U52 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U53 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U54 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n119);
   U55 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U56 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U57 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U58 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n79, ZN => n120);
   U59 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U60 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U61 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n122);
   U62 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U63 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U64 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U65 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U66 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U67 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U68 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U69 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U70 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U71 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U72 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U73 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U74 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U75 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U76 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U77 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U78 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U79 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U80 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U81 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U82 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U83 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U84 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U85 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U86 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U87 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U88 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U89 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U90 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U91 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U92 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U93 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U94 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n81, ZN => n146);
   U95 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U96 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U97 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n81, ZN => n148);
   U98 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U99 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U100 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n81, ZN => n150);
   U101 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U102 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U103 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n81, ZN => n152);
   U104 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U105 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U106 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n81, ZN => n154);
   U107 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U108 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U109 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n81, ZN => n156);
   U110 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U111 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U112 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n81, ZN => n158);
   U113 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U114 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U115 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n81, ZN => n160);
   U116 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U117 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U118 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n167);
   U119 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U120 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n109);
   U121 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U122 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U123 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n101);
   U124 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U125 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U126 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n103);
   U127 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U128 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U129 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n105);
   U130 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U131 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U132 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n107);
   U133 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_5 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_5;

architecture SYN_Behavioral of MUX5to1_NBIT32_5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U39 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n115);
   U40 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U41 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U42 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n117);
   U43 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U44 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U45 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n119);
   U46 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U47 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U48 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U49 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n79, ZN => n120);
   U50 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U51 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U52 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n122);
   U53 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U54 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U55 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U56 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U57 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U58 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U59 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U60 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U61 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U62 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U63 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U64 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U65 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U66 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U67 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U68 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U69 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U70 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U71 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U72 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U73 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U74 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U75 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U76 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U77 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U78 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U79 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U80 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U81 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U82 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U83 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U84 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U85 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U86 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U87 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U88 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n81, ZN => n146);
   U89 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U90 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U91 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n81, ZN => n148);
   U92 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U93 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U94 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n81, ZN => n150);
   U95 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U96 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U97 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n81, ZN => n152);
   U98 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U99 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U100 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n81, ZN => n154);
   U101 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U102 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U103 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n81, ZN => n156);
   U104 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U105 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U106 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n81, ZN => n158);
   U107 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U108 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U109 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n81, ZN => n160);
   U110 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U111 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U112 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n167);
   U113 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U114 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n113);
   U115 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U116 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U117 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n101);
   U118 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U119 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U120 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n103);
   U121 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U122 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U123 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n105);
   U124 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U125 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U126 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n107);
   U127 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U128 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U129 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n109);
   U130 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U131 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U132 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n111);
   U133 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_4 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_4;

architecture SYN_Behavioral of MUX5to1_NBIT32_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U39 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n119);
   U40 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U41 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U42 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U43 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n79, ZN => n120);
   U44 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U45 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U46 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n122);
   U47 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U48 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U49 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U50 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U51 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U52 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U53 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U54 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U55 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U56 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U57 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U58 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U59 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U60 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U61 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U62 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U63 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U64 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U65 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U66 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U67 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U68 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U69 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U70 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U71 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U72 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U73 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U74 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U75 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U76 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U77 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U78 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U79 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U80 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U81 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U82 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n81, ZN => n146);
   U83 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U84 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U85 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n81, ZN => n148);
   U86 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U87 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U88 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n81, ZN => n150);
   U89 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U90 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U91 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n81, ZN => n152);
   U92 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U93 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U94 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n81, ZN => n154);
   U95 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U96 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U97 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n81, ZN => n156);
   U98 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U99 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U100 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n81, ZN => n158);
   U101 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U102 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U103 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n81, ZN => n160);
   U104 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U105 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U106 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n167);
   U107 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U108 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n117);
   U109 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U110 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U111 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n101);
   U112 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U113 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U114 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n103);
   U115 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U116 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U117 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n105);
   U118 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U119 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U120 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n107);
   U121 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U122 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U123 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n109);
   U124 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U125 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U126 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n111);
   U127 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U128 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U129 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n113);
   U130 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U131 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U132 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n115);
   U133 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_3 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_3;

architecture SYN_Behavioral of MUX5to1_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U39 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U40 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n122);
   U41 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U42 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U43 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U44 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U45 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U46 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U47 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U48 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U49 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U50 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U51 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U52 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U53 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U54 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U55 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U56 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U57 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U58 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U59 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U60 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U61 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U62 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U63 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U64 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U65 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U66 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U67 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U68 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U69 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U70 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U71 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U72 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U73 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U74 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U75 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U76 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n81, ZN => n146);
   U77 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U78 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U79 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n81, ZN => n148);
   U80 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U81 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U82 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n81, ZN => n150);
   U83 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U84 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U85 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n81, ZN => n152);
   U86 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U87 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U88 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n81, ZN => n154);
   U89 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U90 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U91 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n81, ZN => n156);
   U92 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U93 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U94 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n81, ZN => n158);
   U95 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U96 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U97 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, C1
                           => D(30), C2 => n81, ZN => n160);
   U98 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U99 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U100 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n167);
   U101 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U102 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U103 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, 
                           C1 => D(10), C2 => n79, ZN => n120);
   U104 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U105 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN 
                           => n101);
   U106 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U107 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U108 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n103);
   U109 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U110 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U111 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n105);
   U112 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U113 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U114 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n107);
   U115 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U116 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U117 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n109);
   U118 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U119 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U120 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n111);
   U121 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U122 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U123 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n113);
   U124 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U125 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U126 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n115);
   U127 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U128 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U129 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n117);
   U130 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U131 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U132 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN =>
                           n119);
   U133 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_2 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_2;

architecture SYN_Behavioral of MUX5to1_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U39 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U40 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n126);
   U41 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U42 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U43 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U44 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U45 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U46 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U47 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U48 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U49 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U50 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U51 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U52 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U53 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U54 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U55 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U56 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U57 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U58 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U59 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U60 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U61 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U62 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U63 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U64 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U65 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U66 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U67 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U68 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U69 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U70 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n81, ZN => n146);
   U71 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U72 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U73 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n81, ZN => n148);
   U74 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U75 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U76 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n81, ZN => n150);
   U77 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U78 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U79 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n81, ZN => n152);
   U80 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U81 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U82 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n81, ZN => n154);
   U83 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U84 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U85 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n81, ZN => n156);
   U86 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U87 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U88 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n81, ZN => n158);
   U89 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U90 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U91 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, C1
                           => D(30), C2 => n81, ZN => n160);
   U92 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U93 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U94 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, C1
                           => D(31), C2 => n81, ZN => n167);
   U95 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U96 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U97 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n124);
   U98 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U99 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN =>
                           n101);
   U100 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U101 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U102 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN 
                           => n103);
   U103 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U104 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U105 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN 
                           => n105);
   U106 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U107 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U108 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n107);
   U109 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U110 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U111 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n109);
   U112 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U113 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U114 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n111);
   U115 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U116 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U117 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n113);
   U118 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U119 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U120 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n115);
   U121 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U122 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U123 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n117);
   U124 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U125 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U126 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN =>
                           n119);
   U127 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U128 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U129 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U130 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, 
                           C1 => D(10), C2 => n79, ZN => n120);
   U131 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U132 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U133 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, 
                           C1 => D(11), C2 => n80, ZN => n122);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_1 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_1;

architecture SYN_Behavioral of MUX5to1_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n1, n2, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n164, Z => n82);
   U5 : BUF_X1 port map( A => n163, Z => n78);
   U6 : BUF_X1 port map( A => n165, Z => n83);
   U7 : BUF_X1 port map( A => n166, Z => n90);
   U8 : BUF_X1 port map( A => n162, Z => n74);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n99, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n99);
   U16 : BUF_X1 port map( A => n78, Z => n76);
   U17 : BUF_X1 port map( A => n78, Z => n75);
   U18 : BUF_X1 port map( A => n83, Z => n85);
   U19 : BUF_X1 port map( A => n83, Z => n84);
   U20 : BUF_X1 port map( A => n82, Z => n79);
   U21 : BUF_X1 port map( A => n82, Z => n80);
   U22 : BUF_X1 port map( A => n83, Z => n86);
   U23 : BUF_X1 port map( A => n82, Z => n81);
   U24 : BUF_X1 port map( A => n78, Z => n77);
   U25 : INV_X1 port map( A => SEL(1), ZN => n97);
   U26 : NOR3_X1 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n164);
   U27 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n163);
   U28 : AND3_X1 port map( A1 => n98, A2 => n97, A3 => SEL(2), ZN => n165);
   U29 : BUF_X1 port map( A => n90, Z => n87);
   U30 : BUF_X1 port map( A => n90, Z => n88);
   U31 : BUF_X1 port map( A => n74, Z => n2);
   U32 : BUF_X1 port map( A => n74, Z => n1);
   U33 : BUF_X1 port map( A => n74, Z => n73);
   U34 : BUF_X1 port map( A => n90, Z => n89);
   U35 : INV_X1 port map( A => SEL(0), ZN => n98);
   U36 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n166);
   U37 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n162
                           );
   U38 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => N41);
   U39 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n131);
   U40 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n130);
   U41 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => N42);
   U42 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n133);
   U43 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n132);
   U44 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => N43);
   U45 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n135);
   U46 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n134);
   U47 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => N44);
   U48 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n137);
   U49 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n136);
   U50 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => N45);
   U51 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n139);
   U52 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n138);
   U53 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => N46);
   U54 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n141);
   U55 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, C1
                           => D(20), C2 => n80, ZN => n140);
   U56 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => N47);
   U57 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n143);
   U58 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, C1
                           => D(21), C2 => n80, ZN => n142);
   U59 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => N48);
   U60 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n145);
   U61 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, C1
                           => D(22), C2 => n80, ZN => n144);
   U62 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => N49);
   U63 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n147);
   U64 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, C1
                           => D(23), C2 => n81, ZN => n146);
   U65 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => N50);
   U66 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n149);
   U67 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, C1
                           => D(24), C2 => n81, ZN => n148);
   U68 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => N51);
   U69 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n151);
   U70 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, C1
                           => D(25), C2 => n81, ZN => n150);
   U71 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => N52);
   U72 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n153);
   U73 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, C1
                           => D(26), C2 => n81, ZN => n152);
   U74 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => N53);
   U75 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n155);
   U76 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, C1
                           => D(27), C2 => n81, ZN => n154);
   U77 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => N54);
   U78 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n157);
   U79 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, C1
                           => D(28), C2 => n81, ZN => n156);
   U80 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => N55);
   U81 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n159);
   U82 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, C1
                           => D(29), C2 => n81, ZN => n158);
   U83 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => N56);
   U84 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n161);
   U85 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, C1
                           => D(30), C2 => n81, ZN => n160);
   U86 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => N57);
   U87 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n168);
   U88 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, C1
                           => D(31), C2 => n81, ZN => n167);
   U89 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => N40);
   U90 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n129);
   U91 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n128);
   U92 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => N26);
   U93 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN =>
                           n101);
   U94 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n100);
   U95 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => N27);
   U96 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN =>
                           n103);
   U97 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n102);
   U98 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => N28);
   U99 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN =>
                           n105);
   U100 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n104);
   U101 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => N29);
   U102 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN 
                           => n107);
   U103 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n106);
   U104 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => N30);
   U105 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN 
                           => n109);
   U106 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n108);
   U107 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => N31);
   U108 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN 
                           => n111);
   U109 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n110);
   U110 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => N32);
   U111 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN 
                           => n113);
   U112 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n112);
   U113 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => N33);
   U114 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN 
                           => n115);
   U115 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n114);
   U116 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => N34);
   U117 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN =>
                           n117);
   U118 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n116);
   U119 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => N35);
   U120 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN =>
                           n119);
   U121 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n118);
   U122 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => N36);
   U123 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n121);
   U124 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, 
                           C1 => D(10), C2 => n79, ZN => n120);
   U125 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => N37);
   U126 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n123);
   U127 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, 
                           C1 => D(11), C2 => n80, ZN => n122);
   U128 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => N38);
   U129 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n125);
   U130 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, 
                           C1 => D(12), C2 => n80, ZN => n124);
   U131 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => N39);
   U132 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n127);
   U133 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, 
                           C1 => D(13), C2 => n80, ZN => n126);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_8 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_8;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n80, ZN => Y(1));
   U2 : BUF_X1 port map( A => n68, Z => n1);
   U3 : BUF_X1 port map( A => n68, Z => n2);
   U4 : BUF_X1 port map( A => n68, Z => n3);
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => SEL, ZN => 
                           n80);
   U6 : INV_X1 port map( A => n91, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => SEL, ZN => 
                           n91);
   U8 : INV_X1 port map( A => n94, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => SEL, ZN => 
                           n94);
   U10 : INV_X1 port map( A => n95, ZN => Y(4));
   U11 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => SEL, ZN => 
                           n95);
   U12 : INV_X1 port map( A => n96, ZN => Y(5));
   U13 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => SEL, ZN => 
                           n96);
   U14 : INV_X1 port map( A => n97, ZN => Y(6));
   U15 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => SEL, ZN => 
                           n97);
   U16 : INV_X1 port map( A => n98, ZN => Y(7));
   U17 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => SEL, ZN => 
                           n98);
   U18 : INV_X1 port map( A => n99, ZN => Y(8));
   U19 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => SEL, ZN => 
                           n99);
   U20 : INV_X1 port map( A => n100, ZN => Y(9));
   U21 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => SEL, B2 => B(9), ZN => 
                           n100);
   U22 : INV_X1 port map( A => n70, ZN => Y(10));
   U23 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => SEL, ZN 
                           => n70);
   U24 : INV_X1 port map( A => n71, ZN => Y(11));
   U25 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => SEL, ZN 
                           => n71);
   U26 : INV_X1 port map( A => n72, ZN => Y(12));
   U27 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => SEL, ZN 
                           => n72);
   U28 : INV_X1 port map( A => n73, ZN => Y(13));
   U29 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => SEL, ZN 
                           => n73);
   U30 : INV_X1 port map( A => n74, ZN => Y(14));
   U31 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => SEL, ZN 
                           => n74);
   U32 : INV_X1 port map( A => n75, ZN => Y(15));
   U33 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => SEL, ZN 
                           => n75);
   U34 : INV_X1 port map( A => n76, ZN => Y(16));
   U35 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => SEL, ZN 
                           => n76);
   U36 : INV_X1 port map( A => n77, ZN => Y(17));
   U37 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => SEL, ZN 
                           => n77);
   U38 : INV_X1 port map( A => n78, ZN => Y(18));
   U39 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => SEL, ZN 
                           => n78);
   U40 : INV_X1 port map( A => n79, ZN => Y(19));
   U41 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => SEL, ZN 
                           => n79);
   U42 : INV_X1 port map( A => n81, ZN => Y(20));
   U43 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => SEL, ZN 
                           => n81);
   U44 : INV_X1 port map( A => n82, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => SEL, ZN 
                           => n82);
   U46 : INV_X1 port map( A => n83, ZN => Y(22));
   U47 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => SEL, ZN 
                           => n83);
   U48 : INV_X1 port map( A => n84, ZN => Y(23));
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => SEL, ZN 
                           => n84);
   U50 : INV_X1 port map( A => n85, ZN => Y(24));
   U51 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => SEL, ZN 
                           => n85);
   U52 : INV_X1 port map( A => n86, ZN => Y(25));
   U53 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => SEL, ZN 
                           => n86);
   U54 : INV_X1 port map( A => n87, ZN => Y(26));
   U55 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => SEL, ZN 
                           => n87);
   U56 : INV_X1 port map( A => n88, ZN => Y(27));
   U57 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => SEL, ZN 
                           => n88);
   U58 : INV_X1 port map( A => n89, ZN => Y(28));
   U59 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => SEL, ZN 
                           => n89);
   U60 : INV_X1 port map( A => n90, ZN => Y(29));
   U61 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => SEL, ZN 
                           => n90);
   U62 : INV_X1 port map( A => n92, ZN => Y(30));
   U63 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => SEL, ZN 
                           => n92);
   U64 : INV_X1 port map( A => n69, ZN => Y(0));
   U65 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => SEL, ZN => 
                           n69);
   U66 : INV_X1 port map( A => SEL, ZN => n68);
   U67 : INV_X1 port map( A => n93, ZN => Y(31));
   U68 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => SEL, ZN 
                           => n93);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_7;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net46339, net46337, net46335, net46331, n1, n32, n33, n54, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88 : std_logic;

begin
   
   U1 : INV_X2 port map( A => net46335, ZN => net46331);
   U2 : INV_X1 port map( A => n79, ZN => Y(2));
   U3 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U4 : CLKBUF_X1 port map( A => net46339, Z => net46337);
   U5 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U6 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U7 : CLKBUF_X1 port map( A => net46339, Z => net46335);
   U8 : INV_X1 port map( A => n1, ZN => net46339);
   U9 : INV_X1 port map( A => n68, ZN => Y(19));
   U10 : INV_X1 port map( A => n67, ZN => Y(18));
   U11 : INV_X1 port map( A => n66, ZN => Y(17));
   U12 : INV_X1 port map( A => n65, ZN => Y(16));
   U13 : INV_X1 port map( A => n64, ZN => Y(15));
   U14 : INV_X1 port map( A => n63, ZN => Y(14));
   U15 : INV_X1 port map( A => n62, ZN => Y(13));
   U16 : INV_X1 port map( A => n54, ZN => Y(12));
   U17 : INV_X1 port map( A => n33, ZN => Y(11));
   U18 : INV_X1 port map( A => n32, ZN => Y(10));
   U19 : INV_X1 port map( A => n88, ZN => Y(9));
   U20 : INV_X1 port map( A => n87, ZN => Y(8));
   U21 : INV_X1 port map( A => n86, ZN => Y(7));
   U22 : INV_X1 port map( A => n85, ZN => Y(6));
   U23 : INV_X1 port map( A => n84, ZN => Y(5));
   U24 : INV_X1 port map( A => n83, ZN => Y(4));
   U25 : INV_X1 port map( A => n82, ZN => Y(3));
   U26 : INV_X1 port map( A => n81, ZN => Y(31));
   U27 : INV_X1 port map( A => n80, ZN => Y(30));
   U28 : INV_X1 port map( A => n78, ZN => Y(29));
   U29 : INV_X1 port map( A => n77, ZN => Y(28));
   U30 : INV_X1 port map( A => n76, ZN => Y(27));
   U31 : INV_X1 port map( A => n75, ZN => Y(26));
   U32 : INV_X1 port map( A => n74, ZN => Y(25));
   U33 : INV_X1 port map( A => n73, ZN => Y(24));
   U34 : INV_X1 port map( A => n72, ZN => Y(23));
   U35 : INV_X1 port map( A => n71, ZN => Y(22));
   U36 : INV_X1 port map( A => n70, ZN => Y(21));
   U37 : INV_X1 port map( A => n69, ZN => Y(20));
   U38 : AOI22_X1 port map( A1 => A(2), A2 => net46339, B1 => B(2), B2 => n1, 
                           ZN => n79);
   U39 : AOI22_X1 port map( A1 => A(19), A2 => net46335, B1 => B(19), B2 => 
                           net46331, ZN => n68);
   U40 : AOI22_X1 port map( A1 => A(18), A2 => net46335, B1 => B(18), B2 => 
                           net46331, ZN => n67);
   U41 : AOI22_X1 port map( A1 => A(17), A2 => net46335, B1 => B(17), B2 => 
                           net46331, ZN => n66);
   U42 : AOI22_X1 port map( A1 => A(16), A2 => net46335, B1 => B(16), B2 => 
                           net46331, ZN => n65);
   U43 : AOI22_X1 port map( A1 => A(15), A2 => net46335, B1 => B(15), B2 => 
                           net46331, ZN => n64);
   U44 : AOI22_X1 port map( A1 => A(14), A2 => net46335, B1 => B(14), B2 => 
                           net46331, ZN => n63);
   U45 : AOI22_X1 port map( A1 => A(13), A2 => net46335, B1 => B(13), B2 => 
                           net46331, ZN => n62);
   U46 : AOI22_X1 port map( A1 => A(12), A2 => net46335, B1 => B(12), B2 => 
                           net46331, ZN => n54);
   U47 : AOI22_X1 port map( A1 => A(11), A2 => net46335, B1 => B(11), B2 => 
                           net46331, ZN => n33);
   U48 : AOI22_X1 port map( A1 => A(10), A2 => net46335, B1 => B(10), B2 => 
                           net46331, ZN => n32);
   U49 : AOI22_X1 port map( A1 => A(9), A2 => net46337, B1 => net46331, B2 => 
                           B(9), ZN => n88);
   U50 : AOI22_X1 port map( A1 => A(8), A2 => net46337, B1 => B(8), B2 => 
                           net46331, ZN => n87);
   U51 : AOI22_X1 port map( A1 => A(7), A2 => net46337, B1 => B(7), B2 => 
                           net46331, ZN => n86);
   U52 : AOI22_X1 port map( A1 => A(6), A2 => net46337, B1 => B(6), B2 => 
                           net46331, ZN => n85);
   U53 : AOI22_X1 port map( A1 => A(5), A2 => net46337, B1 => B(5), B2 => 
                           net46331, ZN => n84);
   U54 : AOI22_X1 port map( A1 => A(4), A2 => net46337, B1 => B(4), B2 => 
                           net46331, ZN => n83);
   U55 : AOI22_X1 port map( A1 => A(3), A2 => net46337, B1 => B(3), B2 => 
                           net46331, ZN => n82);
   U56 : AOI22_X1 port map( A1 => A(31), A2 => net46337, B1 => B(31), B2 => 
                           net46331, ZN => n81);
   U57 : AOI22_X1 port map( A1 => A(30), A2 => net46335, B1 => B(30), B2 => 
                           net46331, ZN => n80);
   U58 : AOI22_X1 port map( A1 => A(29), A2 => net46335, B1 => B(29), B2 => 
                           net46331, ZN => n78);
   U59 : AOI22_X1 port map( A1 => A(28), A2 => net46335, B1 => B(28), B2 => 
                           net46331, ZN => n77);
   U60 : AOI22_X1 port map( A1 => A(27), A2 => net46335, B1 => B(27), B2 => 
                           net46331, ZN => n76);
   U61 : AOI22_X1 port map( A1 => A(26), A2 => net46335, B1 => B(26), B2 => 
                           net46331, ZN => n75);
   U62 : AOI22_X1 port map( A1 => A(25), A2 => net46335, B1 => B(25), B2 => 
                           net46331, ZN => n74);
   U63 : AOI22_X1 port map( A1 => A(24), A2 => net46335, B1 => B(24), B2 => 
                           net46331, ZN => n73);
   U64 : AOI22_X1 port map( A1 => A(23), A2 => net46335, B1 => B(23), B2 => 
                           net46331, ZN => n72);
   U65 : AOI22_X1 port map( A1 => A(22), A2 => net46335, B1 => B(22), B2 => 
                           net46331, ZN => n71);
   U66 : AOI22_X1 port map( A1 => A(21), A2 => net46335, B1 => B(21), B2 => 
                           net46331, ZN => n70);
   U67 : AOI22_X1 port map( A1 => A(20), A2 => net46335, B1 => B(20), B2 => 
                           net46331, ZN => n69);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_6;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n9, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : INV_X1 port map( A => n8, ZN => n6);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n5, Z => n8);
   U7 : INV_X1 port map( A => n85, ZN => Y(1));
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n6, B1 => B(1), B2 => n1, ZN => 
                           n85);
   U9 : INV_X1 port map( A => n96, ZN => Y(2));
   U10 : AOI22_X1 port map( A1 => A(2), A2 => n7, B1 => B(2), B2 => n2, ZN => 
                           n96);
   U11 : INV_X1 port map( A => n99, ZN => Y(3));
   U12 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => n3, ZN => 
                           n99);
   U13 : INV_X1 port map( A => n100, ZN => Y(4));
   U14 : AOI22_X1 port map( A1 => A(4), A2 => n7, B1 => B(4), B2 => n3, ZN => 
                           n100);
   U15 : INV_X1 port map( A => n101, ZN => Y(5));
   U16 : AOI22_X1 port map( A1 => A(5), A2 => n6, B1 => B(5), B2 => n3, ZN => 
                           n101);
   U17 : INV_X1 port map( A => n102, ZN => Y(6));
   U18 : AOI22_X1 port map( A1 => A(6), A2 => n7, B1 => B(6), B2 => n3, ZN => 
                           n102);
   U19 : INV_X1 port map( A => n103, ZN => Y(7));
   U20 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n3, ZN => 
                           n103);
   U21 : INV_X1 port map( A => n104, ZN => Y(8));
   U22 : AOI22_X1 port map( A1 => A(8), A2 => n7, B1 => B(8), B2 => n3, ZN => 
                           n104);
   U23 : INV_X1 port map( A => n105, ZN => Y(9));
   U24 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n3, B2 => B(9), ZN => 
                           n105);
   U25 : INV_X1 port map( A => n75, ZN => Y(10));
   U26 : AOI22_X1 port map( A1 => A(10), A2 => n6, B1 => B(10), B2 => n1, ZN =>
                           n75);
   U27 : INV_X1 port map( A => n77, ZN => Y(12));
   U28 : AOI22_X1 port map( A1 => A(12), A2 => n6, B1 => B(12), B2 => n1, ZN =>
                           n77);
   U29 : INV_X1 port map( A => n78, ZN => Y(13));
   U30 : AOI22_X1 port map( A1 => A(13), A2 => n6, B1 => B(13), B2 => n1, ZN =>
                           n78);
   U31 : INV_X1 port map( A => n79, ZN => Y(14));
   U32 : AOI22_X1 port map( A1 => A(14), A2 => n6, B1 => B(14), B2 => n1, ZN =>
                           n79);
   U33 : INV_X1 port map( A => n80, ZN => Y(15));
   U34 : AOI22_X1 port map( A1 => A(15), A2 => n6, B1 => B(15), B2 => n1, ZN =>
                           n80);
   U35 : INV_X1 port map( A => n76, ZN => Y(11));
   U36 : AOI22_X1 port map( A1 => A(11), A2 => n6, B1 => B(11), B2 => n1, ZN =>
                           n76);
   U37 : INV_X1 port map( A => n93, ZN => Y(27));
   U38 : AOI22_X1 port map( A1 => A(27), A2 => n7, B1 => B(27), B2 => n2, ZN =>
                           n93);
   U39 : INV_X1 port map( A => n86, ZN => Y(20));
   U40 : AOI22_X1 port map( A1 => A(20), A2 => n7, B1 => B(20), B2 => n1, ZN =>
                           n86);
   U41 : INV_X1 port map( A => n90, ZN => Y(24));
   U42 : AOI22_X1 port map( A1 => A(24), A2 => n7, B1 => B(24), B2 => n2, ZN =>
                           n90);
   U43 : INV_X1 port map( A => n81, ZN => Y(16));
   U44 : AOI22_X1 port map( A1 => A(16), A2 => n6, B1 => B(16), B2 => n1, ZN =>
                           n81);
   U45 : INV_X1 port map( A => n82, ZN => Y(17));
   U46 : AOI22_X1 port map( A1 => A(17), A2 => n6, B1 => B(17), B2 => n1, ZN =>
                           n82);
   U47 : INV_X1 port map( A => n83, ZN => Y(18));
   U48 : AOI22_X1 port map( A1 => A(18), A2 => n6, B1 => B(18), B2 => n1, ZN =>
                           n83);
   U49 : INV_X1 port map( A => n84, ZN => Y(19));
   U50 : AOI22_X1 port map( A1 => A(19), A2 => n6, B1 => B(19), B2 => n1, ZN =>
                           n84);
   U51 : INV_X1 port map( A => n87, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n7, B1 => B(21), B2 => n2, ZN =>
                           n87);
   U53 : INV_X1 port map( A => n88, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n7, B1 => B(22), B2 => n2, ZN =>
                           n88);
   U55 : INV_X1 port map( A => n89, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n7, B1 => B(23), B2 => n2, ZN =>
                           n89);
   U57 : INV_X1 port map( A => n91, ZN => Y(25));
   U58 : AOI22_X1 port map( A1 => A(25), A2 => n7, B1 => B(25), B2 => n2, ZN =>
                           n91);
   U59 : INV_X1 port map( A => n92, ZN => Y(26));
   U60 : AOI22_X1 port map( A1 => A(26), A2 => n7, B1 => B(26), B2 => n2, ZN =>
                           n92);
   U61 : INV_X1 port map( A => n94, ZN => Y(28));
   U62 : AOI22_X1 port map( A1 => A(28), A2 => n7, B1 => B(28), B2 => n2, ZN =>
                           n94);
   U63 : INV_X1 port map( A => n95, ZN => Y(29));
   U64 : AOI22_X1 port map( A1 => A(29), A2 => n7, B1 => B(29), B2 => n2, ZN =>
                           n95);
   U65 : INV_X1 port map( A => n97, ZN => Y(30));
   U66 : AOI22_X1 port map( A1 => A(30), A2 => n7, B1 => B(30), B2 => n2, ZN =>
                           n97);
   U67 : INV_X1 port map( A => n98, ZN => Y(31));
   U68 : AOI22_X1 port map( A1 => A(31), A2 => n7, B1 => B(31), B2 => n2, ZN =>
                           n98);
   U69 : BUF_X1 port map( A => SEL, Z => n5);
   U70 : INV_X1 port map( A => n8, ZN => n7);
   U71 : CLKBUF_X1 port map( A => n5, Z => n9);
   U72 : AOI22_X1 port map( A1 => A(0), A2 => n6, B1 => B(0), B2 => n3, ZN => 
                           n74);
   U73 : INV_X1 port map( A => n74, ZN => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_5;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => n6);
   U2 : BUF_X1 port map( A => n8, Z => n2);
   U3 : BUF_X1 port map( A => n8, Z => n1);
   U4 : INV_X1 port map( A => n7, ZN => n5);
   U5 : BUF_X1 port map( A => n8, Z => n3);
   U6 : BUF_X1 port map( A => n4, Z => n7);
   U7 : BUF_X1 port map( A => n4, Z => n8);
   U8 : INV_X1 port map( A => n73, ZN => Y(0));
   U9 : INV_X1 port map( A => n84, ZN => Y(1));
   U10 : INV_X1 port map( A => n99, ZN => Y(4));
   U11 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U12 : INV_X1 port map( A => n98, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U14 : INV_X1 port map( A => n101, ZN => Y(6));
   U15 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U16 : INV_X1 port map( A => n76, ZN => Y(12));
   U17 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U18 : INV_X1 port map( A => n100, ZN => Y(5));
   U19 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U20 : INV_X1 port map( A => n102, ZN => Y(7));
   U21 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U22 : INV_X1 port map( A => n103, ZN => Y(8));
   U23 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U24 : INV_X1 port map( A => n75, ZN => Y(11));
   U25 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U26 : INV_X1 port map( A => n79, ZN => Y(15));
   U27 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U28 : INV_X1 port map( A => n77, ZN => Y(13));
   U29 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U30 : INV_X1 port map( A => n78, ZN => Y(14));
   U31 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U32 : INV_X1 port map( A => n74, ZN => Y(10));
   U33 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U34 : INV_X1 port map( A => n104, ZN => Y(9));
   U35 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U36 : INV_X1 port map( A => n85, ZN => Y(20));
   U37 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n1, ZN =>
                           n85);
   U38 : INV_X1 port map( A => n97, ZN => Y(31));
   U39 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n2, ZN =>
                           n97);
   U40 : INV_X1 port map( A => n80, ZN => Y(16));
   U41 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U42 : INV_X1 port map( A => n81, ZN => Y(17));
   U43 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U44 : INV_X1 port map( A => n89, ZN => Y(24));
   U45 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U46 : INV_X1 port map( A => n82, ZN => Y(18));
   U47 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U48 : INV_X1 port map( A => n83, ZN => Y(19));
   U49 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U50 : INV_X1 port map( A => n90, ZN => Y(25));
   U51 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U52 : INV_X1 port map( A => n91, ZN => Y(26));
   U53 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U54 : INV_X1 port map( A => n86, ZN => Y(21));
   U55 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U56 : INV_X1 port map( A => n93, ZN => Y(28));
   U57 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U58 : INV_X1 port map( A => n92, ZN => Y(27));
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U60 : INV_X1 port map( A => n87, ZN => Y(22));
   U61 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U62 : INV_X1 port map( A => n88, ZN => Y(23));
   U63 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U64 : INV_X1 port map( A => n94, ZN => Y(29));
   U65 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U66 : INV_X1 port map( A => n96, ZN => Y(30));
   U67 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U68 : BUF_X1 port map( A => SEL, Z => n4);
   U69 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U70 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U71 : INV_X1 port map( A => n95, ZN => Y(2));
   U72 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n3, ZN => 
                           n73);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_4;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n7);
   U2 : BUF_X1 port map( A => n4, Z => n8);
   U3 : BUF_X1 port map( A => n8, Z => n1);
   U4 : BUF_X1 port map( A => n8, Z => n2);
   U5 : INV_X1 port map( A => n7, ZN => n5);
   U6 : INV_X1 port map( A => n7, ZN => n6);
   U7 : BUF_X1 port map( A => n8, Z => n3);
   U8 : BUF_X1 port map( A => SEL, Z => n4);
   U9 : INV_X1 port map( A => n73, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n73);
   U11 : INV_X1 port map( A => n84, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U13 : INV_X1 port map( A => n95, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U15 : INV_X1 port map( A => n98, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U17 : INV_X1 port map( A => n99, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U19 : INV_X1 port map( A => n100, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U21 : INV_X1 port map( A => n101, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U23 : INV_X1 port map( A => n102, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U25 : INV_X1 port map( A => n103, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U27 : INV_X1 port map( A => n104, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U29 : INV_X1 port map( A => n74, ZN => Y(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U31 : INV_X1 port map( A => n75, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U33 : INV_X1 port map( A => n76, ZN => Y(12));
   U34 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U35 : INV_X1 port map( A => n77, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U37 : INV_X1 port map( A => n78, ZN => Y(14));
   U38 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U39 : INV_X1 port map( A => n79, ZN => Y(15));
   U40 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U41 : INV_X1 port map( A => n80, ZN => Y(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U43 : INV_X1 port map( A => n81, ZN => Y(17));
   U44 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U45 : INV_X1 port map( A => n82, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U47 : INV_X1 port map( A => n83, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U49 : INV_X1 port map( A => n85, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U51 : INV_X1 port map( A => n86, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U53 : INV_X1 port map( A => n87, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U55 : INV_X1 port map( A => n88, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U57 : INV_X1 port map( A => n89, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U59 : INV_X1 port map( A => n90, ZN => Y(25));
   U60 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U61 : INV_X1 port map( A => n91, ZN => Y(26));
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U63 : INV_X1 port map( A => n92, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U65 : INV_X1 port map( A => n93, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U67 : INV_X1 port map( A => n94, ZN => Y(29));
   U68 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U69 : INV_X1 port map( A => n96, ZN => Y(30));
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U71 : INV_X1 port map( A => n97, ZN => Y(31));
   U72 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n3, ZN =>
                           n97);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_3;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n8);
   U2 : BUF_X1 port map( A => n4, Z => n7);
   U3 : INV_X1 port map( A => n7, ZN => n5);
   U4 : INV_X1 port map( A => n7, ZN => n6);
   U5 : BUF_X1 port map( A => n8, Z => n1);
   U6 : BUF_X1 port map( A => n8, Z => n2);
   U7 : BUF_X1 port map( A => n8, Z => n3);
   U8 : INV_X1 port map( A => n102, ZN => Y(7));
   U9 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U10 : INV_X1 port map( A => n74, ZN => Y(10));
   U11 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U12 : INV_X1 port map( A => n75, ZN => Y(11));
   U13 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U14 : INV_X1 port map( A => n76, ZN => Y(12));
   U15 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U16 : INV_X1 port map( A => n77, ZN => Y(13));
   U17 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U18 : INV_X1 port map( A => n78, ZN => Y(14));
   U19 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U20 : INV_X1 port map( A => n79, ZN => Y(15));
   U21 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U22 : INV_X1 port map( A => n80, ZN => Y(16));
   U23 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U24 : INV_X1 port map( A => n81, ZN => Y(17));
   U25 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U26 : INV_X1 port map( A => n82, ZN => Y(18));
   U27 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U28 : INV_X1 port map( A => n83, ZN => Y(19));
   U29 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U30 : INV_X1 port map( A => n85, ZN => Y(20));
   U31 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U32 : INV_X1 port map( A => n86, ZN => Y(21));
   U33 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U34 : INV_X1 port map( A => n87, ZN => Y(22));
   U35 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U36 : INV_X1 port map( A => n88, ZN => Y(23));
   U37 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U38 : INV_X1 port map( A => n89, ZN => Y(24));
   U39 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U40 : INV_X1 port map( A => n90, ZN => Y(25));
   U41 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U42 : INV_X1 port map( A => n91, ZN => Y(26));
   U43 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U44 : INV_X1 port map( A => n92, ZN => Y(27));
   U45 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U46 : INV_X1 port map( A => n93, ZN => Y(28));
   U47 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U48 : INV_X1 port map( A => n94, ZN => Y(29));
   U49 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U50 : INV_X1 port map( A => n96, ZN => Y(30));
   U51 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U52 : INV_X1 port map( A => n97, ZN => Y(31));
   U53 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n3, ZN =>
                           n97);
   U54 : INV_X1 port map( A => n104, ZN => Y(9));
   U55 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U56 : INV_X1 port map( A => n84, ZN => Y(1));
   U57 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U58 : INV_X1 port map( A => n95, ZN => Y(2));
   U59 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U60 : INV_X1 port map( A => n98, ZN => Y(3));
   U61 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U62 : INV_X1 port map( A => n99, ZN => Y(4));
   U63 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U64 : INV_X1 port map( A => n100, ZN => Y(5));
   U65 : AOI22_X1 port map( A1 => A(5), A2 => n6, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U66 : INV_X1 port map( A => n101, ZN => Y(6));
   U67 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U68 : INV_X1 port map( A => n103, ZN => Y(8));
   U69 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U70 : INV_X1 port map( A => n73, ZN => Y(0));
   U71 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n73);
   U72 : BUF_X1 port map( A => SEL, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_2;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n7);
   U2 : BUF_X1 port map( A => n4, Z => n8);
   U3 : BUF_X1 port map( A => n8, Z => n1);
   U4 : BUF_X1 port map( A => n8, Z => n2);
   U5 : INV_X1 port map( A => n7, ZN => n5);
   U6 : INV_X1 port map( A => n7, ZN => n6);
   U7 : BUF_X1 port map( A => n8, Z => n3);
   U8 : BUF_X1 port map( A => SEL, Z => n4);
   U9 : INV_X1 port map( A => n73, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => n1, ZN => 
                           n73);
   U11 : INV_X1 port map( A => n84, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U13 : INV_X1 port map( A => n95, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U15 : INV_X1 port map( A => n98, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U17 : INV_X1 port map( A => n99, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U19 : INV_X1 port map( A => n100, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U21 : INV_X1 port map( A => n101, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U23 : INV_X1 port map( A => n102, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U25 : INV_X1 port map( A => n103, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U27 : INV_X1 port map( A => n104, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U29 : INV_X1 port map( A => n74, ZN => Y(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U31 : INV_X1 port map( A => n75, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U33 : INV_X1 port map( A => n76, ZN => Y(12));
   U34 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U35 : INV_X1 port map( A => n77, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n5, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U37 : INV_X1 port map( A => n78, ZN => Y(14));
   U38 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U39 : INV_X1 port map( A => n79, ZN => Y(15));
   U40 : AOI22_X1 port map( A1 => A(15), A2 => n5, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U41 : INV_X1 port map( A => n80, ZN => Y(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U43 : INV_X1 port map( A => n81, ZN => Y(17));
   U44 : AOI22_X1 port map( A1 => A(17), A2 => n5, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U45 : INV_X1 port map( A => n82, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U47 : INV_X1 port map( A => n83, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n5, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U49 : INV_X1 port map( A => n85, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n6, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U51 : INV_X1 port map( A => n86, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => n6, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U53 : INV_X1 port map( A => n87, ZN => Y(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n6, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U55 : INV_X1 port map( A => n88, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => A(23), A2 => n6, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U57 : INV_X1 port map( A => n89, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A(24), A2 => n6, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U59 : INV_X1 port map( A => n90, ZN => Y(25));
   U60 : AOI22_X1 port map( A1 => A(25), A2 => n6, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U61 : INV_X1 port map( A => n91, ZN => Y(26));
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n6, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U63 : INV_X1 port map( A => n92, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n6, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U65 : INV_X1 port map( A => n93, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n6, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U67 : INV_X1 port map( A => n94, ZN => Y(29));
   U68 : AOI22_X1 port map( A1 => A(29), A2 => n6, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U69 : INV_X1 port map( A => n96, ZN => Y(30));
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U71 : INV_X1 port map( A => n97, ZN => Y(31));
   U72 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n3, ZN =>
                           n97);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_1;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n4, Z => n8);
   U2 : BUF_X1 port map( A => n4, Z => n7);
   U3 : BUF_X1 port map( A => SEL, Z => n4);
   U4 : INV_X1 port map( A => n7, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : BUF_X1 port map( A => n8, Z => n2);
   U7 : BUF_X1 port map( A => n8, Z => n1);
   U8 : BUF_X1 port map( A => n8, Z => n3);
   U9 : INV_X1 port map( A => n95, ZN => Y(2));
   U10 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n2, ZN => 
                           n95);
   U11 : INV_X1 port map( A => n74, ZN => Y(10));
   U12 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n1, ZN =>
                           n74);
   U13 : INV_X1 port map( A => n75, ZN => Y(11));
   U14 : AOI22_X1 port map( A1 => A(11), A2 => n6, B1 => B(11), B2 => n1, ZN =>
                           n75);
   U15 : INV_X1 port map( A => n76, ZN => Y(12));
   U16 : AOI22_X1 port map( A1 => A(12), A2 => n6, B1 => B(12), B2 => n1, ZN =>
                           n76);
   U17 : INV_X1 port map( A => n77, ZN => Y(13));
   U18 : AOI22_X1 port map( A1 => A(13), A2 => n6, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U19 : INV_X1 port map( A => n78, ZN => Y(14));
   U20 : AOI22_X1 port map( A1 => A(14), A2 => n5, B1 => B(14), B2 => n1, ZN =>
                           n78);
   U21 : INV_X1 port map( A => n79, ZN => Y(15));
   U22 : AOI22_X1 port map( A1 => A(15), A2 => n6, B1 => B(15), B2 => n1, ZN =>
                           n79);
   U23 : INV_X1 port map( A => n80, ZN => Y(16));
   U24 : AOI22_X1 port map( A1 => A(16), A2 => n5, B1 => B(16), B2 => n1, ZN =>
                           n80);
   U25 : INV_X1 port map( A => n81, ZN => Y(17));
   U26 : AOI22_X1 port map( A1 => A(17), A2 => n6, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U27 : INV_X1 port map( A => n82, ZN => Y(18));
   U28 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n1, ZN =>
                           n82);
   U29 : INV_X1 port map( A => n83, ZN => Y(19));
   U30 : AOI22_X1 port map( A1 => A(19), A2 => n6, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U31 : INV_X1 port map( A => n85, ZN => Y(20));
   U32 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U33 : INV_X1 port map( A => n86, ZN => Y(21));
   U34 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n2, ZN =>
                           n86);
   U35 : INV_X1 port map( A => n87, ZN => Y(22));
   U36 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n2, ZN =>
                           n87);
   U37 : INV_X1 port map( A => n88, ZN => Y(23));
   U38 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n2, ZN =>
                           n88);
   U39 : INV_X1 port map( A => n89, ZN => Y(24));
   U40 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n2, ZN =>
                           n89);
   U41 : INV_X1 port map( A => n90, ZN => Y(25));
   U42 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n2, ZN =>
                           n90);
   U43 : INV_X1 port map( A => n91, ZN => Y(26));
   U44 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n2, ZN =>
                           n91);
   U45 : INV_X1 port map( A => n92, ZN => Y(27));
   U46 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n2, ZN =>
                           n92);
   U47 : INV_X1 port map( A => n93, ZN => Y(28));
   U48 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n2, ZN =>
                           n93);
   U49 : INV_X1 port map( A => n94, ZN => Y(29));
   U50 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n2, ZN =>
                           n94);
   U51 : INV_X1 port map( A => n96, ZN => Y(30));
   U52 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n2, ZN =>
                           n96);
   U53 : INV_X1 port map( A => n104, ZN => Y(9));
   U54 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n3, B2 => B(9), ZN => 
                           n104);
   U55 : INV_X1 port map( A => n98, ZN => Y(3));
   U56 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => n3, ZN => 
                           n98);
   U57 : INV_X1 port map( A => n99, ZN => Y(4));
   U58 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n3, ZN => 
                           n99);
   U59 : INV_X1 port map( A => n100, ZN => Y(5));
   U60 : AOI22_X1 port map( A1 => A(5), A2 => n6, B1 => B(5), B2 => n3, ZN => 
                           n100);
   U61 : INV_X1 port map( A => n101, ZN => Y(6));
   U62 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n3, ZN => 
                           n101);
   U63 : INV_X1 port map( A => n102, ZN => Y(7));
   U64 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n3, ZN => 
                           n102);
   U65 : INV_X1 port map( A => n103, ZN => Y(8));
   U66 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n3, ZN => 
                           n103);
   U67 : INV_X1 port map( A => n97, ZN => Y(31));
   U68 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n3, ZN =>
                           n97);
   U69 : AOI22_X1 port map( A1 => A(1), A2 => n6, B1 => B(1), B2 => n1, ZN => 
                           n84);
   U70 : AOI22_X1 port map( A1 => A(0), A2 => n6, B1 => B(0), B2 => n1, ZN => 
                           n73);
   U71 : INV_X1 port map( A => n84, ZN => Y(1));
   U72 : INV_X1 port map( A => n73, ZN => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_3 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_3;

architecture SYN_Behavioral of MUX3to1_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12_port, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n27, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n28, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n73, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n83, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n16, D => n84, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n16, D => n85, Q => Y(0));
   U3 : BUF_X1 port map( A => N12, Z => n17);
   U4 : BUF_X1 port map( A => n119, Z => n8);
   U5 : BUF_X1 port map( A => n120, Z => n12_port);
   U6 : BUF_X1 port map( A => n118, Z => n1);
   U7 : BUF_X1 port map( A => n17, Z => n15);
   U8 : BUF_X1 port map( A => n17, Z => n14);
   U9 : BUF_X1 port map( A => n17, Z => n16);
   U10 : BUF_X1 port map( A => n18, Z => n13);
   U11 : BUF_X1 port map( A => N12, Z => n18);
   U12 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U13 : BUF_X1 port map( A => n8, Z => n6);
   U14 : BUF_X1 port map( A => n8, Z => n5);
   U15 : BUF_X1 port map( A => n1, Z => n2);
   U16 : BUF_X1 port map( A => n1, Z => n3);
   U17 : BUF_X1 port map( A => n12_port, Z => n9);
   U18 : BUF_X1 port map( A => n12_port, Z => n10);
   U19 : BUF_X1 port map( A => n8, Z => n7);
   U20 : BUF_X1 port map( A => n1, Z => n4);
   U21 : BUF_X1 port map( A => n12_port, Z => n11);
   U22 : NOR2_X1 port map( A1 => n86, A2 => SEL(0), ZN => n119);
   U23 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n120);
   U24 : INV_X1 port map( A => SEL(1), ZN => n86);
   U25 : AND2_X1 port map( A1 => SEL(0), A2 => n86, ZN => n118);
   U26 : INV_X1 port map( A => n87, ZN => n85);
   U27 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n87);
   U28 : INV_X1 port map( A => n88, ZN => n84);
   U29 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n88);
   U30 : INV_X1 port map( A => n89, ZN => n83);
   U31 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n89);
   U32 : INV_X1 port map( A => n90, ZN => n82);
   U33 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n90);
   U34 : INV_X1 port map( A => n91, ZN => n81);
   U35 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n91);
   U36 : INV_X1 port map( A => n92, ZN => n80);
   U37 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n92);
   U38 : INV_X1 port map( A => n93, ZN => n79);
   U39 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n93);
   U40 : INV_X1 port map( A => n94, ZN => n78);
   U41 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n94);
   U42 : INV_X1 port map( A => n95, ZN => n77);
   U43 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n95);
   U44 : INV_X1 port map( A => n96, ZN => n76);
   U45 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n96);
   U46 : INV_X1 port map( A => n97, ZN => n75);
   U47 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n97);
   U48 : INV_X1 port map( A => n98, ZN => n74);
   U49 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n98);
   U50 : INV_X1 port map( A => n99, ZN => n73);
   U51 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n99);
   U52 : INV_X1 port map( A => n100, ZN => n72);
   U53 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n100);
   U54 : INV_X1 port map( A => n101, ZN => n71);
   U55 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n101);
   U56 : INV_X1 port map( A => n102, ZN => n70);
   U57 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n102);
   U58 : INV_X1 port map( A => n103, ZN => n69);
   U59 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n103);
   U60 : INV_X1 port map( A => n104, ZN => n33);
   U61 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n104);
   U62 : INV_X1 port map( A => n105, ZN => n32);
   U63 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n105);
   U64 : INV_X1 port map( A => n106, ZN => n31);
   U65 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n106);
   U66 : INV_X1 port map( A => n107, ZN => n30);
   U67 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n107);
   U68 : INV_X1 port map( A => n108, ZN => n29);
   U69 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n108);
   U70 : INV_X1 port map( A => n109, ZN => n28);
   U71 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n109);
   U72 : INV_X1 port map( A => n110, ZN => n27);
   U73 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n110);
   U74 : INV_X1 port map( A => n111, ZN => n26);
   U75 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n111);
   U76 : INV_X1 port map( A => n112, ZN => n25);
   U77 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n112);
   U78 : INV_X1 port map( A => n113, ZN => n24);
   U79 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n113);
   U80 : INV_X1 port map( A => n114, ZN => n23);
   U81 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n114);
   U82 : INV_X1 port map( A => n115, ZN => n22);
   U83 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n115);
   U84 : INV_X1 port map( A => n116, ZN => n21);
   U85 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n116);
   U86 : INV_X1 port map( A => n117, ZN => n20);
   U87 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n117);
   U88 : INV_X1 port map( A => n121, ZN => n19);
   U89 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n121);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_2 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_2;

architecture SYN_Behavioral of MUX3to1_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12_port, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n27, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n28, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n73, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n83, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n16, D => n84, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n16, D => n85, Q => Y(0));
   U3 : BUF_X1 port map( A => N12, Z => n17);
   U4 : BUF_X1 port map( A => n119, Z => n8);
   U5 : BUF_X1 port map( A => n120, Z => n12_port);
   U6 : BUF_X1 port map( A => n118, Z => n1);
   U7 : BUF_X1 port map( A => n17, Z => n15);
   U8 : BUF_X1 port map( A => n17, Z => n14);
   U9 : BUF_X1 port map( A => n17, Z => n16);
   U10 : BUF_X1 port map( A => n18, Z => n13);
   U11 : BUF_X1 port map( A => N12, Z => n18);
   U12 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U13 : BUF_X1 port map( A => n8, Z => n6);
   U14 : BUF_X1 port map( A => n8, Z => n5);
   U15 : BUF_X1 port map( A => n1, Z => n2);
   U16 : BUF_X1 port map( A => n1, Z => n3);
   U17 : BUF_X1 port map( A => n12_port, Z => n9);
   U18 : BUF_X1 port map( A => n12_port, Z => n10);
   U19 : BUF_X1 port map( A => n8, Z => n7);
   U20 : BUF_X1 port map( A => n1, Z => n4);
   U21 : BUF_X1 port map( A => n12_port, Z => n11);
   U22 : NOR2_X1 port map( A1 => n86, A2 => SEL(0), ZN => n119);
   U23 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n120);
   U24 : INV_X1 port map( A => SEL(1), ZN => n86);
   U25 : AND2_X1 port map( A1 => SEL(0), A2 => n86, ZN => n118);
   U26 : INV_X1 port map( A => n87, ZN => n85);
   U27 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n87);
   U28 : INV_X1 port map( A => n88, ZN => n84);
   U29 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n88);
   U30 : INV_X1 port map( A => n89, ZN => n83);
   U31 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n89);
   U32 : INV_X1 port map( A => n90, ZN => n82);
   U33 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n90);
   U34 : INV_X1 port map( A => n91, ZN => n81);
   U35 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n91);
   U36 : INV_X1 port map( A => n92, ZN => n80);
   U37 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n92);
   U38 : INV_X1 port map( A => n93, ZN => n79);
   U39 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n93);
   U40 : INV_X1 port map( A => n94, ZN => n78);
   U41 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n94);
   U42 : INV_X1 port map( A => n95, ZN => n77);
   U43 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n95);
   U44 : INV_X1 port map( A => n96, ZN => n76);
   U45 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n96);
   U46 : INV_X1 port map( A => n97, ZN => n75);
   U47 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n97);
   U48 : INV_X1 port map( A => n98, ZN => n74);
   U49 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n98);
   U50 : INV_X1 port map( A => n99, ZN => n73);
   U51 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n99);
   U52 : INV_X1 port map( A => n100, ZN => n72);
   U53 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n100);
   U54 : INV_X1 port map( A => n101, ZN => n71);
   U55 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n101);
   U56 : INV_X1 port map( A => n102, ZN => n70);
   U57 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n102);
   U58 : INV_X1 port map( A => n103, ZN => n69);
   U59 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n103);
   U60 : INV_X1 port map( A => n104, ZN => n33);
   U61 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n104);
   U62 : INV_X1 port map( A => n105, ZN => n32);
   U63 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n105);
   U64 : INV_X1 port map( A => n106, ZN => n31);
   U65 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n106);
   U66 : INV_X1 port map( A => n107, ZN => n30);
   U67 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n107);
   U68 : INV_X1 port map( A => n108, ZN => n29);
   U69 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n108);
   U70 : INV_X1 port map( A => n109, ZN => n28);
   U71 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n109);
   U72 : INV_X1 port map( A => n110, ZN => n27);
   U73 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n110);
   U74 : INV_X1 port map( A => n111, ZN => n26);
   U75 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n111);
   U76 : INV_X1 port map( A => n112, ZN => n25);
   U77 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n112);
   U78 : INV_X1 port map( A => n113, ZN => n24);
   U79 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n113);
   U80 : INV_X1 port map( A => n114, ZN => n23);
   U81 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n114);
   U82 : INV_X1 port map( A => n115, ZN => n22);
   U83 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n115);
   U84 : INV_X1 port map( A => n116, ZN => n21);
   U85 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n116);
   U86 : INV_X1 port map( A => n117, ZN => n20);
   U87 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n117);
   U88 : INV_X1 port map( A => n121, ZN => n19);
   U89 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n121);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_1 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_1;

architecture SYN_Behavioral of MUX3to1_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12_port, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n13, D => n19, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n13, D => n20, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n13, D => n21, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n13, D => n22, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n13, D => n23, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n13, D => n24, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n13, D => n25, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n13, D => n26, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n13, D => n27, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n13, D => n28, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n14, D => n29, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n14, D => n30, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n14, D => n31, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n14, D => n32, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n14, D => n33, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n14, D => n69, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n14, D => n70, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n14, D => n71, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n14, D => n72, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n14, D => n73, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n15, D => n74, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n15, D => n75, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n15, D => n76, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n15, D => n77, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n15, D => n78, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n15, D => n79, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n15, D => n80, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n15, D => n81, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n15, D => n82, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n15, D => n83, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n16, D => n84, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n16, D => n85, Q => Y(0));
   U3 : BUF_X1 port map( A => N12, Z => n17);
   U4 : BUF_X1 port map( A => n119, Z => n8);
   U5 : BUF_X1 port map( A => n120, Z => n12_port);
   U6 : BUF_X1 port map( A => n118, Z => n1);
   U7 : BUF_X1 port map( A => n17, Z => n15);
   U8 : BUF_X1 port map( A => n17, Z => n14);
   U9 : BUF_X1 port map( A => n17, Z => n16);
   U10 : BUF_X1 port map( A => n18, Z => n13);
   U11 : BUF_X1 port map( A => N12, Z => n18);
   U12 : OR3_X1 port map( A1 => n2, A2 => n9, A3 => n7, ZN => N12);
   U13 : BUF_X1 port map( A => n8, Z => n6);
   U14 : BUF_X1 port map( A => n8, Z => n5);
   U15 : BUF_X1 port map( A => n1, Z => n2);
   U16 : BUF_X1 port map( A => n1, Z => n3);
   U17 : BUF_X1 port map( A => n12_port, Z => n9);
   U18 : BUF_X1 port map( A => n12_port, Z => n10);
   U19 : BUF_X1 port map( A => n8, Z => n7);
   U20 : BUF_X1 port map( A => n1, Z => n4);
   U21 : BUF_X1 port map( A => n12_port, Z => n11);
   U22 : NOR2_X1 port map( A1 => n86, A2 => SEL(0), ZN => n119);
   U23 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n120);
   U24 : INV_X1 port map( A => SEL(1), ZN => n86);
   U25 : AND2_X1 port map( A1 => SEL(0), A2 => n86, ZN => n118);
   U26 : INV_X1 port map( A => n87, ZN => n85);
   U27 : AOI222_X1 port map( A1 => A(0), A2 => n9, B1 => C(0), B2 => n7, C1 => 
                           B(0), C2 => n2, ZN => n87);
   U28 : INV_X1 port map( A => n88, ZN => n84);
   U29 : AOI222_X1 port map( A1 => A(1), A2 => n9, B1 => C(1), B2 => n7, C1 => 
                           B(1), C2 => n2, ZN => n88);
   U30 : INV_X1 port map( A => n89, ZN => n83);
   U31 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => C(2), B2 => n7, C1 => 
                           B(2), C2 => n2, ZN => n89);
   U32 : INV_X1 port map( A => n90, ZN => n82);
   U33 : AOI222_X1 port map( A1 => A(3), A2 => n9, B1 => C(3), B2 => n7, C1 => 
                           B(3), C2 => n2, ZN => n90);
   U34 : INV_X1 port map( A => n91, ZN => n81);
   U35 : AOI222_X1 port map( A1 => A(4), A2 => n9, B1 => C(4), B2 => n7, C1 => 
                           B(4), C2 => n2, ZN => n91);
   U36 : INV_X1 port map( A => n92, ZN => n80);
   U37 : AOI222_X1 port map( A1 => A(5), A2 => n9, B1 => C(5), B2 => n7, C1 => 
                           B(5), C2 => n2, ZN => n92);
   U38 : INV_X1 port map( A => n93, ZN => n79);
   U39 : AOI222_X1 port map( A1 => A(6), A2 => n9, B1 => C(6), B2 => n7, C1 => 
                           B(6), C2 => n2, ZN => n93);
   U40 : INV_X1 port map( A => n94, ZN => n78);
   U41 : AOI222_X1 port map( A1 => A(7), A2 => n9, B1 => C(7), B2 => n7, C1 => 
                           B(7), C2 => n2, ZN => n94);
   U42 : INV_X1 port map( A => n95, ZN => n77);
   U43 : AOI222_X1 port map( A1 => A(8), A2 => n9, B1 => C(8), B2 => n6, C1 => 
                           B(8), C2 => n2, ZN => n95);
   U44 : INV_X1 port map( A => n96, ZN => n76);
   U45 : AOI222_X1 port map( A1 => A(9), A2 => n9, B1 => C(9), B2 => n6, C1 => 
                           B(9), C2 => n2, ZN => n96);
   U46 : INV_X1 port map( A => n97, ZN => n75);
   U47 : AOI222_X1 port map( A1 => A(10), A2 => n9, B1 => C(10), B2 => n6, C1 
                           => B(10), C2 => n2, ZN => n97);
   U48 : INV_X1 port map( A => n98, ZN => n74);
   U49 : AOI222_X1 port map( A1 => A(11), A2 => n10, B1 => C(11), B2 => n6, C1 
                           => B(11), C2 => n3, ZN => n98);
   U50 : INV_X1 port map( A => n99, ZN => n73);
   U51 : AOI222_X1 port map( A1 => A(12), A2 => n10, B1 => C(12), B2 => n6, C1 
                           => B(12), C2 => n3, ZN => n99);
   U52 : INV_X1 port map( A => n100, ZN => n72);
   U53 : AOI222_X1 port map( A1 => A(13), A2 => n10, B1 => C(13), B2 => n6, C1 
                           => B(13), C2 => n3, ZN => n100);
   U54 : INV_X1 port map( A => n101, ZN => n71);
   U55 : AOI222_X1 port map( A1 => A(14), A2 => n10, B1 => C(14), B2 => n6, C1 
                           => B(14), C2 => n3, ZN => n101);
   U56 : INV_X1 port map( A => n102, ZN => n70);
   U57 : AOI222_X1 port map( A1 => A(15), A2 => n10, B1 => C(15), B2 => n6, C1 
                           => B(15), C2 => n3, ZN => n102);
   U58 : INV_X1 port map( A => n103, ZN => n69);
   U59 : AOI222_X1 port map( A1 => A(16), A2 => n10, B1 => C(16), B2 => n6, C1 
                           => B(16), C2 => n3, ZN => n103);
   U60 : INV_X1 port map( A => n104, ZN => n33);
   U61 : AOI222_X1 port map( A1 => A(17), A2 => n10, B1 => C(17), B2 => n6, C1 
                           => B(17), C2 => n3, ZN => n104);
   U62 : INV_X1 port map( A => n105, ZN => n32);
   U63 : AOI222_X1 port map( A1 => A(18), A2 => n10, B1 => C(18), B2 => n6, C1 
                           => B(18), C2 => n3, ZN => n105);
   U64 : INV_X1 port map( A => n106, ZN => n31);
   U65 : AOI222_X1 port map( A1 => A(19), A2 => n10, B1 => C(19), B2 => n6, C1 
                           => B(19), C2 => n3, ZN => n106);
   U66 : INV_X1 port map( A => n107, ZN => n30);
   U67 : AOI222_X1 port map( A1 => A(20), A2 => n10, B1 => C(20), B2 => n5, C1 
                           => B(20), C2 => n3, ZN => n107);
   U68 : INV_X1 port map( A => n108, ZN => n29);
   U69 : AOI222_X1 port map( A1 => A(21), A2 => n10, B1 => C(21), B2 => n5, C1 
                           => B(21), C2 => n3, ZN => n108);
   U70 : INV_X1 port map( A => n109, ZN => n28);
   U71 : AOI222_X1 port map( A1 => A(22), A2 => n10, B1 => C(22), B2 => n5, C1 
                           => B(22), C2 => n3, ZN => n109);
   U72 : INV_X1 port map( A => n110, ZN => n27);
   U73 : AOI222_X1 port map( A1 => A(23), A2 => n11, B1 => C(23), B2 => n5, C1 
                           => B(23), C2 => n4, ZN => n110);
   U74 : INV_X1 port map( A => n111, ZN => n26);
   U75 : AOI222_X1 port map( A1 => A(24), A2 => n11, B1 => C(24), B2 => n5, C1 
                           => B(24), C2 => n4, ZN => n111);
   U76 : INV_X1 port map( A => n112, ZN => n25);
   U77 : AOI222_X1 port map( A1 => A(25), A2 => n11, B1 => C(25), B2 => n5, C1 
                           => B(25), C2 => n4, ZN => n112);
   U78 : INV_X1 port map( A => n113, ZN => n24);
   U79 : AOI222_X1 port map( A1 => A(26), A2 => n11, B1 => C(26), B2 => n5, C1 
                           => B(26), C2 => n4, ZN => n113);
   U80 : INV_X1 port map( A => n114, ZN => n23);
   U81 : AOI222_X1 port map( A1 => A(27), A2 => n11, B1 => C(27), B2 => n5, C1 
                           => B(27), C2 => n4, ZN => n114);
   U82 : INV_X1 port map( A => n115, ZN => n22);
   U83 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => C(28), B2 => n5, C1 
                           => B(28), C2 => n4, ZN => n115);
   U84 : INV_X1 port map( A => n116, ZN => n21);
   U85 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => C(29), B2 => n5, C1 
                           => B(29), C2 => n4, ZN => n116);
   U86 : INV_X1 port map( A => n117, ZN => n20);
   U87 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => C(30), B2 => n5, C1 
                           => B(30), C2 => n4, ZN => n117);
   U88 : INV_X1 port map( A => n121, ZN => n19);
   U89 : AOI222_X1 port map( A1 => A(31), A2 => n11, B1 => C(31), B2 => n5, C1 
                           => B(31), C2 => n4, ZN => n121);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Sum : out std_logic_vector 
         (31 downto 0));

end PC_adder_1;

architecture SYN_Behavioral of PC_adder_1 is

   component PC_adder_1_DW01_add_0_DW01_add_128
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1139 : std_logic;

begin
   
   n2 <= '0';
   add_16 : PC_adder_1_DW01_add_0_DW01_add_128 port map( A(31) => A(31), A(30) 
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => n2, SUM(31) => Sum(31),
                           SUM(30) => Sum(30), SUM(29) => Sum(29), SUM(28) => 
                           Sum(28), SUM(27) => Sum(27), SUM(26) => Sum(26), 
                           SUM(25) => Sum(25), SUM(24) => Sum(24), SUM(23) => 
                           Sum(23), SUM(22) => Sum(22), SUM(21) => Sum(21), 
                           SUM(20) => Sum(20), SUM(19) => Sum(19), SUM(18) => 
                           Sum(18), SUM(17) => Sum(17), SUM(16) => Sum(16), 
                           SUM(15) => Sum(15), SUM(14) => Sum(14), SUM(13) => 
                           Sum(13), SUM(12) => Sum(12), SUM(11) => Sum(11), 
                           SUM(10) => Sum(10), SUM(9) => Sum(9), SUM(8) => 
                           Sum(8), SUM(7) => Sum(7), SUM(6) => Sum(6), SUM(5) 
                           => Sum(5), SUM(4) => Sum(4), SUM(3) => Sum(3), 
                           SUM(2) => Sum(2), SUM(1) => Sum(1), SUM(0) => Sum(0)
                           , CO => n_1139);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FFD_1;

architecture SYN_BEHAVIORAL of FFD_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n5, n6, n7, n8 : std_logic;

begin
   
   Q_reg : SDFFR_X1 port map( D => n5, SI => n6, SE => n3, CK => CK, RN => n7, 
                           Q => Q, QN => n1);
   U2 : INV_X1 port map( A => n1, ZN => n2);
   U3 : INV_X1 port map( A => n8, ZN => n3);
   n5 <= '1';
   n6 <= '0';
   U6 : INV_X1 port map( A => RESET, ZN => n7);
   U7 : MUX2_X1 port map( A => n2, B => D, S => ENABLE, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_17 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_17;

architecture SYN_Behavioral of REG_NBIT32_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n143);
   reg_reg_30_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n144);
   reg_reg_29_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n145);
   reg_reg_26_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n148);
   reg_reg_25_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n149);
   reg_reg_24_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n150);
   reg_reg_23_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n151);
   reg_reg_22_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n152);
   reg_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n153);
   reg_reg_20_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n154);
   reg_reg_19_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n155);
   reg_reg_18_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n156);
   reg_reg_17_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n157);
   reg_reg_16_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n158);
   reg_reg_15_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n159);
   reg_reg_14_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n160);
   reg_reg_13_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n161);
   reg_reg_12_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n162);
   reg_reg_11_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n163);
   reg_reg_10_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n164);
   reg_reg_9_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n165);
   reg_reg_8_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n167);
   reg_reg_6_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n168);
   reg_reg_5_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n169);
   reg_reg_4_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n170);
   reg_reg_3_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n171);
   reg_reg_2_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n172);
   reg_reg_1_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n173);
   reg_reg_0_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n174);
   reg_reg_28_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n110, Q => 
                           data_out(28), QN => n146);
   reg_reg_27_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n110, Q => 
                           data_out(27), QN => n147);
   U2 : BUF_X1 port map( A => n110, Z => n109);
   U3 : BUF_X1 port map( A => n96, Z => n105);
   U4 : BUF_X1 port map( A => n96, Z => n104);
   U5 : BUF_X1 port map( A => n109, Z => n106);
   U6 : BUF_X1 port map( A => n109, Z => n107);
   U7 : BUF_X1 port map( A => n109, Z => n108);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n103);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n101);
   U14 : INV_X1 port map( A => reset, ZN => n110);
   U15 : BUF_X1 port map( A => enable, Z => n96);
   U16 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U17 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n178);
   U18 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U19 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n179);
   U20 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U21 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n199);
   U22 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n197, ZN => n133);
   U23 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n197);
   U24 : OAI21_X1 port map( B1 => n164, B2 => n100, A => n196, ZN => n132);
   U25 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n196);
   U26 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U27 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n195);
   U28 : OAI21_X1 port map( B1 => n162, B2 => n101, A => n194, ZN => n130);
   U29 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n194);
   U30 : OAI21_X1 port map( B1 => n161, B2 => n100, A => n193, ZN => n129);
   U31 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n193);
   U32 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U33 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n192);
   U34 : OAI21_X1 port map( B1 => n159, B2 => n101, A => n191, ZN => n127);
   U35 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n191);
   U36 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U37 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n190);
   U38 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U39 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n189);
   U40 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U41 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n188);
   U42 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U43 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n187);
   U44 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U45 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n186);
   U46 : OAI21_X1 port map( B1 => n153, B2 => n102, A => n185, ZN => n121);
   U47 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n185);
   U48 : OAI21_X1 port map( B1 => n152, B2 => n101, A => n184, ZN => n120);
   U49 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n184);
   U50 : OAI21_X1 port map( B1 => n151, B2 => n102, A => n183, ZN => n119);
   U51 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n183);
   U52 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U53 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n182);
   U54 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U55 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n181);
   U56 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U57 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n180);
   U58 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U59 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n177);
   U60 : OAI21_X1 port map( B1 => n144, B2 => n103, A => n176, ZN => n112);
   U61 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n176);
   U62 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U63 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n175);
   U64 : OAI21_X1 port map( B1 => n173, B2 => n102, A => n205, ZN => n141);
   U65 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n205);
   U66 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U67 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n204);
   U68 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U69 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n203);
   U70 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U71 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n202);
   U72 : OAI21_X1 port map( B1 => n169, B2 => n101, A => n201, ZN => n137);
   U73 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n201);
   U74 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U75 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n200);
   U76 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n198, ZN => n134);
   U77 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n198);
   U78 : OAI21_X1 port map( B1 => n174, B2 => n103, A => n206, ZN => n142);
   U79 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n206);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_16 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_16;

architecture SYN_Behavioral of REG_NBIT32_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, 
      n28, n29, n30, n31, n32, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_28_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n25, Q => 
                           data_out_28_port, QN => n_1140);
   reg_reg_26_inst : DFFR_X1 port map( D => n50, CK => clk, RN => n25, Q => 
                           data_out_26_port, QN => n_1141);
   reg_reg_25_inst : DFFR_X1 port map( D => n51, CK => clk, RN => n26, Q => 
                           data_out_25_port, QN => n_1142);
   reg_reg_24_inst : DFFR_X1 port map( D => n52, CK => clk, RN => n26, Q => 
                           data_out_24_port, QN => n_1143);
   reg_reg_23_inst : DFFR_X1 port map( D => n53, CK => clk, RN => n26, Q => 
                           data_out_23_port, QN => n_1144);
   reg_reg_22_inst : DFFR_X1 port map( D => n54, CK => clk, RN => n26, Q => 
                           data_out_22_port, QN => n_1145);
   reg_reg_21_inst : DFFR_X1 port map( D => n55, CK => clk, RN => n26, Q => 
                           data_out_21_port, QN => n_1146);
   reg_reg_20_inst : DFFR_X1 port map( D => n56, CK => clk, RN => n26, Q => 
                           data_out_20_port, QN => n_1147);
   reg_reg_19_inst : DFFR_X1 port map( D => n57, CK => clk, RN => n26, Q => 
                           data_out_19_port, QN => n_1148);
   reg_reg_18_inst : DFFR_X1 port map( D => n58, CK => clk, RN => n26, Q => 
                           data_out_18_port, QN => n_1149);
   reg_reg_17_inst : DFFR_X1 port map( D => n59, CK => clk, RN => n26, Q => 
                           data_out_17_port, QN => n_1150);
   reg_reg_16_inst : DFFR_X1 port map( D => n60, CK => clk, RN => n26, Q => 
                           data_out_16_port, QN => n_1151);
   reg_reg_15_inst : DFFR_X1 port map( D => n61, CK => clk, RN => n24, Q => 
                           data_out_15_port, QN => n89);
   reg_reg_14_inst : DFFR_X1 port map( D => n62, CK => clk, RN => n24, Q => 
                           data_out_14_port, QN => n90);
   reg_reg_13_inst : DFFR_X1 port map( D => n63, CK => clk, RN => n24, Q => 
                           data_out_13_port, QN => n91);
   reg_reg_12_inst : DFFR_X1 port map( D => n64, CK => clk, RN => n24, Q => 
                           data_out_12_port, QN => n92);
   reg_reg_11_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n24, Q => 
                           data_out_11_port, QN => n93);
   reg_reg_10_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n24, Q => 
                           data_out_10_port, QN => n94);
   reg_reg_9_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n24, Q => 
                           data_out_9_port, QN => n95);
   reg_reg_8_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n24, Q => 
                           data_out_8_port, QN => n96);
   reg_reg_7_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n24, Q => 
                           data_out_7_port, QN => n97);
   reg_reg_6_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n24, Q => 
                           data_out_6_port, QN => n98);
   reg_reg_5_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n24, Q => 
                           data_out_5_port, QN => n99);
   reg_reg_4_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n25, Q => 
                           data_out_4_port, QN => n100);
   reg_reg_3_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n25, Q => 
                           data_out_3_port, QN => n101);
   reg_reg_2_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n25, Q => 
                           data_out_2_port, QN => n102);
   reg_reg_1_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n25, Q => 
                           data_out_1_port, QN => n103);
   reg_reg_0_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n25, Q => 
                           data_out_0_port, QN => n104);
   reg_reg_27_inst : DFFR_X1 port map( D => n49, CK => clk, RN => n28, Q => 
                           data_out_27_port, QN => n_1152);
   reg_reg_29_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n28, Q => 
                           data_out_29_port, QN => n_1153);
   reg_reg_30_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n28, Q => 
                           data_out_30_port, QN => n_1154);
   reg_reg_31_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n28, Q => 
                           data_out_31_port, QN => n_1155);
   U2 : BUF_X1 port map( A => n17, Z => n22);
   U3 : BUF_X1 port map( A => n28, Z => n27);
   U4 : BUF_X1 port map( A => n22, Z => n19);
   U5 : BUF_X1 port map( A => n22, Z => n20);
   U6 : BUF_X1 port map( A => n22, Z => n21);
   U7 : BUF_X1 port map( A => n27, Z => n24);
   U8 : BUF_X1 port map( A => n27, Z => n25);
   U9 : BUF_X1 port map( A => n27, Z => n26);
   U10 : BUF_X1 port map( A => n23, Z => n18);
   U11 : BUF_X1 port map( A => n17, Z => n23);
   U12 : INV_X1 port map( A => reset, ZN => n28);
   U13 : BUF_X1 port map( A => enable, Z => n17);
   U14 : OAI21_X1 port map( B1 => n103, B2 => n19, A => n119, ZN => n87);
   U15 : NAND2_X1 port map( A1 => data_in(1), A2 => n19, ZN => n119);
   U16 : OAI21_X1 port map( B1 => n102, B2 => n19, A => n118, ZN => n86);
   U17 : NAND2_X1 port map( A1 => data_in(2), A2 => n19, ZN => n118);
   U18 : OAI21_X1 port map( B1 => n101, B2 => n19, A => n117, ZN => n85);
   U19 : NAND2_X1 port map( A1 => data_in(3), A2 => n19, ZN => n117);
   U20 : OAI21_X1 port map( B1 => n104, B2 => n19, A => n120, ZN => n88);
   U21 : NAND2_X1 port map( A1 => n20, A2 => data_in(0), ZN => n120);
   U22 : OAI21_X1 port map( B1 => n89, B2 => n20, A => n105, ZN => n61);
   U23 : NAND2_X1 port map( A1 => data_in(15), A2 => n18, ZN => n105);
   U24 : OAI21_X1 port map( B1 => n95, B2 => n20, A => n111, ZN => n79);
   U25 : NAND2_X1 port map( A1 => data_in(9), A2 => n18, ZN => n111);
   U26 : OAI21_X1 port map( B1 => n94, B2 => n20, A => n110, ZN => n78);
   U27 : NAND2_X1 port map( A1 => data_in(10), A2 => n18, ZN => n110);
   U28 : OAI21_X1 port map( B1 => n93, B2 => n20, A => n109, ZN => n77);
   U29 : NAND2_X1 port map( A1 => data_in(11), A2 => n18, ZN => n109);
   U30 : OAI21_X1 port map( B1 => n92, B2 => n20, A => n108, ZN => n64);
   U31 : NAND2_X1 port map( A1 => data_in(12), A2 => n18, ZN => n108);
   U32 : OAI21_X1 port map( B1 => n91, B2 => n20, A => n107, ZN => n63);
   U33 : NAND2_X1 port map( A1 => data_in(13), A2 => n18, ZN => n107);
   U34 : OAI21_X1 port map( B1 => n90, B2 => n20, A => n106, ZN => n62);
   U35 : NAND2_X1 port map( A1 => data_in(14), A2 => n18, ZN => n106);
   U36 : OAI21_X1 port map( B1 => n100, B2 => n19, A => n116, ZN => n84);
   U37 : NAND2_X1 port map( A1 => data_in(4), A2 => n18, ZN => n116);
   U38 : OAI21_X1 port map( B1 => n99, B2 => n19, A => n115, ZN => n83);
   U39 : NAND2_X1 port map( A1 => data_in(5), A2 => n18, ZN => n115);
   U40 : OAI21_X1 port map( B1 => n98, B2 => n19, A => n114, ZN => n82);
   U41 : NAND2_X1 port map( A1 => data_in(6), A2 => n18, ZN => n114);
   U42 : OAI21_X1 port map( B1 => n97, B2 => n19, A => n113, ZN => n81);
   U43 : NAND2_X1 port map( A1 => data_in(7), A2 => n18, ZN => n113);
   U44 : OAI21_X1 port map( B1 => n96, B2 => n19, A => n112, ZN => n80);
   U45 : NAND2_X1 port map( A1 => data_in(8), A2 => n18, ZN => n112);
   U46 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => n21, Z
                           => n60);
   U47 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => n21, Z
                           => n59);
   U48 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => n21, Z
                           => n58);
   U49 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => n21, Z
                           => n57);
   U50 : MUX2_X1 port map( A => data_out_20_port, B => data_in(20), S => n21, Z
                           => n56);
   U51 : MUX2_X1 port map( A => data_out_21_port, B => data_in(21), S => n21, Z
                           => n55);
   U52 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => n21, Z
                           => n54);
   U53 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => n21, Z
                           => n53);
   U54 : MUX2_X1 port map( A => data_out_24_port, B => data_in(24), S => n21, Z
                           => n52);
   U55 : MUX2_X1 port map( A => data_out_25_port, B => data_in(25), S => n21, Z
                           => n51);
   U56 : MUX2_X1 port map( A => data_out_26_port, B => data_in(26), S => n20, Z
                           => n50);
   U57 : MUX2_X1 port map( A => data_out_27_port, B => data_in(27), S => n20, Z
                           => n49);
   U58 : MUX2_X1 port map( A => data_out_28_port, B => data_in(28), S => n20, Z
                           => n32);
   U59 : MUX2_X1 port map( A => data_out_29_port, B => data_in(29), S => n20, Z
                           => n31);
   U60 : MUX2_X1 port map( A => data_out_30_port, B => data_in(30), S => n20, Z
                           => n30);
   U61 : MUX2_X1 port map( A => data_out_31_port, B => data_in(31), S => n20, Z
                           => n29);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_15 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_15;

architecture SYN_Behavioral of REG_NBIT32_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_14 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_14;

architecture SYN_Behavioral of REG_NBIT32_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_13 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_13;

architecture SYN_Behavioral of REG_NBIT32_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n27, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n105, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n105, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n105, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n105, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n105, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n107, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n105, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n105, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n105, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n105, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n105, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n105, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n106, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n106, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n106, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n106, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n106, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n106, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n106, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n106, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n106, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n107, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n107, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n107, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n107, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n107, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n107, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n107, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n107, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n107, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n27, Z => n104);
   U3 : BUF_X1 port map( A => n27, Z => n103);
   U4 : BUF_X1 port map( A => n108, Z => n106);
   U5 : BUF_X1 port map( A => n108, Z => n105);
   U6 : BUF_X1 port map( A => n108, Z => n107);
   U7 : INV_X1 port map( A => reset, ZN => n108);
   U8 : BUF_X1 port map( A => n104, Z => n98);
   U9 : BUF_X1 port map( A => n104, Z => n96);
   U10 : BUF_X1 port map( A => n104, Z => n99);
   U11 : BUF_X1 port map( A => n103, Z => n100);
   U12 : BUF_X1 port map( A => n103, Z => n101);
   U13 : BUF_X1 port map( A => n103, Z => n102);
   U14 : BUF_X1 port map( A => enable, Z => n27);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n101, A => n204, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n102, A2 => data_in(0), ZN => n204);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n101, A => n203, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n99, ZN => n203);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n101, A => n202, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n99, ZN => n202);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n101, A => n201, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n99, ZN => n201);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n101, A => n200, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n99, ZN => n200);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n100, A => n199, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n98, ZN => n199);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n100, A => n198, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n99, ZN => n198);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n197, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n197);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n99, A => n196, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n98, ZN => n196);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n99, A => n195, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n98, ZN => n195);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n99, A => n194, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n98, ZN => n194);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n193, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n98, ZN => n193);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n99, A => n192, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n98, ZN => n192);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n99, A => n191, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n98, ZN => n191);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n190, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n98, ZN => n190);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n99, A => n189, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n98, ZN => n189);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n100, A => n188, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n98, ZN => n188);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n100, A => n187, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n98, ZN => n187);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n100, A => n186, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n98, ZN => n186);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n100, A => n185, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n96, ZN => n185);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n100, A => n184, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n96, ZN => n184);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n100, A => n183, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n96, ZN => n183);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n100, A => n182, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n96, ZN => n182);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n101, A => n181, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n96, ZN => n181);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n101, A => n180, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n96, ZN => n180);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n101, A => n179, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n96, ZN => n179);
   U67 : OAI21_X1 port map( B1 => n146, B2 => n101, A => n178, ZN => n114);
   U68 : NAND2_X1 port map( A1 => data_in(27), A2 => n96, ZN => n178);
   U69 : OAI21_X1 port map( B1 => n145, B2 => n101, A => n177, ZN => n113);
   U70 : NAND2_X1 port map( A1 => data_in(28), A2 => n96, ZN => n177);
   U71 : OAI21_X1 port map( B1 => n144, B2 => n101, A => n176, ZN => n112);
   U72 : NAND2_X1 port map( A1 => data_in(29), A2 => n96, ZN => n176);
   U73 : OAI21_X1 port map( B1 => n143, B2 => n101, A => n175, ZN => n111);
   U74 : NAND2_X1 port map( A1 => data_in(30), A2 => n96, ZN => n175);
   U75 : OAI21_X1 port map( B1 => n142, B2 => n102, A => n174, ZN => n110);
   U76 : NAND2_X1 port map( A1 => data_in(31), A2 => n96, ZN => n174);
   U77 : INV_X1 port map( A => n147, ZN => n109);
   U78 : MUX2_X1 port map( A => n109, B => data_in(26), S => n102, Z => n115);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_12 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_12;

architecture SYN_Behavioral of REG_NBIT32_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_31_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n8, Q => 
                           data_out_31_port, QN => n103);
   reg_reg_30_inst : DFFR_X1 port map( D => n33, CK => clk, RN => n8, Q => 
                           data_out_30_port, QN => n104);
   reg_reg_29_inst : DFFR_X1 port map( D => n34, CK => clk, RN => n8, Q => 
                           data_out_29_port, QN => n105);
   reg_reg_28_inst : DFFR_X1 port map( D => n35, CK => clk, RN => n8, Q => 
                           data_out_28_port, QN => n106);
   reg_reg_27_inst : DFFR_X1 port map( D => n36, CK => clk, RN => n8, Q => 
                           data_out_27_port, QN => n107);
   reg_reg_26_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n8, Q => 
                           data_out_26_port, QN => n108);
   reg_reg_25_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n8, Q => 
                           data_out_25_port, QN => n109);
   reg_reg_24_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n8, Q => 
                           data_out_24_port, QN => n110);
   reg_reg_23_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n8, Q => 
                           data_out_23_port, QN => n111);
   reg_reg_22_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n8, Q => 
                           data_out_22_port, QN => n112);
   reg_reg_21_inst : DFFR_X1 port map( D => n42, CK => clk, RN => n8, Q => 
                           data_out_21_port, QN => n113);
   reg_reg_20_inst : DFFR_X1 port map( D => n43, CK => clk, RN => n9, Q => 
                           data_out_20_port, QN => n114);
   reg_reg_19_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n9, Q => 
                           data_out_19_port, QN => n115);
   reg_reg_18_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n9, Q => 
                           data_out_18_port, QN => n116);
   reg_reg_17_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n9, Q => 
                           data_out_17_port, QN => n117);
   reg_reg_16_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n9, Q => 
                           data_out_16_port, QN => n118);
   reg_reg_15_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n9, Q => 
                           data_out_15_port, QN => n119);
   reg_reg_14_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n9, Q => 
                           data_out_14_port, QN => n120);
   reg_reg_13_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n9, Q => 
                           data_out_13_port, QN => n121);
   reg_reg_12_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n9, Q => 
                           data_out_12_port, QN => n122);
   reg_reg_11_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n9, Q => 
                           data_out_11_port, QN => n_1156);
   reg_reg_10_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n9, Q => 
                           data_out_10_port, QN => n_1157);
   reg_reg_9_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n10, Q => 
                           data_out_9_port, QN => n_1158);
   reg_reg_8_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n10, Q => 
                           data_out_8_port, QN => n_1159);
   reg_reg_7_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n10, Q => 
                           data_out_7_port, QN => n_1160);
   reg_reg_6_inst : DFFR_X1 port map( D => n96, CK => clk, RN => n10, Q => 
                           data_out_6_port, QN => n_1161);
   reg_reg_5_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n10, Q => 
                           data_out_5_port, QN => n_1162);
   reg_reg_4_inst : DFFR_X1 port map( D => n98, CK => clk, RN => n10, Q => 
                           data_out_4_port, QN => n_1163);
   reg_reg_3_inst : DFFR_X1 port map( D => n99, CK => clk, RN => n10, Q => 
                           data_out_3_port, QN => n_1164);
   reg_reg_2_inst : DFFR_X1 port map( D => n100, CK => clk, RN => n10, Q => 
                           data_out_2_port, QN => n_1165);
   reg_reg_1_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n10, Q => 
                           data_out_1_port, QN => n_1166);
   reg_reg_0_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n10, Q => 
                           data_out_0_port, QN => n_1167);
   U2 : BUF_X1 port map( A => n1, Z => n6);
   U3 : BUF_X1 port map( A => n11, Z => n9);
   U4 : BUF_X1 port map( A => n11, Z => n8);
   U5 : BUF_X1 port map( A => n11, Z => n10);
   U6 : INV_X1 port map( A => reset, ZN => n11);
   U7 : BUF_X1 port map( A => n6, Z => n3);
   U8 : BUF_X1 port map( A => n6, Z => n4);
   U9 : BUF_X1 port map( A => n6, Z => n5);
   U10 : BUF_X1 port map( A => n7, Z => n2);
   U11 : BUF_X1 port map( A => n1, Z => n7);
   U12 : BUF_X1 port map( A => enable, Z => n1);
   U13 : OAI21_X1 port map( B1 => n122, B2 => n4, A => n142, ZN => n90);
   U14 : NAND2_X1 port map( A1 => data_in(12), A2 => n3, ZN => n142);
   U15 : OAI21_X1 port map( B1 => n121, B2 => n4, A => n141, ZN => n89);
   U16 : NAND2_X1 port map( A1 => data_in(13), A2 => n3, ZN => n141);
   U17 : OAI21_X1 port map( B1 => n120, B2 => n3, A => n140, ZN => n88);
   U18 : NAND2_X1 port map( A1 => data_in(14), A2 => n3, ZN => n140);
   U19 : OAI21_X1 port map( B1 => n119, B2 => n3, A => n139, ZN => n87);
   U20 : NAND2_X1 port map( A1 => data_in(15), A2 => n3, ZN => n139);
   U21 : OAI21_X1 port map( B1 => n118, B2 => n3, A => n138, ZN => n86);
   U22 : NAND2_X1 port map( A1 => data_in(16), A2 => n3, ZN => n138);
   U23 : OAI21_X1 port map( B1 => n117, B2 => n3, A => n137, ZN => n85);
   U24 : NAND2_X1 port map( A1 => data_in(17), A2 => n3, ZN => n137);
   U25 : OAI21_X1 port map( B1 => n116, B2 => n4, A => n136, ZN => n84);
   U26 : NAND2_X1 port map( A1 => data_in(18), A2 => n3, ZN => n136);
   U27 : OAI21_X1 port map( B1 => n115, B2 => n4, A => n135, ZN => n44);
   U28 : NAND2_X1 port map( A1 => data_in(19), A2 => n2, ZN => n135);
   U29 : OAI21_X1 port map( B1 => n114, B2 => n4, A => n134, ZN => n43);
   U30 : NAND2_X1 port map( A1 => data_in(20), A2 => n2, ZN => n134);
   U31 : OAI21_X1 port map( B1 => n113, B2 => n4, A => n133, ZN => n42);
   U32 : NAND2_X1 port map( A1 => data_in(21), A2 => n2, ZN => n133);
   U33 : OAI21_X1 port map( B1 => n112, B2 => n4, A => n132, ZN => n41);
   U34 : NAND2_X1 port map( A1 => data_in(22), A2 => n2, ZN => n132);
   U35 : OAI21_X1 port map( B1 => n111, B2 => n4, A => n131, ZN => n40);
   U36 : NAND2_X1 port map( A1 => data_in(23), A2 => n2, ZN => n131);
   U37 : OAI21_X1 port map( B1 => n110, B2 => n4, A => n130, ZN => n39);
   U38 : NAND2_X1 port map( A1 => data_in(24), A2 => n2, ZN => n130);
   U39 : OAI21_X1 port map( B1 => n109, B2 => n4, A => n129, ZN => n38);
   U40 : NAND2_X1 port map( A1 => data_in(25), A2 => n2, ZN => n129);
   U41 : OAI21_X1 port map( B1 => n108, B2 => n4, A => n128, ZN => n37);
   U42 : NAND2_X1 port map( A1 => data_in(26), A2 => n2, ZN => n128);
   U43 : OAI21_X1 port map( B1 => n107, B2 => n4, A => n127, ZN => n36);
   U44 : NAND2_X1 port map( A1 => data_in(27), A2 => n2, ZN => n127);
   U45 : OAI21_X1 port map( B1 => n106, B2 => n5, A => n126, ZN => n35);
   U46 : NAND2_X1 port map( A1 => data_in(28), A2 => n2, ZN => n126);
   U47 : OAI21_X1 port map( B1 => n105, B2 => n5, A => n125, ZN => n34);
   U48 : NAND2_X1 port map( A1 => data_in(29), A2 => n2, ZN => n125);
   U49 : OAI21_X1 port map( B1 => n104, B2 => n5, A => n124, ZN => n33);
   U50 : NAND2_X1 port map( A1 => data_in(30), A2 => n2, ZN => n124);
   U51 : OAI21_X1 port map( B1 => n103, B2 => n5, A => n123, ZN => n12);
   U52 : NAND2_X1 port map( A1 => data_in(31), A2 => n3, ZN => n123);
   U53 : MUX2_X1 port map( A => data_out_0_port, B => data_in(0), S => n5, Z =>
                           n102);
   U54 : MUX2_X1 port map( A => data_out_1_port, B => data_in(1), S => n5, Z =>
                           n101);
   U55 : MUX2_X1 port map( A => data_out_2_port, B => data_in(2), S => n5, Z =>
                           n100);
   U56 : MUX2_X1 port map( A => data_out_3_port, B => data_in(3), S => n5, Z =>
                           n99);
   U57 : MUX2_X1 port map( A => data_out_4_port, B => data_in(4), S => n5, Z =>
                           n98);
   U58 : MUX2_X1 port map( A => data_out_5_port, B => data_in(5), S => n5, Z =>
                           n97);
   U59 : MUX2_X1 port map( A => data_out_6_port, B => data_in(6), S => n5, Z =>
                           n96);
   U60 : MUX2_X1 port map( A => data_out_7_port, B => data_in(7), S => n5, Z =>
                           n95);
   U61 : MUX2_X1 port map( A => data_out_8_port, B => data_in(8), S => n5, Z =>
                           n94);
   U62 : MUX2_X1 port map( A => data_out_9_port, B => data_in(9), S => n5, Z =>
                           n93);
   U63 : MUX2_X1 port map( A => data_out_10_port, B => data_in(10), S => n5, Z 
                           => n92);
   U64 : MUX2_X1 port map( A => data_out_11_port, B => data_in(11), S => n5, Z 
                           => n91);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_11 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_11;

architecture SYN_Behavioral of REG_NBIT32_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_10 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_10;

architecture SYN_Behavioral of REG_NBIT32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_9 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_9;

architecture SYN_Behavioral of REG_NBIT32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_8 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_8;

architecture SYN_Behavioral of REG_NBIT32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_7 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_7;

architecture SYN_Behavioral of REG_NBIT32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n100);
   U9 : BUF_X1 port map( A => n104, Z => n101);
   U10 : BUF_X1 port map( A => n105, Z => n99);
   U11 : BUF_X1 port map( A => n105, Z => n98);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U16 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U17 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U18 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U19 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U20 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U21 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U22 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U23 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U24 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U25 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U26 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U27 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U28 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U29 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U30 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U31 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U32 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U33 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U34 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U35 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U36 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U37 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U38 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U39 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U40 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U41 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U42 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U46 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U47 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U48 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U49 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U50 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U51 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U52 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U53 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U54 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U55 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U56 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U57 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U58 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U59 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U60 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U61 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);
   U62 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U63 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U64 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U65 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U66 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U67 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U68 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U69 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U70 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U71 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U72 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U73 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U74 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U75 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U76 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U77 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U78 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_6 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_6;

architecture SYN_Behavioral of REG_NBIT32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : INV_X1 port map( A => reset, ZN => n109);
   U8 : BUF_X1 port map( A => n105, Z => n98);
   U9 : BUF_X1 port map( A => n105, Z => n99);
   U10 : BUF_X1 port map( A => n105, Z => n100);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : BUF_X1 port map( A => n104, Z => n103);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U16 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);
   U17 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U18 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U19 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U20 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U21 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U22 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U23 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U24 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U25 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U26 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U27 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U28 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U29 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U30 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U31 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U32 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U33 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U34 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U35 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U36 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U37 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U38 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U39 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U40 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U41 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U42 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U43 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U44 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U45 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U46 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U47 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U48 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U49 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U50 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U51 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U52 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U53 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U54 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U55 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U56 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U57 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U58 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U59 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U60 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U61 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U62 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U63 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U64 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U65 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U66 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U67 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U68 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U69 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U70 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U71 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U72 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U73 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U74 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U75 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U76 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U77 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U78 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_5 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_5;

architecture SYN_Behavioral of REG_NBIT32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : BUF_X1 port map( A => n105, Z => n98);
   U8 : BUF_X1 port map( A => n105, Z => n99);
   U9 : BUF_X1 port map( A => n105, Z => n100);
   U10 : BUF_X1 port map( A => n104, Z => n103);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : INV_X1 port map( A => reset, ZN => n109);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U16 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U17 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U18 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U19 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U20 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U21 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U22 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U23 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U24 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U25 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U26 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U27 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U28 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U29 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U30 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U31 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U32 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U33 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U34 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U35 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U36 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U37 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U38 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U39 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U40 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U41 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U42 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U43 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U44 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U45 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U46 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U47 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U48 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U49 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U50 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U51 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U52 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U53 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U54 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U55 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U56 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U57 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U58 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U59 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U60 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);
   U61 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U62 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U63 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U64 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U65 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U66 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U67 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U68 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U69 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U70 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U71 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U72 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U73 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U74 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U75 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U76 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U77 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U78 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_4 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_4;

architecture SYN_Behavioral of REG_NBIT32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n108, Q => 
                           data_out(31), QN => n142);
   reg_reg_30_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n108, Q => 
                           data_out(30), QN => n143);
   reg_reg_29_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n108, Q => 
                           data_out(29), QN => n144);
   reg_reg_28_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n108, Q => 
                           data_out(28), QN => n145);
   reg_reg_27_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n108, Q => 
                           data_out(27), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n108, Q => 
                           data_out(26), QN => n147);
   reg_reg_25_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n108, Q => 
                           data_out(25), QN => n148);
   reg_reg_24_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n108, Q => 
                           data_out(24), QN => n149);
   reg_reg_23_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n108, Q => 
                           data_out(23), QN => n150);
   reg_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n108, Q => 
                           data_out(22), QN => n151);
   reg_reg_21_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n107, Q => 
                           data_out(21), QN => n152);
   reg_reg_20_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n107, Q => 
                           data_out(20), QN => n153);
   reg_reg_19_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n107, Q => 
                           data_out(19), QN => n154);
   reg_reg_18_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n107, Q => 
                           data_out(18), QN => n155);
   reg_reg_17_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n107, Q => 
                           data_out(17), QN => n156);
   reg_reg_16_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n107, Q => 
                           data_out(16), QN => n157);
   reg_reg_15_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n107, Q => 
                           data_out(15), QN => n158);
   reg_reg_14_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n107, Q => 
                           data_out(14), QN => n159);
   reg_reg_13_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n107, Q => 
                           data_out(13), QN => n160);
   reg_reg_12_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n107, Q => 
                           data_out(12), QN => n161);
   reg_reg_11_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n107, Q => 
                           data_out(11), QN => n162);
   reg_reg_10_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n106, Q => 
                           data_out(10), QN => n163);
   reg_reg_9_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n106, Q => 
                           data_out(9), QN => n164);
   reg_reg_8_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n106, Q => 
                           data_out(8), QN => n165);
   reg_reg_7_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n106, Q => 
                           data_out(7), QN => n166);
   reg_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n106, Q => 
                           data_out(6), QN => n167);
   reg_reg_5_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n106, Q => 
                           data_out(5), QN => n168);
   reg_reg_4_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n106, Q => 
                           data_out(4), QN => n169);
   reg_reg_3_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n106, Q => 
                           data_out(3), QN => n170);
   reg_reg_2_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n106, Q => 
                           data_out(2), QN => n171);
   reg_reg_1_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n106, Q => 
                           data_out(1), QN => n172);
   reg_reg_0_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n106, Q => 
                           data_out(0), QN => n173);
   U2 : BUF_X1 port map( A => n96, Z => n105);
   U3 : BUF_X1 port map( A => n96, Z => n104);
   U4 : BUF_X1 port map( A => n109, Z => n106);
   U5 : BUF_X1 port map( A => n109, Z => n107);
   U6 : BUF_X1 port map( A => n109, Z => n108);
   U7 : BUF_X1 port map( A => n105, Z => n98);
   U8 : BUF_X1 port map( A => n105, Z => n99);
   U9 : BUF_X1 port map( A => n105, Z => n100);
   U10 : BUF_X1 port map( A => n104, Z => n103);
   U11 : BUF_X1 port map( A => n104, Z => n101);
   U12 : BUF_X1 port map( A => n104, Z => n102);
   U13 : INV_X1 port map( A => reset, ZN => n109);
   U14 : BUF_X1 port map( A => enable, Z => n96);
   U15 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n198, ZN => n134);
   U16 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n198);
   U17 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n196, ZN => n132);
   U18 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n196);
   U19 : OAI21_X1 port map( B1 => n163, B2 => n100, A => n195, ZN => n131);
   U20 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n195);
   U21 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n194, ZN => n130);
   U22 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n194);
   U23 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n193, ZN => n129);
   U24 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n193);
   U25 : OAI21_X1 port map( B1 => n160, B2 => n100, A => n192, ZN => n128);
   U26 : NAND2_X1 port map( A1 => data_in(13), A2 => n99, ZN => n192);
   U27 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n191, ZN => n127);
   U28 : NAND2_X1 port map( A1 => data_in(14), A2 => n99, ZN => n191);
   U29 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n190, ZN => n126);
   U30 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n190);
   U31 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n189, ZN => n125);
   U32 : NAND2_X1 port map( A1 => data_in(16), A2 => n99, ZN => n189);
   U33 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n188, ZN => n124);
   U34 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n188);
   U35 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n187, ZN => n123);
   U36 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n187);
   U37 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n186, ZN => n122);
   U38 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n186);
   U39 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n185, ZN => n121);
   U40 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n185);
   U41 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n184, ZN => n120);
   U42 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n184);
   U43 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n183, ZN => n119);
   U44 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n183);
   U45 : OAI21_X1 port map( B1 => n150, B2 => n102, A => n182, ZN => n118);
   U46 : NAND2_X1 port map( A1 => data_in(23), A2 => n98, ZN => n182);
   U47 : OAI21_X1 port map( B1 => n149, B2 => n102, A => n181, ZN => n117);
   U48 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n181);
   U49 : OAI21_X1 port map( B1 => n148, B2 => n102, A => n180, ZN => n116);
   U50 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n180);
   U51 : OAI21_X1 port map( B1 => n147, B2 => n102, A => n179, ZN => n115);
   U52 : NAND2_X1 port map( A1 => data_in(26), A2 => n98, ZN => n179);
   U53 : OAI21_X1 port map( B1 => n146, B2 => n102, A => n178, ZN => n114);
   U54 : NAND2_X1 port map( A1 => data_in(27), A2 => n98, ZN => n178);
   U55 : OAI21_X1 port map( B1 => n145, B2 => n102, A => n177, ZN => n113);
   U56 : NAND2_X1 port map( A1 => data_in(28), A2 => n98, ZN => n177);
   U57 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n176, ZN => n112);
   U58 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n176);
   U59 : OAI21_X1 port map( B1 => n143, B2 => n103, A => n175, ZN => n111);
   U60 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n175);
   U61 : OAI21_X1 port map( B1 => n142, B2 => n103, A => n174, ZN => n110);
   U62 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n174);
   U63 : OAI21_X1 port map( B1 => n172, B2 => n102, A => n204, ZN => n140);
   U64 : NAND2_X1 port map( A1 => data_in(1), A2 => n100, ZN => n204);
   U65 : OAI21_X1 port map( B1 => n171, B2 => n102, A => n203, ZN => n139);
   U66 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n203);
   U67 : OAI21_X1 port map( B1 => n170, B2 => n102, A => n202, ZN => n138);
   U68 : NAND2_X1 port map( A1 => data_in(3), A2 => n100, ZN => n202);
   U69 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n201, ZN => n137);
   U70 : NAND2_X1 port map( A1 => data_in(4), A2 => n100, ZN => n201);
   U71 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n200, ZN => n136);
   U72 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n200);
   U73 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n199, ZN => n135);
   U74 : NAND2_X1 port map( A1 => data_in(6), A2 => n100, ZN => n199);
   U75 : OAI21_X1 port map( B1 => n165, B2 => n100, A => n197, ZN => n133);
   U76 : NAND2_X1 port map( A1 => data_in(8), A2 => n100, ZN => n197);
   U77 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n205, ZN => n141);
   U78 : NAND2_X1 port map( A1 => n103, A2 => data_in(0), ZN => n205);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_3 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_3;

architecture SYN_Behavioral of REG_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196 : std_logic;

begin
   
   reg_reg_31_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n96, Q => 
                           data_out(31), QN => n133);
   reg_reg_30_inst : DFFR_X1 port map( D => n102, CK => clk, RN => n96, Q => 
                           data_out(30), QN => n134);
   reg_reg_29_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n96, Q => 
                           data_out(29), QN => n135);
   reg_reg_28_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n96, Q => 
                           data_out(28), QN => n136);
   reg_reg_27_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n96, Q => 
                           data_out(27), QN => n137);
   reg_reg_26_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n96, Q => 
                           data_out(26), QN => n138);
   reg_reg_25_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n96, Q => 
                           data_out(25), QN => n139);
   reg_reg_24_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n96, Q => 
                           data_out(24), QN => n140);
   reg_reg_23_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n96, Q => 
                           data_out(23), QN => n141);
   reg_reg_22_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n96, Q => 
                           data_out(22), QN => n142);
   reg_reg_21_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n96, Q => 
                           data_out(21), QN => n143);
   reg_reg_20_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n98, Q => 
                           data_out(20), QN => n144);
   reg_reg_19_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n98, Q => 
                           data_out(19), QN => n145);
   reg_reg_18_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n98, Q => 
                           data_out(18), QN => n146);
   reg_reg_17_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n98, Q => 
                           data_out(17), QN => n147);
   reg_reg_16_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n98, Q => 
                           data_out(16), QN => n148);
   reg_reg_15_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n98, Q => 
                           data_out(15), QN => n149);
   reg_reg_14_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n98, Q => 
                           data_out(14), QN => n150);
   reg_reg_13_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n98, Q => 
                           data_out(13), QN => n151);
   reg_reg_12_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n98, Q => 
                           data_out(12), QN => n152);
   reg_reg_11_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n98, Q => 
                           data_out(11), QN => n153);
   reg_reg_10_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n98, Q => 
                           data_out(10), QN => n154);
   reg_reg_9_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n99, Q => 
                           data_out(9), QN => n155);
   reg_reg_8_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n99, Q => 
                           data_out(8), QN => n156);
   reg_reg_7_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n99, Q => 
                           data_out(7), QN => n157);
   reg_reg_6_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n99, Q => 
                           data_out(6), QN => n158);
   reg_reg_5_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n99, Q => 
                           data_out(5), QN => n159);
   reg_reg_4_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n99, Q => 
                           data_out(4), QN => n160);
   reg_reg_3_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n99, Q => 
                           data_out(3), QN => n161);
   reg_reg_2_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n99, Q => 
                           data_out(2), QN => n162);
   reg_reg_1_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n99, Q => 
                           data_out(1), QN => n163);
   reg_reg_0_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n99, Q => 
                           data_out(0), QN => n164);
   U2 : BUF_X1 port map( A => n100, Z => n98);
   U3 : BUF_X1 port map( A => n100, Z => n96);
   U4 : BUF_X1 port map( A => n100, Z => n99);
   U5 : OAI21_X1 port map( B1 => n145, B2 => enable, A => n177, ZN => n113);
   U6 : NAND2_X1 port map( A1 => data_in(19), A2 => enable, ZN => n177);
   U7 : OAI21_X1 port map( B1 => n157, B2 => enable, A => n189, ZN => n125);
   U8 : NAND2_X1 port map( A1 => data_in(7), A2 => enable, ZN => n189);
   U9 : OAI21_X1 port map( B1 => n153, B2 => enable, A => n185, ZN => n121);
   U10 : NAND2_X1 port map( A1 => data_in(11), A2 => enable, ZN => n185);
   U11 : OAI21_X1 port map( B1 => n148, B2 => enable, A => n180, ZN => n116);
   U12 : NAND2_X1 port map( A1 => data_in(16), A2 => enable, ZN => n180);
   U13 : OAI21_X1 port map( B1 => n147, B2 => enable, A => n179, ZN => n115);
   U14 : NAND2_X1 port map( A1 => data_in(17), A2 => enable, ZN => n179);
   U15 : OAI21_X1 port map( B1 => n146, B2 => enable, A => n178, ZN => n114);
   U16 : NAND2_X1 port map( A1 => data_in(18), A2 => enable, ZN => n178);
   U17 : OAI21_X1 port map( B1 => n160, B2 => enable, A => n192, ZN => n128);
   U18 : NAND2_X1 port map( A1 => data_in(4), A2 => enable, ZN => n192);
   U19 : OAI21_X1 port map( B1 => n159, B2 => enable, A => n191, ZN => n127);
   U20 : NAND2_X1 port map( A1 => data_in(5), A2 => enable, ZN => n191);
   U21 : OAI21_X1 port map( B1 => n158, B2 => enable, A => n190, ZN => n126);
   U22 : NAND2_X1 port map( A1 => data_in(6), A2 => enable, ZN => n190);
   U23 : OAI21_X1 port map( B1 => n156, B2 => enable, A => n188, ZN => n124);
   U24 : NAND2_X1 port map( A1 => data_in(8), A2 => enable, ZN => n188);
   U25 : OAI21_X1 port map( B1 => n155, B2 => enable, A => n187, ZN => n123);
   U26 : NAND2_X1 port map( A1 => data_in(9), A2 => enable, ZN => n187);
   U27 : OAI21_X1 port map( B1 => n154, B2 => enable, A => n186, ZN => n122);
   U28 : NAND2_X1 port map( A1 => data_in(10), A2 => enable, ZN => n186);
   U29 : OAI21_X1 port map( B1 => n152, B2 => enable, A => n184, ZN => n120);
   U30 : NAND2_X1 port map( A1 => data_in(12), A2 => enable, ZN => n184);
   U31 : OAI21_X1 port map( B1 => n151, B2 => enable, A => n183, ZN => n119);
   U32 : NAND2_X1 port map( A1 => data_in(13), A2 => enable, ZN => n183);
   U33 : OAI21_X1 port map( B1 => n150, B2 => enable, A => n182, ZN => n118);
   U34 : NAND2_X1 port map( A1 => data_in(14), A2 => enable, ZN => n182);
   U35 : OAI21_X1 port map( B1 => n149, B2 => enable, A => n181, ZN => n117);
   U36 : NAND2_X1 port map( A1 => data_in(15), A2 => enable, ZN => n181);
   U37 : OAI21_X1 port map( B1 => n144, B2 => enable, A => n176, ZN => n112);
   U38 : NAND2_X1 port map( A1 => data_in(20), A2 => enable, ZN => n176);
   U39 : OAI21_X1 port map( B1 => n143, B2 => enable, A => n175, ZN => n111);
   U40 : NAND2_X1 port map( A1 => data_in(21), A2 => enable, ZN => n175);
   U41 : OAI21_X1 port map( B1 => n142, B2 => enable, A => n174, ZN => n110);
   U42 : NAND2_X1 port map( A1 => data_in(22), A2 => enable, ZN => n174);
   U43 : OAI21_X1 port map( B1 => n141, B2 => enable, A => n173, ZN => n109);
   U44 : NAND2_X1 port map( A1 => data_in(23), A2 => enable, ZN => n173);
   U45 : OAI21_X1 port map( B1 => n140, B2 => enable, A => n172, ZN => n108);
   U46 : NAND2_X1 port map( A1 => data_in(24), A2 => enable, ZN => n172);
   U47 : OAI21_X1 port map( B1 => n139, B2 => enable, A => n171, ZN => n107);
   U48 : NAND2_X1 port map( A1 => data_in(25), A2 => enable, ZN => n171);
   U49 : OAI21_X1 port map( B1 => n138, B2 => enable, A => n170, ZN => n106);
   U50 : NAND2_X1 port map( A1 => data_in(26), A2 => enable, ZN => n170);
   U51 : OAI21_X1 port map( B1 => n137, B2 => enable, A => n169, ZN => n105);
   U52 : NAND2_X1 port map( A1 => data_in(27), A2 => enable, ZN => n169);
   U53 : OAI21_X1 port map( B1 => n136, B2 => enable, A => n168, ZN => n104);
   U54 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n168);
   U55 : OAI21_X1 port map( B1 => n135, B2 => enable, A => n167, ZN => n103);
   U56 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n167);
   U57 : OAI21_X1 port map( B1 => n134, B2 => enable, A => n166, ZN => n102);
   U58 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n166);
   U59 : OAI21_X1 port map( B1 => n133, B2 => enable, A => n165, ZN => n101);
   U60 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n165);
   U61 : OAI21_X1 port map( B1 => n163, B2 => enable, A => n195, ZN => n131);
   U62 : NAND2_X1 port map( A1 => data_in(1), A2 => enable, ZN => n195);
   U63 : OAI21_X1 port map( B1 => n162, B2 => enable, A => n194, ZN => n130);
   U64 : NAND2_X1 port map( A1 => data_in(2), A2 => enable, ZN => n194);
   U65 : OAI21_X1 port map( B1 => n161, B2 => enable, A => n193, ZN => n129);
   U66 : NAND2_X1 port map( A1 => data_in(3), A2 => enable, ZN => n193);
   U67 : OAI21_X1 port map( B1 => n164, B2 => enable, A => n196, ZN => n132);
   U68 : NAND2_X1 port map( A1 => enable, A2 => data_in(0), ZN => n196);
   U69 : INV_X1 port map( A => reset, ZN => n100);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_2 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_2;

architecture SYN_Behavioral of REG_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198 : std_logic;

begin
   
   reg_reg_19_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n99, Q => 
                           data_out(19), QN => n147);
   reg_reg_18_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n99, Q => 
                           data_out(18), QN => n148);
   reg_reg_17_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n99, Q => 
                           data_out(17), QN => n149);
   reg_reg_16_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n99, Q => 
                           data_out(16), QN => n150);
   reg_reg_15_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n99, Q => 
                           data_out(15), QN => n151);
   reg_reg_14_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n99, Q => 
                           data_out(14), QN => n152);
   reg_reg_13_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n99, Q => 
                           data_out(13), QN => n153);
   reg_reg_12_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n99, Q => 
                           data_out(12), QN => n154);
   reg_reg_11_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n99, Q => 
                           data_out(11), QN => n155);
   reg_reg_10_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n99, Q => 
                           data_out(10), QN => n156);
   reg_reg_9_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n100, Q => 
                           data_out(9), QN => n157);
   reg_reg_8_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n100, Q => 
                           data_out(8), QN => n158);
   reg_reg_6_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n100, Q => 
                           data_out(6), QN => n160);
   reg_reg_5_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n100, Q => 
                           data_out(5), QN => n161);
   reg_reg_4_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n100, Q => 
                           data_out(4), QN => n162);
   reg_reg_3_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n100, Q => 
                           data_out(3), QN => n163);
   reg_reg_2_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n100, Q => 
                           data_out(2), QN => n164);
   reg_reg_1_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n100, Q => 
                           data_out(1), QN => n165);
   reg_reg_0_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n100, Q => 
                           data_out(0), QN => n166);
   reg_reg_7_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n102, Q => 
                           data_out(7), QN => n159);
   reg_reg_22_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n102, Q => 
                           data_out(22), QN => n144);
   reg_reg_21_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n102, Q => 
                           data_out(21), QN => n145);
   reg_reg_20_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n102, Q => 
                           data_out(20), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n102, Q => 
                           data_out(26), QN => n140);
   reg_reg_25_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n102, Q => 
                           data_out(25), QN => n141);
   reg_reg_24_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n102, Q => 
                           data_out(24), QN => n142);
   reg_reg_23_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n102, Q => 
                           data_out(23), QN => n143);
   reg_reg_27_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n102, Q => 
                           data_out(27), QN => n139);
   reg_reg_31_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n102, Q => 
                           data_out(31), QN => n135);
   reg_reg_30_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n102, Q => 
                           data_out(30), QN => n136);
   reg_reg_29_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n102, Q => 
                           data_out(29), QN => n137);
   reg_reg_28_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n102, Q => 
                           data_out(28), QN => n138);
   U2 : OR2_X2 port map( A1 => n138, A2 => enable, ZN => n96);
   U3 : NAND2_X1 port map( A1 => n96, A2 => n170, ZN => n106);
   U4 : OR2_X1 port map( A1 => n135, A2 => enable, ZN => n98);
   U5 : NAND2_X1 port map( A1 => n98, A2 => n167, ZN => n103);
   U6 : BUF_X1 port map( A => n102, Z => n101);
   U7 : BUF_X1 port map( A => n101, Z => n100);
   U8 : BUF_X1 port map( A => n101, Z => n99);
   U9 : OAI21_X1 port map( B1 => n143, B2 => enable, A => n175, ZN => n111);
   U10 : NAND2_X1 port map( A1 => data_in(23), A2 => enable, ZN => n175);
   U11 : OAI21_X1 port map( B1 => n146, B2 => enable, A => n178, ZN => n114);
   U12 : NAND2_X1 port map( A1 => data_in(20), A2 => enable, ZN => n178);
   U13 : OAI21_X1 port map( B1 => n145, B2 => enable, A => n177, ZN => n113);
   U14 : NAND2_X1 port map( A1 => data_in(21), A2 => enable, ZN => n177);
   U15 : OAI21_X1 port map( B1 => n144, B2 => enable, A => n176, ZN => n112);
   U16 : NAND2_X1 port map( A1 => data_in(22), A2 => enable, ZN => n176);
   U17 : OAI21_X1 port map( B1 => n139, B2 => enable, A => n171, ZN => n107);
   U18 : NAND2_X1 port map( A1 => data_in(27), A2 => enable, ZN => n171);
   U19 : OAI21_X1 port map( B1 => n142, B2 => enable, A => n174, ZN => n110);
   U20 : NAND2_X1 port map( A1 => data_in(24), A2 => enable, ZN => n174);
   U21 : OAI21_X1 port map( B1 => n141, B2 => enable, A => n173, ZN => n109);
   U22 : NAND2_X1 port map( A1 => data_in(25), A2 => enable, ZN => n173);
   U23 : OAI21_X1 port map( B1 => n140, B2 => enable, A => n172, ZN => n108);
   U24 : NAND2_X1 port map( A1 => data_in(26), A2 => enable, ZN => n172);
   U25 : OAI21_X1 port map( B1 => n137, B2 => enable, A => n169, ZN => n105);
   U26 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n169);
   U27 : OAI21_X1 port map( B1 => n136, B2 => enable, A => n168, ZN => n104);
   U28 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n168);
   U29 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n170);
   U30 : OAI21_X1 port map( B1 => n147, B2 => enable, A => n179, ZN => n115);
   U31 : NAND2_X1 port map( A1 => data_in(19), A2 => enable, ZN => n179);
   U32 : OAI21_X1 port map( B1 => n150, B2 => enable, A => n182, ZN => n118);
   U33 : NAND2_X1 port map( A1 => data_in(16), A2 => enable, ZN => n182);
   U34 : OAI21_X1 port map( B1 => n149, B2 => enable, A => n181, ZN => n117);
   U35 : NAND2_X1 port map( A1 => data_in(17), A2 => enable, ZN => n181);
   U36 : OAI21_X1 port map( B1 => n148, B2 => enable, A => n180, ZN => n116);
   U37 : NAND2_X1 port map( A1 => data_in(18), A2 => enable, ZN => n180);
   U38 : OAI21_X1 port map( B1 => n151, B2 => enable, A => n183, ZN => n119);
   U39 : NAND2_X1 port map( A1 => data_in(15), A2 => enable, ZN => n183);
   U40 : OAI21_X1 port map( B1 => n154, B2 => enable, A => n186, ZN => n122);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => enable, ZN => n186);
   U42 : OAI21_X1 port map( B1 => n153, B2 => enable, A => n185, ZN => n121);
   U43 : NAND2_X1 port map( A1 => data_in(13), A2 => enable, ZN => n185);
   U44 : OAI21_X1 port map( B1 => n152, B2 => enable, A => n184, ZN => n120);
   U45 : NAND2_X1 port map( A1 => data_in(14), A2 => enable, ZN => n184);
   U46 : OAI21_X1 port map( B1 => n155, B2 => enable, A => n187, ZN => n123);
   U47 : NAND2_X1 port map( A1 => data_in(11), A2 => enable, ZN => n187);
   U48 : OAI21_X1 port map( B1 => n158, B2 => enable, A => n190, ZN => n126);
   U49 : NAND2_X1 port map( A1 => data_in(8), A2 => enable, ZN => n190);
   U50 : OAI21_X1 port map( B1 => n157, B2 => enable, A => n189, ZN => n125);
   U51 : NAND2_X1 port map( A1 => data_in(9), A2 => enable, ZN => n189);
   U52 : OAI21_X1 port map( B1 => n156, B2 => enable, A => n188, ZN => n124);
   U53 : NAND2_X1 port map( A1 => data_in(10), A2 => enable, ZN => n188);
   U54 : OAI21_X1 port map( B1 => n159, B2 => enable, A => n191, ZN => n127);
   U55 : NAND2_X1 port map( A1 => data_in(7), A2 => enable, ZN => n191);
   U56 : OAI21_X1 port map( B1 => n162, B2 => enable, A => n194, ZN => n130);
   U57 : NAND2_X1 port map( A1 => data_in(4), A2 => enable, ZN => n194);
   U58 : OAI21_X1 port map( B1 => n161, B2 => enable, A => n193, ZN => n129);
   U59 : NAND2_X1 port map( A1 => data_in(5), A2 => enable, ZN => n193);
   U60 : OAI21_X1 port map( B1 => n160, B2 => enable, A => n192, ZN => n128);
   U61 : NAND2_X1 port map( A1 => data_in(6), A2 => enable, ZN => n192);
   U62 : OAI21_X1 port map( B1 => n163, B2 => enable, A => n195, ZN => n131);
   U63 : NAND2_X1 port map( A1 => data_in(3), A2 => enable, ZN => n195);
   U64 : OAI21_X1 port map( B1 => n164, B2 => enable, A => n196, ZN => n132);
   U65 : NAND2_X1 port map( A1 => data_in(2), A2 => enable, ZN => n196);
   U66 : OAI21_X1 port map( B1 => n165, B2 => enable, A => n197, ZN => n133);
   U67 : NAND2_X1 port map( A1 => data_in(1), A2 => enable, ZN => n197);
   U68 : OAI21_X1 port map( B1 => n166, B2 => enable, A => n198, ZN => n134);
   U69 : NAND2_X1 port map( A1 => enable, A2 => data_in(0), ZN => n198);
   U70 : INV_X1 port map( A => reset, ZN => n102);
   U71 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n167);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_1 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_1;

architecture SYN_Behavioral of REG_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n96, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198 : std_logic;

begin
   
   reg_reg_19_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n99, Q => 
                           data_out(19), QN => n147);
   reg_reg_18_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n99, Q => 
                           data_out(18), QN => n148);
   reg_reg_17_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n99, Q => 
                           data_out(17), QN => n149);
   reg_reg_16_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n99, Q => 
                           data_out(16), QN => n150);
   reg_reg_15_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n99, Q => 
                           data_out(15), QN => n151);
   reg_reg_14_inst : DFFR_X1 port map( D => n120, CK => clk, RN => n99, Q => 
                           data_out(14), QN => n152);
   reg_reg_13_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n99, Q => 
                           data_out(13), QN => n153);
   reg_reg_12_inst : DFFR_X1 port map( D => n122, CK => clk, RN => n99, Q => 
                           data_out(12), QN => n154);
   reg_reg_11_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n99, Q => 
                           data_out(11), QN => n155);
   reg_reg_10_inst : DFFR_X1 port map( D => n124, CK => clk, RN => n99, Q => 
                           data_out(10), QN => n156);
   reg_reg_9_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n100, Q => 
                           data_out(9), QN => n157);
   reg_reg_8_inst : DFFR_X1 port map( D => n126, CK => clk, RN => n100, Q => 
                           data_out(8), QN => n158);
   reg_reg_7_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n100, Q => 
                           data_out(7), QN => n159);
   reg_reg_6_inst : DFFR_X1 port map( D => n128, CK => clk, RN => n100, Q => 
                           data_out(6), QN => n160);
   reg_reg_5_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n100, Q => 
                           data_out(5), QN => n161);
   reg_reg_4_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n100, Q => 
                           data_out(4), QN => n162);
   reg_reg_3_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n100, Q => 
                           data_out(3), QN => n163);
   reg_reg_2_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n100, Q => 
                           data_out(2), QN => n164);
   reg_reg_1_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n100, Q => 
                           data_out(1), QN => n165);
   reg_reg_0_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n100, Q => 
                           data_out(0), QN => n166);
   reg_reg_22_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n102, Q => 
                           data_out(22), QN => n144);
   reg_reg_21_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n102, Q => 
                           data_out(21), QN => n145);
   reg_reg_20_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n102, Q => 
                           data_out(20), QN => n146);
   reg_reg_26_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n102, Q => 
                           data_out(26), QN => n140);
   reg_reg_25_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n102, Q => 
                           data_out(25), QN => n141);
   reg_reg_24_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n102, Q => 
                           data_out(24), QN => n142);
   reg_reg_23_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n102, Q => 
                           data_out(23), QN => n143);
   reg_reg_27_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n102, Q => 
                           data_out(27), QN => n139);
   reg_reg_31_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n102, Q => 
                           data_out(31), QN => n135);
   reg_reg_29_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n102, Q => 
                           data_out(29), QN => n137);
   reg_reg_28_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n102, Q => 
                           data_out(28), QN => n138);
   reg_reg_30_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n102, Q => 
                           data_out(30), QN => n136);
   U2 : OR2_X1 port map( A1 => n136, A2 => enable, ZN => n96);
   U3 : NAND2_X1 port map( A1 => n96, A2 => n168, ZN => n104);
   U4 : OR2_X1 port map( A1 => n135, A2 => enable, ZN => n98);
   U5 : NAND2_X1 port map( A1 => n167, A2 => n98, ZN => n103);
   U6 : BUF_X1 port map( A => n102, Z => n101);
   U7 : BUF_X1 port map( A => n101, Z => n99);
   U8 : BUF_X1 port map( A => n101, Z => n100);
   U9 : OAI21_X1 port map( B1 => n138, B2 => enable, A => n170, ZN => n106);
   U10 : NAND2_X1 port map( A1 => data_in(28), A2 => enable, ZN => n170);
   U11 : OAI21_X1 port map( B1 => n137, B2 => enable, A => n169, ZN => n105);
   U12 : NAND2_X1 port map( A1 => data_in(29), A2 => enable, ZN => n169);
   U13 : NAND2_X1 port map( A1 => data_in(30), A2 => enable, ZN => n168);
   U14 : NAND2_X1 port map( A1 => data_in(31), A2 => enable, ZN => n167);
   U15 : OAI21_X1 port map( B1 => n143, B2 => enable, A => n175, ZN => n111);
   U16 : NAND2_X1 port map( A1 => data_in(23), A2 => enable, ZN => n175);
   U17 : OAI21_X1 port map( B1 => n139, B2 => enable, A => n171, ZN => n107);
   U18 : NAND2_X1 port map( A1 => data_in(27), A2 => enable, ZN => n171);
   U19 : OAI21_X1 port map( B1 => n142, B2 => enable, A => n174, ZN => n110);
   U20 : NAND2_X1 port map( A1 => data_in(24), A2 => enable, ZN => n174);
   U21 : OAI21_X1 port map( B1 => n141, B2 => enable, A => n173, ZN => n109);
   U22 : NAND2_X1 port map( A1 => data_in(25), A2 => enable, ZN => n173);
   U23 : OAI21_X1 port map( B1 => n140, B2 => enable, A => n172, ZN => n108);
   U24 : NAND2_X1 port map( A1 => data_in(26), A2 => enable, ZN => n172);
   U25 : OAI21_X1 port map( B1 => n146, B2 => enable, A => n178, ZN => n114);
   U26 : NAND2_X1 port map( A1 => data_in(20), A2 => enable, ZN => n178);
   U27 : OAI21_X1 port map( B1 => n145, B2 => enable, A => n177, ZN => n113);
   U28 : NAND2_X1 port map( A1 => data_in(21), A2 => enable, ZN => n177);
   U29 : OAI21_X1 port map( B1 => n144, B2 => enable, A => n176, ZN => n112);
   U30 : NAND2_X1 port map( A1 => data_in(22), A2 => enable, ZN => n176);
   U31 : OAI21_X1 port map( B1 => n147, B2 => enable, A => n179, ZN => n115);
   U32 : NAND2_X1 port map( A1 => data_in(19), A2 => enable, ZN => n179);
   U33 : OAI21_X1 port map( B1 => n150, B2 => enable, A => n182, ZN => n118);
   U34 : NAND2_X1 port map( A1 => data_in(16), A2 => enable, ZN => n182);
   U35 : OAI21_X1 port map( B1 => n149, B2 => enable, A => n181, ZN => n117);
   U36 : NAND2_X1 port map( A1 => data_in(17), A2 => enable, ZN => n181);
   U37 : OAI21_X1 port map( B1 => n148, B2 => enable, A => n180, ZN => n116);
   U38 : NAND2_X1 port map( A1 => data_in(18), A2 => enable, ZN => n180);
   U39 : OAI21_X1 port map( B1 => n151, B2 => enable, A => n183, ZN => n119);
   U40 : NAND2_X1 port map( A1 => data_in(15), A2 => enable, ZN => n183);
   U41 : OAI21_X1 port map( B1 => n154, B2 => enable, A => n186, ZN => n122);
   U42 : NAND2_X1 port map( A1 => data_in(12), A2 => enable, ZN => n186);
   U43 : OAI21_X1 port map( B1 => n153, B2 => enable, A => n185, ZN => n121);
   U44 : NAND2_X1 port map( A1 => data_in(13), A2 => enable, ZN => n185);
   U45 : OAI21_X1 port map( B1 => n152, B2 => enable, A => n184, ZN => n120);
   U46 : NAND2_X1 port map( A1 => data_in(14), A2 => enable, ZN => n184);
   U47 : OAI21_X1 port map( B1 => n155, B2 => enable, A => n187, ZN => n123);
   U48 : NAND2_X1 port map( A1 => data_in(11), A2 => enable, ZN => n187);
   U49 : OAI21_X1 port map( B1 => n158, B2 => enable, A => n190, ZN => n126);
   U50 : NAND2_X1 port map( A1 => data_in(8), A2 => enable, ZN => n190);
   U51 : OAI21_X1 port map( B1 => n157, B2 => enable, A => n189, ZN => n125);
   U52 : NAND2_X1 port map( A1 => data_in(9), A2 => enable, ZN => n189);
   U53 : OAI21_X1 port map( B1 => n156, B2 => enable, A => n188, ZN => n124);
   U54 : NAND2_X1 port map( A1 => data_in(10), A2 => enable, ZN => n188);
   U55 : OAI21_X1 port map( B1 => n159, B2 => enable, A => n191, ZN => n127);
   U56 : NAND2_X1 port map( A1 => data_in(7), A2 => enable, ZN => n191);
   U57 : OAI21_X1 port map( B1 => n162, B2 => enable, A => n194, ZN => n130);
   U58 : NAND2_X1 port map( A1 => data_in(4), A2 => enable, ZN => n194);
   U59 : OAI21_X1 port map( B1 => n161, B2 => enable, A => n193, ZN => n129);
   U60 : NAND2_X1 port map( A1 => data_in(5), A2 => enable, ZN => n193);
   U61 : OAI21_X1 port map( B1 => n160, B2 => enable, A => n192, ZN => n128);
   U62 : NAND2_X1 port map( A1 => data_in(6), A2 => enable, ZN => n192);
   U63 : OAI21_X1 port map( B1 => n163, B2 => enable, A => n195, ZN => n131);
   U64 : NAND2_X1 port map( A1 => data_in(3), A2 => enable, ZN => n195);
   U65 : OAI21_X1 port map( B1 => n164, B2 => enable, A => n196, ZN => n132);
   U66 : NAND2_X1 port map( A1 => data_in(2), A2 => enable, ZN => n196);
   U67 : OAI21_X1 port map( B1 => n165, B2 => enable, A => n197, ZN => n133);
   U68 : NAND2_X1 port map( A1 => data_in(1), A2 => enable, ZN => n197);
   U69 : OAI21_X1 port map( B1 => n166, B2 => enable, A => n198, ZN => n134);
   U70 : NAND2_X1 port map( A1 => enable, A2 => data_in(0), ZN => n198);
   U71 : INV_X1 port map( A => reset, ZN => n102);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX2to1_NBIT4_0;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => Y(3));
   U2 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U3 : INV_X1 port map( A => n7, ZN => Y(2));
   U4 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U5 : INV_X1 port map( A => n8, ZN => Y(1));
   U6 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U7 : INV_X1 port map( A => n9, ZN => Y(0));
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCAN_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCAN_NBIT4_0;

architecture SYN_BEHAVIORAL of RCAN_NBIT4_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_49_2_carry_1_port, add_1_root_add_49_2_carry_2_port, 
      add_1_root_add_49_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_49_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_49_2_carry_1_port, S => S(0));
   add_1_root_add_49_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_49_2_carry_1_port, CO => 
                           add_1_root_add_49_2_carry_2_port, S => S(1));
   add_1_root_add_49_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_49_2_carry_2_port, CO => 
                           add_1_root_add_49_2_carry_3_port, S => S(2));
   add_1_root_add_49_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_49_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_SEL_N_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CARRY_SEL_N_NBIT4_0;

architecture SYN_STRUCTURAL of CARRY_SEL_N_NBIT4_0 is

   component MUX2to1_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCAN_NBIT4_127
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCAN_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S0_3_port, S0_2_port, S0_1_port, S0_0_port, n_1168, n_1169 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCAN_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1168);
   RCA0 : RCAN_NBIT4_127 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1169);
   MUX21 : MUX2to1_NBIT4_0 port map( A(3) => S0_3_port, A(2) => S0_2_port, A(1)
                           => S0_1_port, A(0) => S0_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_block_0 is

   port( A, B : in std_logic_vector (1 downto 0);  PGout : out std_logic_vector
         (1 downto 0));

end PG_block_0;

architecture SYN_BEHAVIORAL of PG_block_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => PGout(1));
   U2 : INV_X1 port map( A => n2, ZN => PGout(0));
   U3 : AOI21_X1 port map( B1 => B(0), B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity G_block_0 is

   port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : out 
         std_logic);

end G_block_0;

architecture SYN_BEHAVIORAL of G_block_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gout);
   U2 : AOI21_X1 port map( B1 => B, B2 => A(1), A => A(0), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_network_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
         std_logic_vector (31 downto 0));

end PG_network_NBIT32_0;

architecture SYN_BEHAVIORAL of PG_network_NBIT32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U33 : XOR2_X1 port map( A => B(9), B => A(9), Z => Pout(9));
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => Pout(8));
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => Pout(7));
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => Pout(6));
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => Pout(5));
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => Pout(4));
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => Pout(3));
   U40 : XOR2_X1 port map( A => B(31), B => A(31), Z => Pout(31));
   U41 : XOR2_X1 port map( A => B(30), B => A(30), Z => Pout(30));
   U42 : XOR2_X1 port map( A => B(2), B => A(2), Z => Pout(2));
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => Pout(29));
   U44 : XOR2_X1 port map( A => B(28), B => A(28), Z => Pout(28));
   U45 : XOR2_X1 port map( A => B(27), B => A(27), Z => Pout(27));
   U46 : XOR2_X1 port map( A => B(26), B => A(26), Z => Pout(26));
   U47 : XOR2_X1 port map( A => B(25), B => A(25), Z => Pout(25));
   U48 : XOR2_X1 port map( A => B(24), B => A(24), Z => Pout(24));
   U49 : XOR2_X1 port map( A => B(23), B => A(23), Z => Pout(23));
   U50 : XOR2_X1 port map( A => B(22), B => A(22), Z => Pout(22));
   U51 : XOR2_X1 port map( A => B(21), B => A(21), Z => Pout(21));
   U52 : XOR2_X1 port map( A => B(20), B => A(20), Z => Pout(20));
   U53 : XOR2_X1 port map( A => B(1), B => A(1), Z => Pout(1));
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => Pout(19));
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => Pout(18));
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => Pout(17));
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => Pout(16));
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => Pout(15));
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => Pout(14));
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => Pout(13));
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => Pout(12));
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => Pout(11));
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => Pout(10));
   U64 : XOR2_X1 port map( A => B(0), B => A(0), Z => Pout(0));
   U1 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Gout(1));
   U2 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Gout(18));
   U3 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Gout(4));
   U4 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Gout(21));
   U5 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Gout(20));
   U6 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Gout(22));
   U7 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Gout(17));
   U8 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Gout(16));
   U9 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Gout(10));
   U10 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Gout(11));
   U11 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Gout(8));
   U12 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Gout(14));
   U13 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Gout(13));
   U14 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Gout(12));
   U15 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Gout(6));
   U16 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Gout(26));
   U17 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Gout(27));
   U18 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Gout(25));
   U19 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Gout(24));
   U20 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Gout(31));
   U21 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Gout(30));
   U22 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Gout(28));
   U23 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Gout(29));
   U24 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Gout(19));
   U25 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Gout(2));
   U26 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Gout(23));
   U27 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Gout(9));
   U28 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Gout(5));
   U29 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Gout(3));
   U30 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Gout(15));
   U31 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Gout(7));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Gout(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_0 is

   port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
         std_logic_vector (2 downto 0));

end ENCODER_0;

architecture SYN_BEHAVIORAL of ENCODER_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n1, n2 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => INPUT(0), B => INPUT(1), Z => n4);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n3, A3 => n4, ZN => OUTPUT(2));
   U2 : OAI21_X1 port map( B1 => INPUT(2), B2 => n2, A => n5, ZN => OUTPUT(0));
   U3 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n5, ZN => OUTPUT(1));
   U4 : INV_X1 port map( A => INPUT(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => n5);
   U6 : INV_X1 port map( A => n4, ZN => n2);
   U7 : AND2_X1 port map( A1 => INPUT(1), A2 => INPUT(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND4_0 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end ND4_0;

architecture SYN_ARCH1 of ND4_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ND3_0 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end ND3_0;

architecture SYN_ARCH1 of ND3_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0;

architecture SYN_STRUCTURAL of SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 is

   component CARRY_SEL_N_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SEL_N_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   UCSi_1 : CARRY_SEL_N_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   UCSi_2 : CARRY_SEL_N_NBIT4_63 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   UCSi_3 : CARRY_SEL_N_NBIT4_62 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   UCSi_4 : CARRY_SEL_N_NBIT4_61 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   UCSi_5 : CARRY_SEL_N_NBIT4_60 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   UCSi_6 : CARRY_SEL_N_NBIT4_59 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   UCSi_7 : CARRY_SEL_N_NBIT4_58 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   UCSi_8 : CARRY_SEL_N_NBIT4_57 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_block_64
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_65
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_66
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_67
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_190
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_191
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_68
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component G_block_69
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_192
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_193
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_194
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_70
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_195
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_196
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_197
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_198
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_199
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_200
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_201
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_71
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_block_202
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_203
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_204
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_205
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_206
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_207
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_208
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_209
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_210
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_211
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_212
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_213
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_214
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_215
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_block_0
      port( A, B : in std_logic_vector (1 downto 0);  PGout : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_block_0
      port( A : in std_logic_vector (1 downto 0);  B : in std_logic;  Gout : 
            out std_logic);
   end component;
   
   component PG_network_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  Pout, Gout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, G_1_0_port, G_16_16_port, G_16_15_port, 
      G_16_13_port, G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, 
      G_10_10_port, G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port
      , G_7_7_port, G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port,
      G_3_3_port, G_2_2_port, G_2_0_port, G_32_32_port, G_32_31_port, 
      G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, 
      G_30_29_port, G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, 
      G_28_17_port, G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, 
      G_24_24_port, G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, 
      G_22_22_port, G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, 
      G_20_17_port, G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, 
      P_16_16_port, P_16_15_port, P_16_13_port, P_16_9_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_12_port, P_12_11_port, 
      P_12_9_port, P_11_11_port, P_10_10_port, P_10_9_port, P_9_9_port, 
      P_8_8_port, P_8_7_port, P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, 
      P_5_5_port, P_4_4_port, P_4_3_port, P_3_3_port, P_2_2_port, P_32_32_port,
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, N2, n1, n2_port, n3, n4, n5, n_1170 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgnetwork_0 : PG_network_NBIT32_0 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Pout(31) => P_32_32_port, 
                           Pout(30) => P_31_31_port, Pout(29) => P_30_30_port, 
                           Pout(28) => P_29_29_port, Pout(27) => P_28_28_port, 
                           Pout(26) => P_27_27_port, Pout(25) => P_26_26_port, 
                           Pout(24) => P_25_25_port, Pout(23) => P_24_24_port, 
                           Pout(22) => P_23_23_port, Pout(21) => P_22_22_port, 
                           Pout(20) => P_21_21_port, Pout(19) => P_20_20_port, 
                           Pout(18) => P_19_19_port, Pout(17) => P_18_18_port, 
                           Pout(16) => P_17_17_port, Pout(15) => P_16_16_port, 
                           Pout(14) => P_15_15_port, Pout(13) => P_14_14_port, 
                           Pout(12) => P_13_13_port, Pout(11) => P_12_12_port, 
                           Pout(10) => P_11_11_port, Pout(9) => P_10_10_port, 
                           Pout(8) => P_9_9_port, Pout(7) => P_8_8_port, 
                           Pout(6) => P_7_7_port, Pout(5) => P_6_6_port, 
                           Pout(4) => P_5_5_port, Pout(3) => P_4_4_port, 
                           Pout(2) => P_3_3_port, Pout(1) => P_2_2_port, 
                           Pout(0) => n_1170, Gout(31) => G_32_32_port, 
                           Gout(30) => G_31_31_port, Gout(29) => G_30_30_port, 
                           Gout(28) => G_29_29_port, Gout(27) => G_28_28_port, 
                           Gout(26) => G_27_27_port, Gout(25) => G_26_26_port, 
                           Gout(24) => G_25_25_port, Gout(23) => G_24_24_port, 
                           Gout(22) => G_23_23_port, Gout(21) => G_22_22_port, 
                           Gout(20) => G_21_21_port, Gout(19) => G_20_20_port, 
                           Gout(18) => G_19_19_port, Gout(17) => G_18_18_port, 
                           Gout(16) => G_17_17_port, Gout(15) => G_16_16_port, 
                           Gout(14) => G_15_15_port, Gout(13) => G_14_14_port, 
                           Gout(12) => G_13_13_port, Gout(11) => G_12_12_port, 
                           Gout(10) => G_11_11_port, Gout(9) => G_10_10_port, 
                           Gout(8) => G_9_9_port, Gout(7) => G_8_8_port, 
                           Gout(6) => G_7_7_port, Gout(5) => G_6_6_port, 
                           Gout(4) => G_5_5_port, Gout(3) => G_4_4_port, 
                           Gout(2) => G_3_3_port, Gout(1) => G_2_2_port, 
                           Gout(0) => n5);
   gblock1_1_1 : G_block_0 port map( A(1) => P_2_2_port, A(0) => G_2_2_port, B 
                           => G_1_0_port, Gout => G_2_0_port);
   pgblock1_1_2 : PG_block_0 port map( A(1) => P_4_4_port, A(0) => G_4_4_port, 
                           B(1) => P_3_3_port, B(0) => G_3_3_port, PGout(1) => 
                           P_4_3_port, PGout(0) => G_4_3_port);
   pgblock1_1_3 : PG_block_215 port map( A(1) => P_6_6_port, A(0) => G_6_6_port
                           , B(1) => P_5_5_port, B(0) => G_5_5_port, PGout(1) 
                           => P_6_5_port, PGout(0) => G_6_5_port);
   pgblock1_1_4 : PG_block_214 port map( A(1) => P_8_8_port, A(0) => G_8_8_port
                           , B(1) => P_7_7_port, B(0) => G_7_7_port, PGout(1) 
                           => P_8_7_port, PGout(0) => G_8_7_port);
   pgblock1_1_5 : PG_block_213 port map( A(1) => P_10_10_port, A(0) => 
                           G_10_10_port, B(1) => P_9_9_port, B(0) => G_9_9_port
                           , PGout(1) => P_10_9_port, PGout(0) => G_10_9_port);
   pgblock1_1_6 : PG_block_212 port map( A(1) => P_12_12_port, A(0) => 
                           G_12_12_port, B(1) => P_11_11_port, B(0) => 
                           G_11_11_port, PGout(1) => P_12_11_port, PGout(0) => 
                           G_12_11_port);
   pgblock1_1_7 : PG_block_211 port map( A(1) => P_14_14_port, A(0) => 
                           G_14_14_port, B(1) => P_13_13_port, B(0) => 
                           G_13_13_port, PGout(1) => P_14_13_port, PGout(0) => 
                           G_14_13_port);
   pgblock1_1_8 : PG_block_210 port map( A(1) => P_16_16_port, A(0) => 
                           G_16_16_port, B(1) => P_15_15_port, B(0) => 
                           G_15_15_port, PGout(1) => P_16_15_port, PGout(0) => 
                           G_16_15_port);
   pgblock1_1_9 : PG_block_209 port map( A(1) => P_18_18_port, A(0) => 
                           G_18_18_port, B(1) => P_17_17_port, B(0) => 
                           G_17_17_port, PGout(1) => P_18_17_port, PGout(0) => 
                           G_18_17_port);
   pgblock1_1_10 : PG_block_208 port map( A(1) => P_20_20_port, A(0) => 
                           G_20_20_port, B(1) => P_19_19_port, B(0) => 
                           G_19_19_port, PGout(1) => P_20_19_port, PGout(0) => 
                           G_20_19_port);
   pgblock1_1_11 : PG_block_207 port map( A(1) => P_22_22_port, A(0) => 
                           G_22_22_port, B(1) => P_21_21_port, B(0) => 
                           G_21_21_port, PGout(1) => P_22_21_port, PGout(0) => 
                           G_22_21_port);
   pgblock1_1_12 : PG_block_206 port map( A(1) => P_24_24_port, A(0) => 
                           G_24_24_port, B(1) => P_23_23_port, B(0) => 
                           G_23_23_port, PGout(1) => P_24_23_port, PGout(0) => 
                           G_24_23_port);
   pgblock1_1_13 : PG_block_205 port map( A(1) => P_26_26_port, A(0) => 
                           G_26_26_port, B(1) => P_25_25_port, B(0) => 
                           G_25_25_port, PGout(1) => P_26_25_port, PGout(0) => 
                           G_26_25_port);
   pgblock1_1_14 : PG_block_204 port map( A(1) => P_28_28_port, A(0) => 
                           G_28_28_port, B(1) => P_27_27_port, B(0) => 
                           G_27_27_port, PGout(1) => P_28_27_port, PGout(0) => 
                           G_28_27_port);
   pgblock1_1_15 : PG_block_203 port map( A(1) => P_30_30_port, A(0) => 
                           G_30_30_port, B(1) => P_29_29_port, B(0) => 
                           G_29_29_port, PGout(1) => P_30_29_port, PGout(0) => 
                           G_30_29_port);
   pgblock1_1_16 : PG_block_202 port map( A(1) => P_32_32_port, A(0) => 
                           G_32_32_port, B(1) => P_31_31_port, B(0) => 
                           G_31_31_port, PGout(1) => P_32_31_port, PGout(0) => 
                           G_32_31_port);
   gblock1_2_1 : G_block_71 port map( A(1) => P_4_3_port, A(0) => G_4_3_port, B
                           => G_2_0_port, Gout => Co_1_port);
   pgblock1_2_2 : PG_block_201 port map( A(1) => P_8_7_port, A(0) => G_8_7_port
                           , B(1) => P_6_5_port, B(0) => G_6_5_port, PGout(1) 
                           => P_8_5_port, PGout(0) => G_8_5_port);
   pgblock1_2_3 : PG_block_200 port map( A(1) => P_12_11_port, A(0) => 
                           G_12_11_port, B(1) => P_10_9_port, B(0) => 
                           G_10_9_port, PGout(1) => P_12_9_port, PGout(0) => 
                           G_12_9_port);
   pgblock1_2_4 : PG_block_199 port map( A(1) => P_16_15_port, A(0) => 
                           G_16_15_port, B(1) => P_14_13_port, B(0) => 
                           G_14_13_port, PGout(1) => P_16_13_port, PGout(0) => 
                           G_16_13_port);
   pgblock1_2_5 : PG_block_198 port map( A(1) => P_20_19_port, A(0) => 
                           G_20_19_port, B(1) => P_18_17_port, B(0) => 
                           G_18_17_port, PGout(1) => P_20_17_port, PGout(0) => 
                           G_20_17_port);
   pgblock1_2_6 : PG_block_197 port map( A(1) => P_24_23_port, A(0) => 
                           G_24_23_port, B(1) => P_22_21_port, B(0) => 
                           G_22_21_port, PGout(1) => P_24_21_port, PGout(0) => 
                           G_24_21_port);
   pgblock1_2_7 : PG_block_196 port map( A(1) => P_28_27_port, A(0) => 
                           G_28_27_port, B(1) => P_26_25_port, B(0) => 
                           G_26_25_port, PGout(1) => P_28_25_port, PGout(0) => 
                           G_28_25_port);
   pgblock1_2_8 : PG_block_195 port map( A(1) => P_32_31_port, A(0) => 
                           G_32_31_port, B(1) => P_30_29_port, B(0) => 
                           G_30_29_port, PGout(1) => P_32_29_port, PGout(0) => 
                           G_32_29_port);
   gblock1_3_1 : G_block_70 port map( A(1) => P_8_5_port, A(0) => G_8_5_port, B
                           => Co_1_port, Gout => Co_2_port);
   pgblock1_3_2 : PG_block_194 port map( A(1) => P_16_13_port, A(0) => 
                           G_16_13_port, B(1) => P_12_9_port, B(0) => 
                           G_12_9_port, PGout(1) => P_16_9_port, PGout(0) => 
                           G_16_9_port);
   pgblock1_3_3 : PG_block_193 port map( A(1) => P_24_21_port, A(0) => 
                           G_24_21_port, B(1) => P_20_17_port, B(0) => 
                           G_20_17_port, PGout(1) => P_24_17_port, PGout(0) => 
                           G_24_17_port);
   pgblock1_3_4 : PG_block_192 port map( A(1) => P_32_29_port, A(0) => 
                           G_32_29_port, B(1) => P_28_25_port, B(0) => 
                           G_28_25_port, PGout(1) => P_32_25_port, PGout(0) => 
                           G_32_25_port);
   gblock2_4_3 : G_block_69 port map( A(1) => P_12_9_port, A(0) => G_12_9_port,
                           B => Co_2_port, Gout => Co_3_port);
   gblock2_4_4 : G_block_68 port map( A(1) => P_16_9_port, A(0) => G_16_9_port,
                           B => Co_2_port, Gout => Co_4_port);
   pgblock2_4_28_2 : PG_block_191 port map( A(1) => P_28_25_port, A(0) => 
                           G_28_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_28_17_port, PGout(0) => 
                           G_28_17_port);
   pgblock2_4_32_2 : PG_block_190 port map( A(1) => P_32_25_port, A(0) => 
                           G_32_25_port, B(1) => P_24_17_port, B(0) => 
                           G_24_17_port, PGout(1) => P_32_17_port, PGout(0) => 
                           G_32_17_port);
   gblock2_5_5 : G_block_67 port map( A(1) => P_20_17_port, A(0) => 
                           G_20_17_port, B => Co_4_port, Gout => Co_5_port);
   gblock2_5_6 : G_block_66 port map( A(1) => P_24_17_port, A(0) => 
                           G_24_17_port, B => Co_4_port, Gout => Co_6_port);
   gblock2_5_7 : G_block_65 port map( A(1) => P_28_17_port, A(0) => 
                           G_28_17_port, B => Co_4_port, Gout => Co_7_port);
   gblock2_5_8 : G_block_64 port map( A(1) => P_32_17_port, A(0) => 
                           G_32_17_port, B => Co_4_port, Gout => Co_8_port);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n2_port, ZN => n3);
   U2 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => n1);
   U3 : NAND2_X1 port map( A1 => n5, A2 => Cin, ZN => n2_port);
   U4 : OR2_X1 port map( A1 => n3, A2 => n4, ZN => G_1_0_port);
   U5 : AND2_X1 port map( A1 => n5, A2 => N2, ZN => n4);
   U6 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => N2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUL is

   port( CLOCK : in std_logic;  A, B : in std_logic_vector (15 downto 0);  Y : 
         out std_logic_vector (31 downto 0));

end MUL;

architecture SYN_BEHAVIORAL of MUL is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_1
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_4
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_2
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_5
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_6
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component REG_NBIT32_3
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_7
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component MUX5to1_NBIT32_1
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_2
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_3
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_4
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_5
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_6
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_7
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX5to1_NBIT32_8
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component ENCODER_1
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_2
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_3
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_4
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_5
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_6
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_7
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component ENCODER_0
      port( INPUT : in std_logic_vector (2 downto 0);  OUTPUT : out 
            std_logic_vector (2 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, A_neg_15_30_port, A_neg_15_29_port, 
      A_neg_15_28_port, A_neg_15_27_port, A_neg_15_26_port, A_neg_15_25_port, 
      A_neg_15_24_port, A_neg_15_23_port, A_neg_15_22_port, A_neg_15_21_port, 
      A_neg_15_20_port, A_neg_15_19_port, A_neg_15_18_port, A_neg_15_17_port, 
      A_neg_15_16_port, A_neg_14_29_port, A_neg_14_28_port, A_neg_14_27_port, 
      A_neg_14_26_port, A_neg_14_25_port, A_neg_14_24_port, A_neg_14_23_port, 
      A_neg_14_22_port, A_neg_14_21_port, A_neg_14_20_port, A_neg_14_19_port, 
      A_neg_14_18_port, A_neg_14_17_port, A_neg_14_16_port, A_neg_14_15_port, 
      A_neg_13_28_port, A_neg_13_27_port, A_neg_13_26_port, A_neg_13_25_port, 
      A_neg_13_24_port, A_neg_13_23_port, A_neg_13_22_port, A_neg_13_21_port, 
      A_neg_13_20_port, A_neg_13_19_port, A_neg_13_18_port, A_neg_13_17_port, 
      A_neg_13_16_port, A_neg_13_15_port, A_neg_13_14_port, A_neg_12_27_port, 
      A_neg_12_26_port, A_neg_12_25_port, A_neg_12_24_port, A_neg_12_23_port, 
      A_neg_12_22_port, A_neg_12_21_port, A_neg_12_20_port, A_neg_12_19_port, 
      A_neg_12_18_port, A_neg_12_17_port, A_neg_12_16_port, A_neg_12_15_port, 
      A_neg_12_14_port, A_neg_12_13_port, A_neg_11_26_port, A_neg_11_25_port, 
      A_neg_11_24_port, A_neg_11_23_port, A_neg_11_22_port, A_neg_11_21_port, 
      A_neg_11_20_port, A_neg_11_19_port, A_neg_11_18_port, A_neg_11_17_port, 
      A_neg_11_16_port, A_neg_11_15_port, A_neg_11_14_port, A_neg_11_13_port, 
      A_neg_11_12_port, A_neg_10_25_port, A_neg_10_24_port, A_neg_10_23_port, 
      A_neg_10_22_port, A_neg_10_21_port, A_neg_10_20_port, A_neg_10_19_port, 
      A_neg_10_18_port, A_neg_10_17_port, A_neg_10_16_port, A_neg_10_15_port, 
      A_neg_10_14_port, A_neg_10_13_port, A_neg_10_12_port, A_neg_10_11_port, 
      A_neg_9_24_port, A_neg_9_23_port, A_neg_9_22_port, A_neg_9_21_port, 
      A_neg_9_20_port, A_neg_9_19_port, A_neg_9_18_port, A_neg_9_17_port, 
      A_neg_9_16_port, A_neg_9_15_port, A_neg_9_14_port, A_neg_9_13_port, 
      A_neg_9_12_port, A_neg_9_11_port, A_neg_9_10_port, A_neg_8_23_port, 
      A_neg_8_22_port, A_neg_8_21_port, A_neg_8_20_port, A_neg_8_19_port, 
      A_neg_8_18_port, A_neg_8_17_port, A_neg_8_16_port, A_neg_8_15_port, 
      A_neg_8_14_port, A_neg_8_13_port, A_neg_8_12_port, A_neg_8_11_port, 
      A_neg_8_10_port, A_neg_8_9_port, A_neg_7_22_port, A_neg_7_21_port, 
      A_neg_7_20_port, A_neg_7_19_port, A_neg_7_18_port, A_neg_7_17_port, 
      A_neg_7_16_port, A_neg_7_15_port, A_neg_7_14_port, A_neg_7_13_port, 
      A_neg_7_12_port, A_neg_7_11_port, A_neg_7_10_port, A_neg_7_9_port, 
      A_neg_7_8_port, A_neg_6_21_port, A_neg_6_20_port, A_neg_6_19_port, 
      A_neg_6_18_port, A_neg_6_17_port, A_neg_6_16_port, A_neg_6_15_port, 
      A_neg_6_14_port, A_neg_6_13_port, A_neg_6_12_port, A_neg_6_11_port, 
      A_neg_6_10_port, A_neg_6_9_port, A_neg_6_8_port, A_neg_6_7_port, 
      A_neg_5_20_port, A_neg_5_19_port, A_neg_5_18_port, A_neg_5_17_port, 
      A_neg_5_16_port, A_neg_5_15_port, A_neg_5_14_port, A_neg_5_13_port, 
      A_neg_5_12_port, A_neg_5_11_port, A_neg_5_10_port, A_neg_5_9_port, 
      A_neg_5_8_port, A_neg_5_7_port, A_neg_5_6_port, A_neg_4_19_port, 
      A_neg_4_18_port, A_neg_4_17_port, A_neg_4_16_port, A_neg_4_15_port, 
      A_neg_4_14_port, A_neg_4_13_port, A_neg_4_12_port, A_neg_4_11_port, 
      A_neg_4_10_port, A_neg_4_9_port, A_neg_4_8_port, A_neg_4_7_port, 
      A_neg_4_6_port, A_neg_4_5_port, A_neg_3_18_port, A_neg_3_17_port, 
      A_neg_3_16_port, A_neg_3_15_port, A_neg_3_14_port, A_neg_3_13_port, 
      A_neg_3_12_port, A_neg_3_11_port, A_neg_3_10_port, A_neg_3_9_port, 
      A_neg_3_8_port, A_neg_3_7_port, A_neg_3_6_port, A_neg_3_5_port, 
      A_neg_3_4_port, A_neg_2_17_port, A_neg_2_16_port, A_neg_2_15_port, 
      A_neg_2_14_port, A_neg_2_13_port, A_neg_2_12_port, A_neg_2_11_port, 
      A_neg_2_10_port, A_neg_2_9_port, A_neg_2_8_port, A_neg_2_7_port, 
      A_neg_2_6_port, A_neg_2_5_port, A_neg_2_4_port, A_neg_2_3_port, 
      A_neg_1_16_port, A_neg_1_15_port, A_neg_1_14_port, A_neg_1_13_port, 
      A_neg_1_12_port, A_neg_1_11_port, A_neg_1_10_port, A_neg_1_9_port, 
      A_neg_1_8_port, A_neg_1_7_port, A_neg_1_6_port, A_neg_1_5_port, 
      A_neg_1_4_port, A_neg_1_3_port, A_neg_1_2_port, A_neg_0_15_port, 
      A_neg_0_14_port, A_neg_0_13_port, A_neg_0_12_port, A_neg_0_11_port, 
      A_neg_0_10_port, A_neg_0_9_port, A_neg_0_8_port, A_neg_0_7_port, 
      A_neg_0_6_port, A_neg_0_5_port, A_neg_0_4_port, A_neg_0_3_port, 
      A_neg_0_2_port, A_neg_0_1_port, mux_out_7_31_port, mux_out_7_30_port, 
      mux_out_7_29_port, mux_out_7_28_port, mux_out_7_27_port, 
      mux_out_7_26_port, mux_out_7_25_port, mux_out_7_24_port, 
      mux_out_7_23_port, mux_out_7_22_port, mux_out_7_21_port, 
      mux_out_7_20_port, mux_out_7_19_port, mux_out_7_18_port, 
      mux_out_7_17_port, mux_out_7_16_port, mux_out_7_15_port, 
      mux_out_7_14_port, mux_out_7_13_port, mux_out_7_12_port, 
      mux_out_7_11_port, mux_out_7_10_port, mux_out_7_9_port, mux_out_7_8_port,
      mux_out_7_7_port, mux_out_7_6_port, mux_out_7_5_port, mux_out_7_4_port, 
      mux_out_7_3_port, mux_out_7_2_port, mux_out_7_1_port, mux_out_7_0_port, 
      mux_out_6_31_port, mux_out_6_30_port, mux_out_6_29_port, 
      mux_out_6_28_port, mux_out_6_27_port, mux_out_6_26_port, 
      mux_out_6_25_port, mux_out_6_24_port, mux_out_6_23_port, 
      mux_out_6_22_port, mux_out_6_21_port, mux_out_6_20_port, 
      mux_out_6_19_port, mux_out_6_18_port, mux_out_6_17_port, 
      mux_out_6_16_port, mux_out_6_15_port, mux_out_6_14_port, 
      mux_out_6_13_port, mux_out_6_12_port, mux_out_6_11_port, 
      mux_out_6_10_port, mux_out_6_9_port, mux_out_6_8_port, mux_out_6_7_port, 
      mux_out_6_6_port, mux_out_6_5_port, mux_out_6_4_port, mux_out_6_3_port, 
      mux_out_6_2_port, mux_out_6_1_port, mux_out_6_0_port, mux_out_5_31_port, 
      mux_out_5_30_port, mux_out_5_29_port, mux_out_5_28_port, 
      mux_out_5_27_port, mux_out_5_26_port, mux_out_5_25_port, 
      mux_out_5_24_port, mux_out_5_23_port, mux_out_5_22_port, 
      mux_out_5_21_port, mux_out_5_20_port, mux_out_5_19_port, 
      mux_out_5_18_port, mux_out_5_17_port, mux_out_5_16_port, 
      mux_out_5_15_port, mux_out_5_14_port, mux_out_5_13_port, 
      mux_out_5_12_port, mux_out_5_11_port, mux_out_5_10_port, mux_out_5_9_port
      , mux_out_5_8_port, mux_out_5_7_port, mux_out_5_6_port, mux_out_5_5_port,
      mux_out_5_4_port, mux_out_5_3_port, mux_out_5_2_port, mux_out_5_1_port, 
      mux_out_5_0_port, mux_out_4_31_port, mux_out_4_30_port, mux_out_4_29_port
      , mux_out_4_28_port, mux_out_4_27_port, mux_out_4_26_port, 
      mux_out_4_25_port, mux_out_4_24_port, mux_out_4_23_port, 
      mux_out_4_22_port, mux_out_4_21_port, mux_out_4_20_port, 
      mux_out_4_19_port, mux_out_4_18_port, mux_out_4_17_port, 
      mux_out_4_16_port, mux_out_4_15_port, mux_out_4_14_port, 
      mux_out_4_13_port, mux_out_4_12_port, mux_out_4_11_port, 
      mux_out_4_10_port, mux_out_4_9_port, mux_out_4_8_port, mux_out_4_7_port, 
      mux_out_4_6_port, mux_out_4_5_port, mux_out_4_4_port, mux_out_4_3_port, 
      mux_out_4_2_port, mux_out_4_1_port, mux_out_4_0_port, mux_out_3_31_port, 
      mux_out_3_30_port, mux_out_3_29_port, mux_out_3_28_port, 
      mux_out_3_27_port, mux_out_3_26_port, mux_out_3_25_port, 
      mux_out_3_24_port, mux_out_3_23_port, mux_out_3_22_port, 
      mux_out_3_21_port, mux_out_3_20_port, mux_out_3_19_port, 
      mux_out_3_18_port, mux_out_3_17_port, mux_out_3_16_port, 
      mux_out_3_15_port, mux_out_3_14_port, mux_out_3_13_port, 
      mux_out_3_12_port, mux_out_3_11_port, mux_out_3_10_port, mux_out_3_9_port
      , mux_out_3_8_port, mux_out_3_7_port, mux_out_3_6_port, mux_out_3_5_port,
      mux_out_3_4_port, mux_out_3_3_port, mux_out_3_2_port, mux_out_3_1_port, 
      mux_out_3_0_port, mux_out_2_31_port, mux_out_2_30_port, mux_out_2_29_port
      , mux_out_2_28_port, mux_out_2_27_port, mux_out_2_26_port, 
      mux_out_2_25_port, mux_out_2_24_port, mux_out_2_23_port, 
      mux_out_2_22_port, mux_out_2_21_port, mux_out_2_20_port, 
      mux_out_2_19_port, mux_out_2_18_port, mux_out_2_17_port, 
      mux_out_2_16_port, mux_out_2_15_port, mux_out_2_14_port, 
      mux_out_2_13_port, mux_out_2_12_port, mux_out_2_11_port, 
      mux_out_2_10_port, mux_out_2_9_port, mux_out_2_8_port, mux_out_2_7_port, 
      mux_out_2_6_port, mux_out_2_5_port, mux_out_2_4_port, mux_out_2_3_port, 
      mux_out_2_2_port, mux_out_2_1_port, mux_out_2_0_port, addends_7_31_port, 
      addends_7_30_port, addends_7_29_port, addends_7_28_port, 
      addends_7_27_port, addends_7_26_port, addends_7_25_port, 
      addends_7_24_port, addends_7_23_port, addends_7_22_port, 
      addends_7_21_port, addends_7_20_port, addends_7_19_port, 
      addends_7_18_port, addends_7_17_port, addends_7_16_port, 
      addends_7_15_port, addends_7_14_port, addends_7_13_port, 
      addends_7_12_port, addends_7_11_port, addends_7_10_port, addends_7_9_port
      , addends_7_8_port, addends_7_7_port, addends_7_6_port, addends_7_5_port,
      addends_7_4_port, addends_7_3_port, addends_7_2_port, addends_7_1_port, 
      addends_7_0_port, addends_6_31_port, addends_6_30_port, addends_6_29_port
      , addends_6_28_port, addends_6_27_port, addends_6_26_port, 
      addends_6_25_port, addends_6_24_port, addends_6_23_port, 
      addends_6_22_port, addends_6_21_port, addends_6_20_port, 
      addends_6_19_port, addends_6_18_port, addends_6_17_port, 
      addends_6_16_port, addends_6_15_port, addends_6_14_port, 
      addends_6_13_port, addends_6_12_port, addends_6_11_port, 
      addends_6_10_port, addends_6_9_port, addends_6_8_port, addends_6_7_port, 
      addends_6_6_port, addends_6_5_port, addends_6_4_port, addends_6_3_port, 
      addends_6_2_port, addends_6_1_port, addends_6_0_port, addends_5_31_port, 
      addends_5_30_port, addends_5_29_port, addends_5_28_port, 
      addends_5_27_port, addends_5_26_port, addends_5_25_port, 
      addends_5_24_port, addends_5_23_port, addends_5_22_port, 
      addends_5_21_port, addends_5_20_port, addends_5_19_port, 
      addends_5_18_port, addends_5_17_port, addends_5_16_port, 
      addends_5_15_port, addends_5_14_port, addends_5_13_port, 
      addends_5_12_port, addends_5_11_port, addends_5_10_port, addends_5_9_port
      , addends_5_8_port, addends_5_7_port, addends_5_6_port, addends_5_5_port,
      addends_5_4_port, addends_5_3_port, addends_5_2_port, addends_5_1_port, 
      addends_5_0_port, addends_4_31_port, addends_4_30_port, addends_4_29_port
      , addends_4_28_port, addends_4_27_port, addends_4_26_port, 
      addends_4_25_port, addends_4_24_port, addends_4_23_port, 
      addends_4_22_port, addends_4_21_port, addends_4_20_port, 
      addends_4_19_port, addends_4_18_port, addends_4_17_port, 
      addends_4_16_port, addends_4_15_port, addends_4_14_port, 
      addends_4_13_port, addends_4_12_port, addends_4_11_port, 
      addends_4_10_port, addends_4_9_port, addends_4_8_port, addends_4_7_port, 
      addends_4_6_port, addends_4_5_port, addends_4_4_port, addends_4_3_port, 
      addends_4_2_port, addends_4_1_port, addends_4_0_port, addends_3_31_port, 
      addends_3_30_port, addends_3_29_port, addends_3_28_port, 
      addends_3_27_port, addends_3_26_port, addends_3_25_port, 
      addends_3_24_port, addends_3_23_port, addends_3_22_port, 
      addends_3_21_port, addends_3_20_port, addends_3_19_port, 
      addends_3_18_port, addends_3_17_port, addends_3_16_port, 
      addends_3_15_port, addends_3_14_port, addends_3_13_port, 
      addends_3_12_port, addends_3_11_port, addends_3_10_port, addends_3_9_port
      , addends_3_8_port, addends_3_7_port, addends_3_6_port, addends_3_5_port,
      addends_3_4_port, addends_3_3_port, addends_3_2_port, addends_3_1_port, 
      addends_3_0_port, addends_2_31_port, addends_2_30_port, addends_2_29_port
      , addends_2_28_port, addends_2_27_port, addends_2_26_port, 
      addends_2_25_port, addends_2_24_port, addends_2_23_port, 
      addends_2_22_port, addends_2_21_port, addends_2_20_port, 
      addends_2_19_port, addends_2_18_port, addends_2_17_port, 
      addends_2_16_port, addends_2_15_port, addends_2_14_port, 
      addends_2_13_port, addends_2_12_port, addends_2_11_port, 
      addends_2_10_port, addends_2_9_port, addends_2_8_port, addends_2_7_port, 
      addends_2_6_port, addends_2_5_port, addends_2_4_port, addends_2_3_port, 
      addends_2_2_port, addends_2_1_port, addends_2_0_port, addends_1_31_port, 
      addends_1_30_port, addends_1_29_port, addends_1_28_port, 
      addends_1_27_port, addends_1_26_port, addends_1_25_port, 
      addends_1_24_port, addends_1_23_port, addends_1_22_port, 
      addends_1_21_port, addends_1_20_port, addends_1_19_port, 
      addends_1_18_port, addends_1_17_port, addends_1_16_port, 
      addends_1_15_port, addends_1_14_port, addends_1_13_port, 
      addends_1_12_port, addends_1_11_port, addends_1_10_port, addends_1_9_port
      , addends_1_8_port, addends_1_7_port, addends_1_6_port, addends_1_5_port,
      addends_1_4_port, addends_1_3_port, addends_1_2_port, addends_1_1_port, 
      addends_1_0_port, addends_0_31_port, addends_0_30_port, addends_0_29_port
      , addends_0_28_port, addends_0_27_port, addends_0_26_port, 
      addends_0_25_port, addends_0_24_port, addends_0_23_port, 
      addends_0_22_port, addends_0_21_port, addends_0_20_port, 
      addends_0_19_port, addends_0_18_port, addends_0_17_port, 
      addends_0_16_port, addends_0_15_port, addends_0_14_port, 
      addends_0_13_port, addends_0_12_port, addends_0_11_port, 
      addends_0_10_port, addends_0_9_port, addends_0_8_port, addends_0_7_port, 
      addends_0_6_port, addends_0_5_port, addends_0_4_port, addends_0_3_port, 
      addends_0_2_port, addends_0_1_port, addends_0_0_port, pipe1_3_31_port, 
      pipe1_3_30_port, pipe1_3_29_port, pipe1_3_28_port, pipe1_3_27_port, 
      pipe1_3_26_port, pipe1_3_25_port, pipe1_3_24_port, pipe1_3_23_port, 
      pipe1_3_22_port, pipe1_3_21_port, pipe1_3_20_port, pipe1_3_19_port, 
      pipe1_3_18_port, pipe1_3_17_port, pipe1_3_16_port, pipe1_3_15_port, 
      pipe1_3_14_port, pipe1_3_13_port, pipe1_3_12_port, pipe1_3_11_port, 
      pipe1_3_10_port, pipe1_3_9_port, pipe1_3_8_port, pipe1_3_7_port, 
      pipe1_3_6_port, pipe1_3_5_port, pipe1_3_4_port, pipe1_3_3_port, 
      pipe1_3_2_port, pipe1_3_1_port, pipe1_3_0_port, pipe1_2_31_port, 
      pipe1_2_30_port, pipe1_2_29_port, pipe1_2_28_port, pipe1_2_27_port, 
      pipe1_2_26_port, pipe1_2_25_port, pipe1_2_24_port, pipe1_2_23_port, 
      pipe1_2_22_port, pipe1_2_21_port, pipe1_2_20_port, pipe1_2_19_port, 
      pipe1_2_18_port, pipe1_2_17_port, pipe1_2_16_port, pipe1_2_15_port, 
      pipe1_2_14_port, pipe1_2_13_port, pipe1_2_12_port, pipe1_2_11_port, 
      pipe1_2_10_port, pipe1_2_9_port, pipe1_2_8_port, pipe1_2_7_port, 
      pipe1_2_6_port, pipe1_2_5_port, pipe1_2_4_port, pipe1_2_3_port, 
      pipe1_2_2_port, pipe1_2_1_port, pipe1_2_0_port, pipe1_1_31_port, 
      pipe1_1_30_port, pipe1_1_29_port, pipe1_1_28_port, pipe1_1_27_port, 
      pipe1_1_26_port, pipe1_1_25_port, pipe1_1_24_port, pipe1_1_23_port, 
      pipe1_1_22_port, pipe1_1_21_port, pipe1_1_20_port, pipe1_1_19_port, 
      pipe1_1_18_port, pipe1_1_17_port, pipe1_1_16_port, pipe1_1_15_port, 
      pipe1_1_14_port, pipe1_1_13_port, pipe1_1_12_port, pipe1_1_11_port, 
      pipe1_1_10_port, pipe1_1_9_port, pipe1_1_8_port, pipe1_1_7_port, 
      pipe1_1_6_port, pipe1_1_5_port, pipe1_1_4_port, pipe1_1_3_port, 
      pipe1_1_2_port, pipe1_1_1_port, pipe1_1_0_port, pipe1_0_31_port, 
      pipe1_0_30_port, pipe1_0_29_port, pipe1_0_28_port, pipe1_0_27_port, 
      pipe1_0_26_port, pipe1_0_25_port, pipe1_0_24_port, pipe1_0_23_port, 
      pipe1_0_22_port, pipe1_0_21_port, pipe1_0_20_port, pipe1_0_19_port, 
      pipe1_0_18_port, pipe1_0_17_port, pipe1_0_16_port, pipe1_0_15_port, 
      pipe1_0_14_port, pipe1_0_13_port, pipe1_0_12_port, pipe1_0_11_port, 
      pipe1_0_10_port, pipe1_0_9_port, pipe1_0_8_port, pipe1_0_7_port, 
      pipe1_0_6_port, pipe1_0_5_port, pipe1_0_4_port, pipe1_0_3_port, 
      pipe1_0_2_port, pipe1_0_1_port, pipe1_0_0_port, pipe2_1_31_port, 
      pipe2_1_30_port, pipe2_1_29_port, pipe2_1_28_port, pipe2_1_27_port, 
      pipe2_1_26_port, pipe2_1_25_port, pipe2_1_24_port, pipe2_1_23_port, 
      pipe2_1_22_port, pipe2_1_21_port, pipe2_1_20_port, pipe2_1_19_port, 
      pipe2_1_18_port, pipe2_1_17_port, pipe2_1_16_port, pipe2_1_15_port, 
      pipe2_1_14_port, pipe2_1_13_port, pipe2_1_12_port, pipe2_1_11_port, 
      pipe2_1_10_port, pipe2_1_9_port, pipe2_1_8_port, pipe2_1_7_port, 
      pipe2_1_6_port, pipe2_1_5_port, pipe2_1_4_port, pipe2_1_3_port, 
      pipe2_1_2_port, pipe2_1_1_port, pipe2_1_0_port, pipe2_0_31_port, 
      pipe2_0_30_port, pipe2_0_29_port, pipe2_0_28_port, pipe2_0_27_port, 
      pipe2_0_26_port, pipe2_0_25_port, pipe2_0_24_port, pipe2_0_23_port, 
      pipe2_0_22_port, pipe2_0_21_port, pipe2_0_20_port, pipe2_0_19_port, 
      pipe2_0_18_port, pipe2_0_17_port, pipe2_0_16_port, pipe2_0_15_port, 
      pipe2_0_14_port, pipe2_0_13_port, pipe2_0_12_port, pipe2_0_11_port, 
      pipe2_0_10_port, pipe2_0_9_port, pipe2_0_8_port, pipe2_0_7_port, 
      pipe2_0_6_port, pipe2_0_5_port, pipe2_0_4_port, pipe2_0_3_port, 
      pipe2_0_2_port, pipe2_0_1_port, pipe2_0_0_port, selector_23_port, 
      selector_22_port, selector_21_port, selector_20_port, selector_19_port, 
      selector_18_port, selector_17_port, selector_16_port, selector_15_port, 
      selector_14_port, selector_13_port, selector_12_port, selector_11_port, 
      selector_10_port, selector_9_port, selector_8_port, selector_7_port, 
      selector_6_port, selector_5_port, selector_4_port, selector_3_port, 
      selector_2_port, selector_1_port, selector_0_port, reg_in_2_31_port, 
      reg_in_2_30_port, reg_in_2_29_port, reg_in_2_28_port, reg_in_2_27_port, 
      reg_in_2_26_port, reg_in_2_25_port, reg_in_2_24_port, reg_in_2_23_port, 
      reg_in_2_22_port, reg_in_2_21_port, reg_in_2_20_port, reg_in_2_19_port, 
      reg_in_2_18_port, reg_in_2_17_port, reg_in_2_16_port, reg_in_2_15_port, 
      reg_in_2_14_port, reg_in_2_13_port, reg_in_2_12_port, reg_in_2_11_port, 
      reg_in_2_10_port, reg_in_2_9_port, reg_in_2_8_port, reg_in_2_7_port, 
      reg_in_2_6_port, reg_in_2_5_port, reg_in_2_4_port, reg_in_2_3_port, 
      reg_in_2_2_port, reg_in_2_1_port, reg_in_2_0_port, reg_in_1_31_port, 
      reg_in_1_30_port, reg_in_1_29_port, reg_in_1_28_port, reg_in_1_27_port, 
      reg_in_1_26_port, reg_in_1_25_port, reg_in_1_24_port, reg_in_1_23_port, 
      reg_in_1_22_port, reg_in_1_21_port, reg_in_1_20_port, reg_in_1_19_port, 
      reg_in_1_18_port, reg_in_1_17_port, reg_in_1_16_port, reg_in_1_15_port, 
      reg_in_1_14_port, reg_in_1_13_port, reg_in_1_12_port, reg_in_1_11_port, 
      reg_in_1_10_port, reg_in_1_9_port, reg_in_1_8_port, reg_in_1_7_port, 
      reg_in_1_6_port, reg_in_1_5_port, reg_in_1_4_port, reg_in_1_3_port, 
      reg_in_1_2_port, reg_in_1_1_port, reg_in_1_0_port, reg_in_0_31_port, 
      reg_in_0_30_port, reg_in_0_29_port, reg_in_0_28_port, reg_in_0_27_port, 
      reg_in_0_26_port, reg_in_0_25_port, reg_in_0_24_port, reg_in_0_23_port, 
      reg_in_0_22_port, reg_in_0_21_port, reg_in_0_20_port, reg_in_0_19_port, 
      reg_in_0_18_port, reg_in_0_17_port, reg_in_0_16_port, reg_in_0_15_port, 
      reg_in_0_14_port, reg_in_0_13_port, reg_in_0_12_port, reg_in_0_11_port, 
      reg_in_0_10_port, reg_in_0_9_port, reg_in_0_8_port, reg_in_0_7_port, 
      reg_in_0_6_port, reg_in_0_5_port, reg_in_0_4_port, reg_in_0_3_port, 
      reg_in_0_2_port, reg_in_0_1_port, reg_in_0_0_port, reg_out_2_31_port, 
      reg_out_2_30_port, reg_out_2_29_port, reg_out_2_28_port, 
      reg_out_2_27_port, reg_out_2_26_port, reg_out_2_25_port, 
      reg_out_2_24_port, reg_out_2_23_port, reg_out_2_22_port, 
      reg_out_2_21_port, reg_out_2_20_port, reg_out_2_19_port, 
      reg_out_2_18_port, reg_out_2_17_port, reg_out_2_16_port, 
      reg_out_2_15_port, reg_out_2_14_port, reg_out_2_13_port, 
      reg_out_2_12_port, reg_out_2_11_port, reg_out_2_10_port, reg_out_2_9_port
      , reg_out_2_8_port, reg_out_2_7_port, reg_out_2_6_port, reg_out_2_5_port,
      reg_out_2_4_port, reg_out_2_3_port, reg_out_2_2_port, reg_out_2_1_port, 
      reg_out_2_0_port, reg_out_1_31_port, reg_out_1_30_port, reg_out_1_29_port
      , reg_out_1_28_port, reg_out_1_27_port, reg_out_1_26_port, 
      reg_out_1_25_port, reg_out_1_24_port, reg_out_1_23_port, 
      reg_out_1_22_port, reg_out_1_21_port, reg_out_1_20_port, 
      reg_out_1_19_port, reg_out_1_18_port, reg_out_1_17_port, 
      reg_out_1_16_port, reg_out_1_15_port, reg_out_1_14_port, 
      reg_out_1_13_port, reg_out_1_12_port, reg_out_1_11_port, 
      reg_out_1_10_port, reg_out_1_9_port, reg_out_1_8_port, reg_out_1_7_port, 
      reg_out_1_6_port, reg_out_1_5_port, reg_out_1_4_port, reg_out_1_3_port, 
      reg_out_1_2_port, reg_out_1_1_port, reg_out_1_0_port, reg_out_0_31_port, 
      reg_out_0_30_port, reg_out_0_29_port, reg_out_0_28_port, 
      reg_out_0_27_port, reg_out_0_26_port, reg_out_0_25_port, 
      reg_out_0_24_port, reg_out_0_23_port, reg_out_0_22_port, 
      reg_out_0_21_port, reg_out_0_20_port, reg_out_0_19_port, 
      reg_out_0_18_port, reg_out_0_17_port, reg_out_0_16_port, 
      reg_out_0_15_port, reg_out_0_14_port, reg_out_0_13_port, 
      reg_out_0_12_port, reg_out_0_11_port, reg_out_0_10_port, reg_out_0_9_port
      , reg_out_0_8_port, reg_out_0_7_port, reg_out_0_6_port, reg_out_0_5_port,
      reg_out_0_4_port, reg_out_0_3_port, reg_out_0_2_port, reg_out_0_1_port, 
      reg_out_0_0_port, add_out_2_31_port, add_out_2_30_port, add_out_2_29_port
      , add_out_2_28_port, add_out_2_27_port, add_out_2_26_port, 
      add_out_2_25_port, add_out_2_24_port, add_out_2_23_port, 
      add_out_2_22_port, add_out_2_21_port, add_out_2_20_port, 
      add_out_2_19_port, add_out_2_18_port, add_out_2_17_port, 
      add_out_2_16_port, add_out_2_15_port, add_out_2_14_port, 
      add_out_2_13_port, add_out_2_12_port, add_out_2_11_port, 
      add_out_2_10_port, add_out_2_9_port, add_out_2_8_port, add_out_2_7_port, 
      add_out_2_6_port, add_out_2_5_port, add_out_2_4_port, add_out_2_3_port, 
      add_out_2_2_port, add_out_2_1_port, add_out_2_0_port, add_out_1_31_port, 
      add_out_1_30_port, add_out_1_29_port, add_out_1_28_port, 
      add_out_1_27_port, add_out_1_26_port, add_out_1_25_port, 
      add_out_1_24_port, add_out_1_23_port, add_out_1_22_port, 
      add_out_1_21_port, add_out_1_20_port, add_out_1_19_port, 
      add_out_1_18_port, add_out_1_17_port, add_out_1_16_port, 
      add_out_1_15_port, add_out_1_14_port, add_out_1_13_port, 
      add_out_1_12_port, add_out_1_11_port, add_out_1_10_port, add_out_1_9_port
      , add_out_1_8_port, add_out_1_7_port, add_out_1_6_port, add_out_1_5_port,
      add_out_1_4_port, add_out_1_3_port, add_out_1_2_port, add_out_1_1_port, 
      add_out_1_0_port, add_out_0_31_port, add_out_0_30_port, add_out_0_29_port
      , add_out_0_28_port, add_out_0_27_port, add_out_0_26_port, 
      add_out_0_25_port, add_out_0_24_port, add_out_0_23_port, 
      add_out_0_22_port, add_out_0_21_port, add_out_0_20_port, 
      add_out_0_19_port, add_out_0_18_port, add_out_0_17_port, 
      add_out_0_16_port, add_out_0_15_port, add_out_0_14_port, 
      add_out_0_13_port, add_out_0_12_port, add_out_0_11_port, 
      add_out_0_10_port, add_out_0_9_port, add_out_0_8_port, add_out_0_7_port, 
      add_out_0_6_port, add_out_0_5_port, add_out_0_4_port, add_out_0_3_port, 
      add_out_0_2_port, add_out_0_1_port, add_out_0_0_port, 
      sub_126_G16_carry_17_port, sub_126_G16_carry_18_port, 
      sub_126_G16_carry_19_port, sub_126_G16_carry_20_port, 
      sub_126_G16_carry_21_port, sub_126_G16_carry_22_port, 
      sub_126_G16_carry_23_port, sub_126_G16_carry_24_port, 
      sub_126_G16_carry_25_port, sub_126_G16_carry_26_port, 
      sub_126_G16_carry_27_port, sub_126_G16_carry_28_port, 
      sub_126_G16_carry_29_port, sub_126_G16_carry_30_port, 
      sub_126_G15_carry_16_port, sub_126_G15_carry_17_port, 
      sub_126_G15_carry_18_port, sub_126_G15_carry_19_port, 
      sub_126_G15_carry_20_port, sub_126_G15_carry_21_port, 
      sub_126_G15_carry_22_port, sub_126_G15_carry_23_port, 
      sub_126_G15_carry_24_port, sub_126_G15_carry_25_port, 
      sub_126_G15_carry_26_port, sub_126_G15_carry_27_port, 
      sub_126_G15_carry_28_port, sub_126_G15_carry_29_port, 
      sub_126_G14_carry_15_port, sub_126_G14_carry_16_port, 
      sub_126_G14_carry_17_port, sub_126_G14_carry_18_port, 
      sub_126_G14_carry_19_port, sub_126_G14_carry_20_port, 
      sub_126_G14_carry_21_port, sub_126_G14_carry_22_port, 
      sub_126_G14_carry_23_port, sub_126_G14_carry_24_port, 
      sub_126_G14_carry_25_port, sub_126_G14_carry_26_port, 
      sub_126_G14_carry_27_port, sub_126_G14_carry_28_port, 
      sub_126_G13_carry_14_port, sub_126_G13_carry_15_port, 
      sub_126_G13_carry_16_port, sub_126_G13_carry_17_port, 
      sub_126_G13_carry_18_port, sub_126_G13_carry_19_port, 
      sub_126_G13_carry_20_port, sub_126_G13_carry_21_port, 
      sub_126_G13_carry_22_port, sub_126_G13_carry_23_port, 
      sub_126_G13_carry_24_port, sub_126_G13_carry_25_port, 
      sub_126_G13_carry_26_port, sub_126_G13_carry_27_port, 
      sub_126_G12_carry_13_port, sub_126_G12_carry_14_port, 
      sub_126_G12_carry_15_port, sub_126_G12_carry_16_port, 
      sub_126_G12_carry_17_port, sub_126_G12_carry_18_port, 
      sub_126_G12_carry_19_port, sub_126_G12_carry_20_port, 
      sub_126_G12_carry_21_port, sub_126_G12_carry_22_port, 
      sub_126_G12_carry_23_port, sub_126_G12_carry_24_port, 
      sub_126_G12_carry_25_port, sub_126_G12_carry_26_port, 
      sub_126_G11_carry_12_port, sub_126_G11_carry_13_port, 
      sub_126_G11_carry_14_port, sub_126_G11_carry_15_port, 
      sub_126_G11_carry_16_port, sub_126_G11_carry_17_port, 
      sub_126_G11_carry_18_port, sub_126_G11_carry_19_port, 
      sub_126_G11_carry_20_port, sub_126_G11_carry_21_port, 
      sub_126_G11_carry_22_port, sub_126_G11_carry_23_port, 
      sub_126_G11_carry_24_port, sub_126_G11_carry_25_port, 
      sub_126_G10_carry_11_port, sub_126_G10_carry_12_port, 
      sub_126_G10_carry_13_port, sub_126_G10_carry_14_port, 
      sub_126_G10_carry_15_port, sub_126_G10_carry_16_port, 
      sub_126_G10_carry_17_port, sub_126_G10_carry_18_port, 
      sub_126_G10_carry_19_port, sub_126_G10_carry_20_port, 
      sub_126_G10_carry_21_port, sub_126_G10_carry_22_port, 
      sub_126_G10_carry_23_port, sub_126_G10_carry_24_port, 
      sub_126_G9_carry_10_port, sub_126_G9_carry_11_port, 
      sub_126_G9_carry_12_port, sub_126_G9_carry_13_port, 
      sub_126_G9_carry_14_port, sub_126_G9_carry_15_port, 
      sub_126_G9_carry_16_port, sub_126_G9_carry_17_port, 
      sub_126_G9_carry_18_port, sub_126_G9_carry_19_port, 
      sub_126_G9_carry_20_port, sub_126_G9_carry_21_port, 
      sub_126_G9_carry_22_port, sub_126_G9_carry_23_port, 
      sub_126_G8_carry_9_port, sub_126_G8_carry_10_port, 
      sub_126_G8_carry_11_port, sub_126_G8_carry_12_port, 
      sub_126_G8_carry_13_port, sub_126_G8_carry_14_port, 
      sub_126_G8_carry_15_port, sub_126_G8_carry_16_port, 
      sub_126_G8_carry_17_port, sub_126_G8_carry_18_port, 
      sub_126_G8_carry_19_port, sub_126_G8_carry_20_port, 
      sub_126_G8_carry_21_port, sub_126_G8_carry_22_port, 
      sub_126_G7_carry_8_port, sub_126_G7_carry_9_port, 
      sub_126_G7_carry_10_port, sub_126_G7_carry_11_port, 
      sub_126_G7_carry_12_port, sub_126_G7_carry_13_port, 
      sub_126_G7_carry_14_port, sub_126_G7_carry_15_port, 
      sub_126_G7_carry_16_port, sub_126_G7_carry_17_port, 
      sub_126_G7_carry_18_port, sub_126_G7_carry_19_port, 
      sub_126_G7_carry_20_port, sub_126_G7_carry_21_port, 
      sub_126_G6_carry_7_port, sub_126_G6_carry_8_port, sub_126_G6_carry_9_port
      , sub_126_G6_carry_10_port, sub_126_G6_carry_11_port, 
      sub_126_G6_carry_12_port, sub_126_G6_carry_13_port, 
      sub_126_G6_carry_14_port, sub_126_G6_carry_15_port, 
      sub_126_G6_carry_16_port, sub_126_G6_carry_17_port, 
      sub_126_G6_carry_18_port, sub_126_G6_carry_19_port, 
      sub_126_G6_carry_20_port, sub_126_G5_carry_6_port, 
      sub_126_G5_carry_7_port, sub_126_G5_carry_8_port, sub_126_G5_carry_9_port
      , sub_126_G5_carry_10_port, sub_126_G5_carry_11_port, 
      sub_126_G5_carry_12_port, sub_126_G5_carry_13_port, 
      sub_126_G5_carry_14_port, sub_126_G5_carry_15_port, 
      sub_126_G5_carry_16_port, sub_126_G5_carry_17_port, 
      sub_126_G5_carry_18_port, sub_126_G5_carry_19_port, 
      sub_126_G4_carry_5_port, sub_126_G4_carry_6_port, sub_126_G4_carry_7_port
      , sub_126_G4_carry_8_port, sub_126_G4_carry_9_port, 
      sub_126_G4_carry_10_port, sub_126_G4_carry_11_port, 
      sub_126_G4_carry_12_port, sub_126_G4_carry_13_port, 
      sub_126_G4_carry_14_port, sub_126_G4_carry_15_port, 
      sub_126_G4_carry_16_port, sub_126_G4_carry_17_port, 
      sub_126_G4_carry_18_port, sub_126_G3_carry_4_port, 
      sub_126_G3_carry_5_port, sub_126_G3_carry_6_port, sub_126_G3_carry_7_port
      , sub_126_G3_carry_8_port, sub_126_G3_carry_9_port, 
      sub_126_G3_carry_10_port, sub_126_G3_carry_11_port, 
      sub_126_G3_carry_12_port, sub_126_G3_carry_13_port, 
      sub_126_G3_carry_14_port, sub_126_G3_carry_15_port, 
      sub_126_G3_carry_16_port, sub_126_G3_carry_17_port, 
      sub_126_G2_carry_3_port, sub_126_G2_carry_4_port, sub_126_G2_carry_5_port
      , sub_126_G2_carry_6_port, sub_126_G2_carry_7_port, 
      sub_126_G2_carry_8_port, sub_126_G2_carry_9_port, 
      sub_126_G2_carry_10_port, sub_126_G2_carry_11_port, 
      sub_126_G2_carry_12_port, sub_126_G2_carry_13_port, 
      sub_126_G2_carry_14_port, sub_126_G2_carry_15_port, 
      sub_126_G2_carry_16_port, sub_126_carry_2_port, sub_126_carry_3_port, 
      sub_126_carry_4_port, sub_126_carry_5_port, sub_126_carry_6_port, 
      sub_126_carry_7_port, sub_126_carry_8_port, sub_126_carry_9_port, 
      sub_126_carry_10_port, sub_126_carry_11_port, sub_126_carry_12_port, 
      sub_126_carry_13_port, sub_126_carry_14_port, sub_126_carry_15_port, n1, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n_1171, n_1172, n_1173, n_1174,
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   addends_reg_3_31_inst : DFF_X1 port map( D => mux_out_3_31_port, CK => CLOCK
                           , Q => addends_3_31_port, QN => n_1171);
   addends_reg_3_30_inst : DFF_X1 port map( D => mux_out_3_30_port, CK => CLOCK
                           , Q => addends_3_30_port, QN => n_1172);
   addends_reg_3_29_inst : DFF_X1 port map( D => mux_out_3_29_port, CK => CLOCK
                           , Q => addends_3_29_port, QN => n_1173);
   addends_reg_3_28_inst : DFF_X1 port map( D => mux_out_3_28_port, CK => CLOCK
                           , Q => addends_3_28_port, QN => n_1174);
   addends_reg_3_27_inst : DFF_X1 port map( D => mux_out_3_27_port, CK => CLOCK
                           , Q => addends_3_27_port, QN => n_1175);
   addends_reg_3_26_inst : DFF_X1 port map( D => mux_out_3_26_port, CK => CLOCK
                           , Q => addends_3_26_port, QN => n_1176);
   addends_reg_3_25_inst : DFF_X1 port map( D => mux_out_3_25_port, CK => CLOCK
                           , Q => addends_3_25_port, QN => n_1177);
   addends_reg_3_24_inst : DFF_X1 port map( D => mux_out_3_24_port, CK => CLOCK
                           , Q => addends_3_24_port, QN => n_1178);
   addends_reg_3_23_inst : DFF_X1 port map( D => mux_out_3_23_port, CK => CLOCK
                           , Q => addends_3_23_port, QN => n_1179);
   addends_reg_3_22_inst : DFF_X1 port map( D => mux_out_3_22_port, CK => CLOCK
                           , Q => addends_3_22_port, QN => n_1180);
   addends_reg_3_21_inst : DFF_X1 port map( D => mux_out_3_21_port, CK => CLOCK
                           , Q => addends_3_21_port, QN => n_1181);
   addends_reg_3_20_inst : DFF_X1 port map( D => mux_out_3_20_port, CK => CLOCK
                           , Q => addends_3_20_port, QN => n_1182);
   addends_reg_3_19_inst : DFF_X1 port map( D => mux_out_3_19_port, CK => CLOCK
                           , Q => addends_3_19_port, QN => n_1183);
   addends_reg_3_18_inst : DFF_X1 port map( D => mux_out_3_18_port, CK => CLOCK
                           , Q => addends_3_18_port, QN => n_1184);
   addends_reg_3_17_inst : DFF_X1 port map( D => mux_out_3_17_port, CK => CLOCK
                           , Q => addends_3_17_port, QN => n_1185);
   addends_reg_3_16_inst : DFF_X1 port map( D => mux_out_3_16_port, CK => CLOCK
                           , Q => addends_3_16_port, QN => n_1186);
   addends_reg_3_15_inst : DFF_X1 port map( D => mux_out_3_15_port, CK => CLOCK
                           , Q => addends_3_15_port, QN => n_1187);
   addends_reg_3_14_inst : DFF_X1 port map( D => mux_out_3_14_port, CK => CLOCK
                           , Q => addends_3_14_port, QN => n_1188);
   addends_reg_3_13_inst : DFF_X1 port map( D => mux_out_3_13_port, CK => CLOCK
                           , Q => addends_3_13_port, QN => n_1189);
   addends_reg_3_12_inst : DFF_X1 port map( D => mux_out_3_12_port, CK => CLOCK
                           , Q => addends_3_12_port, QN => n_1190);
   addends_reg_3_11_inst : DFF_X1 port map( D => mux_out_3_11_port, CK => CLOCK
                           , Q => addends_3_11_port, QN => n_1191);
   addends_reg_3_10_inst : DFF_X1 port map( D => mux_out_3_10_port, CK => CLOCK
                           , Q => addends_3_10_port, QN => n_1192);
   addends_reg_3_9_inst : DFF_X1 port map( D => mux_out_3_9_port, CK => CLOCK, 
                           Q => addends_3_9_port, QN => n_1193);
   addends_reg_3_8_inst : DFF_X1 port map( D => mux_out_3_8_port, CK => CLOCK, 
                           Q => addends_3_8_port, QN => n_1194);
   addends_reg_3_7_inst : DFF_X1 port map( D => mux_out_3_7_port, CK => CLOCK, 
                           Q => addends_3_7_port, QN => n_1195);
   addends_reg_3_6_inst : DFF_X1 port map( D => mux_out_3_6_port, CK => CLOCK, 
                           Q => addends_3_6_port, QN => n_1196);
   addends_reg_3_5_inst : DFF_X1 port map( D => mux_out_3_5_port, CK => CLOCK, 
                           Q => addends_3_5_port, QN => n_1197);
   addends_reg_3_4_inst : DFF_X1 port map( D => mux_out_3_4_port, CK => CLOCK, 
                           Q => addends_3_4_port, QN => n_1198);
   addends_reg_3_3_inst : DFF_X1 port map( D => mux_out_3_3_port, CK => CLOCK, 
                           Q => addends_3_3_port, QN => n_1199);
   addends_reg_3_2_inst : DFF_X1 port map( D => mux_out_3_2_port, CK => CLOCK, 
                           Q => addends_3_2_port, QN => n_1200);
   addends_reg_3_1_inst : DFF_X1 port map( D => mux_out_3_1_port, CK => CLOCK, 
                           Q => addends_3_1_port, QN => n_1201);
   addends_reg_3_0_inst : DFF_X1 port map( D => mux_out_3_0_port, CK => CLOCK, 
                           Q => addends_3_0_port, QN => n_1202);
   addends_reg_2_31_inst : DFF_X1 port map( D => mux_out_2_31_port, CK => CLOCK
                           , Q => addends_2_31_port, QN => n_1203);
   addends_reg_2_30_inst : DFF_X1 port map( D => mux_out_2_30_port, CK => CLOCK
                           , Q => addends_2_30_port, QN => n_1204);
   addends_reg_2_29_inst : DFF_X1 port map( D => mux_out_2_29_port, CK => CLOCK
                           , Q => addends_2_29_port, QN => n_1205);
   addends_reg_2_28_inst : DFF_X1 port map( D => mux_out_2_28_port, CK => CLOCK
                           , Q => addends_2_28_port, QN => n_1206);
   addends_reg_2_27_inst : DFF_X1 port map( D => mux_out_2_27_port, CK => CLOCK
                           , Q => addends_2_27_port, QN => n_1207);
   addends_reg_2_26_inst : DFF_X1 port map( D => mux_out_2_26_port, CK => CLOCK
                           , Q => addends_2_26_port, QN => n_1208);
   addends_reg_2_25_inst : DFF_X1 port map( D => mux_out_2_25_port, CK => CLOCK
                           , Q => addends_2_25_port, QN => n_1209);
   addends_reg_2_24_inst : DFF_X1 port map( D => mux_out_2_24_port, CK => CLOCK
                           , Q => addends_2_24_port, QN => n_1210);
   addends_reg_2_23_inst : DFF_X1 port map( D => mux_out_2_23_port, CK => CLOCK
                           , Q => addends_2_23_port, QN => n_1211);
   addends_reg_2_22_inst : DFF_X1 port map( D => mux_out_2_22_port, CK => CLOCK
                           , Q => addends_2_22_port, QN => n_1212);
   addends_reg_2_21_inst : DFF_X1 port map( D => mux_out_2_21_port, CK => CLOCK
                           , Q => addends_2_21_port, QN => n_1213);
   addends_reg_2_20_inst : DFF_X1 port map( D => mux_out_2_20_port, CK => CLOCK
                           , Q => addends_2_20_port, QN => n_1214);
   addends_reg_2_19_inst : DFF_X1 port map( D => mux_out_2_19_port, CK => CLOCK
                           , Q => addends_2_19_port, QN => n_1215);
   addends_reg_2_18_inst : DFF_X1 port map( D => mux_out_2_18_port, CK => CLOCK
                           , Q => addends_2_18_port, QN => n_1216);
   addends_reg_2_17_inst : DFF_X1 port map( D => mux_out_2_17_port, CK => CLOCK
                           , Q => addends_2_17_port, QN => n_1217);
   addends_reg_2_16_inst : DFF_X1 port map( D => mux_out_2_16_port, CK => CLOCK
                           , Q => addends_2_16_port, QN => n_1218);
   addends_reg_2_15_inst : DFF_X1 port map( D => mux_out_2_15_port, CK => CLOCK
                           , Q => addends_2_15_port, QN => n_1219);
   addends_reg_2_14_inst : DFF_X1 port map( D => mux_out_2_14_port, CK => CLOCK
                           , Q => addends_2_14_port, QN => n_1220);
   addends_reg_2_13_inst : DFF_X1 port map( D => mux_out_2_13_port, CK => CLOCK
                           , Q => addends_2_13_port, QN => n_1221);
   addends_reg_2_12_inst : DFF_X1 port map( D => mux_out_2_12_port, CK => CLOCK
                           , Q => addends_2_12_port, QN => n_1222);
   addends_reg_2_11_inst : DFF_X1 port map( D => mux_out_2_11_port, CK => CLOCK
                           , Q => addends_2_11_port, QN => n_1223);
   addends_reg_2_10_inst : DFF_X1 port map( D => mux_out_2_10_port, CK => CLOCK
                           , Q => addends_2_10_port, QN => n_1224);
   addends_reg_2_9_inst : DFF_X1 port map( D => mux_out_2_9_port, CK => CLOCK, 
                           Q => addends_2_9_port, QN => n_1225);
   addends_reg_2_8_inst : DFF_X1 port map( D => mux_out_2_8_port, CK => CLOCK, 
                           Q => addends_2_8_port, QN => n_1226);
   addends_reg_2_7_inst : DFF_X1 port map( D => mux_out_2_7_port, CK => CLOCK, 
                           Q => addends_2_7_port, QN => n_1227);
   addends_reg_2_6_inst : DFF_X1 port map( D => mux_out_2_6_port, CK => CLOCK, 
                           Q => addends_2_6_port, QN => n_1228);
   addends_reg_2_5_inst : DFF_X1 port map( D => mux_out_2_5_port, CK => CLOCK, 
                           Q => addends_2_5_port, QN => n_1229);
   addends_reg_2_4_inst : DFF_X1 port map( D => mux_out_2_4_port, CK => CLOCK, 
                           Q => addends_2_4_port, QN => n_1230);
   addends_reg_2_3_inst : DFF_X1 port map( D => mux_out_2_3_port, CK => CLOCK, 
                           Q => addends_2_3_port, QN => n_1231);
   addends_reg_2_2_inst : DFF_X1 port map( D => mux_out_2_2_port, CK => CLOCK, 
                           Q => addends_2_2_port, QN => n_1232);
   addends_reg_2_1_inst : DFF_X1 port map( D => mux_out_2_1_port, CK => CLOCK, 
                           Q => addends_2_1_port, QN => n_1233);
   addends_reg_2_0_inst : DFF_X1 port map( D => mux_out_2_0_port, CK => CLOCK, 
                           Q => addends_2_0_port, QN => n_1234);
   pipe1_reg_3_31_inst : DFF_X1 port map( D => mux_out_7_31_port, CK => CLOCK, 
                           Q => pipe1_3_31_port, QN => n_1235);
   pipe1_reg_3_30_inst : DFF_X1 port map( D => mux_out_7_30_port, CK => CLOCK, 
                           Q => pipe1_3_30_port, QN => n_1236);
   pipe1_reg_3_29_inst : DFF_X1 port map( D => mux_out_7_29_port, CK => CLOCK, 
                           Q => pipe1_3_29_port, QN => n_1237);
   pipe1_reg_3_28_inst : DFF_X1 port map( D => mux_out_7_28_port, CK => CLOCK, 
                           Q => pipe1_3_28_port, QN => n_1238);
   pipe1_reg_3_27_inst : DFF_X1 port map( D => mux_out_7_27_port, CK => CLOCK, 
                           Q => pipe1_3_27_port, QN => n_1239);
   pipe1_reg_3_26_inst : DFF_X1 port map( D => mux_out_7_26_port, CK => CLOCK, 
                           Q => pipe1_3_26_port, QN => n_1240);
   pipe1_reg_3_25_inst : DFF_X1 port map( D => mux_out_7_25_port, CK => CLOCK, 
                           Q => pipe1_3_25_port, QN => n_1241);
   pipe1_reg_3_24_inst : DFF_X1 port map( D => mux_out_7_24_port, CK => CLOCK, 
                           Q => pipe1_3_24_port, QN => n_1242);
   pipe1_reg_3_23_inst : DFF_X1 port map( D => mux_out_7_23_port, CK => CLOCK, 
                           Q => pipe1_3_23_port, QN => n_1243);
   pipe1_reg_3_22_inst : DFF_X1 port map( D => mux_out_7_22_port, CK => CLOCK, 
                           Q => pipe1_3_22_port, QN => n_1244);
   pipe1_reg_3_21_inst : DFF_X1 port map( D => mux_out_7_21_port, CK => CLOCK, 
                           Q => pipe1_3_21_port, QN => n_1245);
   pipe1_reg_3_20_inst : DFF_X1 port map( D => mux_out_7_20_port, CK => CLOCK, 
                           Q => pipe1_3_20_port, QN => n_1246);
   pipe1_reg_3_19_inst : DFF_X1 port map( D => mux_out_7_19_port, CK => CLOCK, 
                           Q => pipe1_3_19_port, QN => n_1247);
   pipe1_reg_3_18_inst : DFF_X1 port map( D => mux_out_7_18_port, CK => CLOCK, 
                           Q => pipe1_3_18_port, QN => n_1248);
   pipe1_reg_3_17_inst : DFF_X1 port map( D => mux_out_7_17_port, CK => CLOCK, 
                           Q => pipe1_3_17_port, QN => n_1249);
   pipe1_reg_3_16_inst : DFF_X1 port map( D => mux_out_7_16_port, CK => CLOCK, 
                           Q => pipe1_3_16_port, QN => n_1250);
   pipe1_reg_3_15_inst : DFF_X1 port map( D => mux_out_7_15_port, CK => CLOCK, 
                           Q => pipe1_3_15_port, QN => n_1251);
   pipe1_reg_3_14_inst : DFF_X1 port map( D => mux_out_7_14_port, CK => CLOCK, 
                           Q => pipe1_3_14_port, QN => n_1252);
   pipe1_reg_3_13_inst : DFF_X1 port map( D => mux_out_7_13_port, CK => CLOCK, 
                           Q => pipe1_3_13_port, QN => n_1253);
   pipe1_reg_3_12_inst : DFF_X1 port map( D => mux_out_7_12_port, CK => CLOCK, 
                           Q => pipe1_3_12_port, QN => n_1254);
   pipe1_reg_3_11_inst : DFF_X1 port map( D => mux_out_7_11_port, CK => CLOCK, 
                           Q => pipe1_3_11_port, QN => n_1255);
   pipe1_reg_3_10_inst : DFF_X1 port map( D => mux_out_7_10_port, CK => CLOCK, 
                           Q => pipe1_3_10_port, QN => n_1256);
   pipe1_reg_3_9_inst : DFF_X1 port map( D => mux_out_7_9_port, CK => CLOCK, Q 
                           => pipe1_3_9_port, QN => n_1257);
   pipe1_reg_3_8_inst : DFF_X1 port map( D => mux_out_7_8_port, CK => CLOCK, Q 
                           => pipe1_3_8_port, QN => n_1258);
   pipe1_reg_3_7_inst : DFF_X1 port map( D => mux_out_7_7_port, CK => CLOCK, Q 
                           => pipe1_3_7_port, QN => n_1259);
   pipe1_reg_3_6_inst : DFF_X1 port map( D => mux_out_7_6_port, CK => CLOCK, Q 
                           => pipe1_3_6_port, QN => n_1260);
   pipe1_reg_3_5_inst : DFF_X1 port map( D => mux_out_7_5_port, CK => CLOCK, Q 
                           => pipe1_3_5_port, QN => n_1261);
   pipe1_reg_3_4_inst : DFF_X1 port map( D => mux_out_7_4_port, CK => CLOCK, Q 
                           => pipe1_3_4_port, QN => n_1262);
   pipe1_reg_3_3_inst : DFF_X1 port map( D => mux_out_7_3_port, CK => CLOCK, Q 
                           => pipe1_3_3_port, QN => n_1263);
   pipe1_reg_3_2_inst : DFF_X1 port map( D => mux_out_7_2_port, CK => CLOCK, Q 
                           => pipe1_3_2_port, QN => n_1264);
   pipe1_reg_3_1_inst : DFF_X1 port map( D => mux_out_7_1_port, CK => CLOCK, Q 
                           => pipe1_3_1_port, QN => n_1265);
   pipe1_reg_3_0_inst : DFF_X1 port map( D => mux_out_7_0_port, CK => CLOCK, Q 
                           => pipe1_3_0_port, QN => n_1266);
   pipe1_reg_2_31_inst : DFF_X1 port map( D => mux_out_6_31_port, CK => CLOCK, 
                           Q => pipe1_2_31_port, QN => n_1267);
   pipe1_reg_2_30_inst : DFF_X1 port map( D => mux_out_6_30_port, CK => CLOCK, 
                           Q => pipe1_2_30_port, QN => n_1268);
   pipe1_reg_2_29_inst : DFF_X1 port map( D => mux_out_6_29_port, CK => CLOCK, 
                           Q => pipe1_2_29_port, QN => n_1269);
   pipe1_reg_2_28_inst : DFF_X1 port map( D => mux_out_6_28_port, CK => CLOCK, 
                           Q => pipe1_2_28_port, QN => n_1270);
   pipe1_reg_2_27_inst : DFF_X1 port map( D => mux_out_6_27_port, CK => CLOCK, 
                           Q => pipe1_2_27_port, QN => n_1271);
   pipe1_reg_2_26_inst : DFF_X1 port map( D => mux_out_6_26_port, CK => CLOCK, 
                           Q => pipe1_2_26_port, QN => n_1272);
   pipe1_reg_2_25_inst : DFF_X1 port map( D => mux_out_6_25_port, CK => CLOCK, 
                           Q => pipe1_2_25_port, QN => n_1273);
   pipe1_reg_2_24_inst : DFF_X1 port map( D => mux_out_6_24_port, CK => CLOCK, 
                           Q => pipe1_2_24_port, QN => n_1274);
   pipe1_reg_2_23_inst : DFF_X1 port map( D => mux_out_6_23_port, CK => CLOCK, 
                           Q => pipe1_2_23_port, QN => n_1275);
   pipe1_reg_2_22_inst : DFF_X1 port map( D => mux_out_6_22_port, CK => CLOCK, 
                           Q => pipe1_2_22_port, QN => n_1276);
   pipe1_reg_2_21_inst : DFF_X1 port map( D => mux_out_6_21_port, CK => CLOCK, 
                           Q => pipe1_2_21_port, QN => n_1277);
   pipe1_reg_2_20_inst : DFF_X1 port map( D => mux_out_6_20_port, CK => CLOCK, 
                           Q => pipe1_2_20_port, QN => n_1278);
   pipe1_reg_2_19_inst : DFF_X1 port map( D => mux_out_6_19_port, CK => CLOCK, 
                           Q => pipe1_2_19_port, QN => n_1279);
   pipe1_reg_2_18_inst : DFF_X1 port map( D => mux_out_6_18_port, CK => CLOCK, 
                           Q => pipe1_2_18_port, QN => n_1280);
   pipe1_reg_2_17_inst : DFF_X1 port map( D => mux_out_6_17_port, CK => CLOCK, 
                           Q => pipe1_2_17_port, QN => n_1281);
   pipe1_reg_2_16_inst : DFF_X1 port map( D => mux_out_6_16_port, CK => CLOCK, 
                           Q => pipe1_2_16_port, QN => n_1282);
   pipe1_reg_2_15_inst : DFF_X1 port map( D => mux_out_6_15_port, CK => CLOCK, 
                           Q => pipe1_2_15_port, QN => n_1283);
   pipe1_reg_2_14_inst : DFF_X1 port map( D => mux_out_6_14_port, CK => CLOCK, 
                           Q => pipe1_2_14_port, QN => n_1284);
   pipe1_reg_2_13_inst : DFF_X1 port map( D => mux_out_6_13_port, CK => CLOCK, 
                           Q => pipe1_2_13_port, QN => n_1285);
   pipe1_reg_2_12_inst : DFF_X1 port map( D => mux_out_6_12_port, CK => CLOCK, 
                           Q => pipe1_2_12_port, QN => n_1286);
   pipe1_reg_2_11_inst : DFF_X1 port map( D => mux_out_6_11_port, CK => CLOCK, 
                           Q => pipe1_2_11_port, QN => n_1287);
   pipe1_reg_2_10_inst : DFF_X1 port map( D => mux_out_6_10_port, CK => CLOCK, 
                           Q => pipe1_2_10_port, QN => n_1288);
   pipe1_reg_2_9_inst : DFF_X1 port map( D => mux_out_6_9_port, CK => CLOCK, Q 
                           => pipe1_2_9_port, QN => n_1289);
   pipe1_reg_2_8_inst : DFF_X1 port map( D => mux_out_6_8_port, CK => CLOCK, Q 
                           => pipe1_2_8_port, QN => n_1290);
   pipe1_reg_2_7_inst : DFF_X1 port map( D => mux_out_6_7_port, CK => CLOCK, Q 
                           => pipe1_2_7_port, QN => n_1291);
   pipe1_reg_2_6_inst : DFF_X1 port map( D => mux_out_6_6_port, CK => CLOCK, Q 
                           => pipe1_2_6_port, QN => n_1292);
   pipe1_reg_2_5_inst : DFF_X1 port map( D => mux_out_6_5_port, CK => CLOCK, Q 
                           => pipe1_2_5_port, QN => n_1293);
   pipe1_reg_2_4_inst : DFF_X1 port map( D => mux_out_6_4_port, CK => CLOCK, Q 
                           => pipe1_2_4_port, QN => n_1294);
   pipe1_reg_2_3_inst : DFF_X1 port map( D => mux_out_6_3_port, CK => CLOCK, Q 
                           => pipe1_2_3_port, QN => n_1295);
   pipe1_reg_2_2_inst : DFF_X1 port map( D => mux_out_6_2_port, CK => CLOCK, Q 
                           => pipe1_2_2_port, QN => n_1296);
   pipe1_reg_2_1_inst : DFF_X1 port map( D => mux_out_6_1_port, CK => CLOCK, Q 
                           => pipe1_2_1_port, QN => n_1297);
   pipe1_reg_2_0_inst : DFF_X1 port map( D => mux_out_6_0_port, CK => CLOCK, Q 
                           => pipe1_2_0_port, QN => n_1298);
   pipe1_reg_1_31_inst : DFF_X1 port map( D => mux_out_5_31_port, CK => CLOCK, 
                           Q => pipe1_1_31_port, QN => n_1299);
   addends_reg_5_31_inst : DFF_X1 port map( D => pipe1_1_31_port, CK => CLOCK, 
                           Q => addends_5_31_port, QN => n_1300);
   pipe1_reg_1_30_inst : DFF_X1 port map( D => mux_out_5_30_port, CK => CLOCK, 
                           Q => pipe1_1_30_port, QN => n_1301);
   addends_reg_5_30_inst : DFF_X1 port map( D => pipe1_1_30_port, CK => CLOCK, 
                           Q => addends_5_30_port, QN => n_1302);
   pipe1_reg_1_29_inst : DFF_X1 port map( D => mux_out_5_29_port, CK => CLOCK, 
                           Q => pipe1_1_29_port, QN => n_1303);
   addends_reg_5_29_inst : DFF_X1 port map( D => pipe1_1_29_port, CK => CLOCK, 
                           Q => addends_5_29_port, QN => n_1304);
   pipe1_reg_1_28_inst : DFF_X1 port map( D => mux_out_5_28_port, CK => CLOCK, 
                           Q => pipe1_1_28_port, QN => n_1305);
   addends_reg_5_28_inst : DFF_X1 port map( D => pipe1_1_28_port, CK => CLOCK, 
                           Q => addends_5_28_port, QN => n_1306);
   pipe1_reg_1_27_inst : DFF_X1 port map( D => mux_out_5_27_port, CK => CLOCK, 
                           Q => pipe1_1_27_port, QN => n_1307);
   addends_reg_5_27_inst : DFF_X1 port map( D => pipe1_1_27_port, CK => CLOCK, 
                           Q => addends_5_27_port, QN => n_1308);
   pipe1_reg_1_26_inst : DFF_X1 port map( D => mux_out_5_26_port, CK => CLOCK, 
                           Q => pipe1_1_26_port, QN => n_1309);
   addends_reg_5_26_inst : DFF_X1 port map( D => pipe1_1_26_port, CK => CLOCK, 
                           Q => addends_5_26_port, QN => n_1310);
   pipe1_reg_1_25_inst : DFF_X1 port map( D => mux_out_5_25_port, CK => CLOCK, 
                           Q => pipe1_1_25_port, QN => n_1311);
   addends_reg_5_25_inst : DFF_X1 port map( D => pipe1_1_25_port, CK => CLOCK, 
                           Q => addends_5_25_port, QN => n_1312);
   pipe1_reg_1_24_inst : DFF_X1 port map( D => mux_out_5_24_port, CK => CLOCK, 
                           Q => pipe1_1_24_port, QN => n_1313);
   addends_reg_5_24_inst : DFF_X1 port map( D => pipe1_1_24_port, CK => CLOCK, 
                           Q => addends_5_24_port, QN => n_1314);
   pipe1_reg_1_23_inst : DFF_X1 port map( D => mux_out_5_23_port, CK => CLOCK, 
                           Q => pipe1_1_23_port, QN => n_1315);
   addends_reg_5_23_inst : DFF_X1 port map( D => pipe1_1_23_port, CK => CLOCK, 
                           Q => addends_5_23_port, QN => n_1316);
   pipe1_reg_1_22_inst : DFF_X1 port map( D => mux_out_5_22_port, CK => CLOCK, 
                           Q => pipe1_1_22_port, QN => n_1317);
   addends_reg_5_22_inst : DFF_X1 port map( D => pipe1_1_22_port, CK => CLOCK, 
                           Q => addends_5_22_port, QN => n_1318);
   pipe1_reg_1_21_inst : DFF_X1 port map( D => mux_out_5_21_port, CK => CLOCK, 
                           Q => pipe1_1_21_port, QN => n_1319);
   addends_reg_5_21_inst : DFF_X1 port map( D => pipe1_1_21_port, CK => CLOCK, 
                           Q => addends_5_21_port, QN => n_1320);
   pipe1_reg_1_20_inst : DFF_X1 port map( D => mux_out_5_20_port, CK => CLOCK, 
                           Q => pipe1_1_20_port, QN => n_1321);
   addends_reg_5_20_inst : DFF_X1 port map( D => pipe1_1_20_port, CK => CLOCK, 
                           Q => addends_5_20_port, QN => n_1322);
   pipe1_reg_1_19_inst : DFF_X1 port map( D => mux_out_5_19_port, CK => CLOCK, 
                           Q => pipe1_1_19_port, QN => n_1323);
   addends_reg_5_19_inst : DFF_X1 port map( D => pipe1_1_19_port, CK => CLOCK, 
                           Q => addends_5_19_port, QN => n_1324);
   pipe1_reg_1_18_inst : DFF_X1 port map( D => mux_out_5_18_port, CK => CLOCK, 
                           Q => pipe1_1_18_port, QN => n_1325);
   addends_reg_5_18_inst : DFF_X1 port map( D => pipe1_1_18_port, CK => CLOCK, 
                           Q => addends_5_18_port, QN => n_1326);
   pipe1_reg_1_17_inst : DFF_X1 port map( D => mux_out_5_17_port, CK => CLOCK, 
                           Q => pipe1_1_17_port, QN => n_1327);
   addends_reg_5_17_inst : DFF_X1 port map( D => pipe1_1_17_port, CK => CLOCK, 
                           Q => addends_5_17_port, QN => n_1328);
   pipe1_reg_1_16_inst : DFF_X1 port map( D => mux_out_5_16_port, CK => CLOCK, 
                           Q => pipe1_1_16_port, QN => n_1329);
   addends_reg_5_16_inst : DFF_X1 port map( D => pipe1_1_16_port, CK => CLOCK, 
                           Q => addends_5_16_port, QN => n_1330);
   pipe1_reg_1_15_inst : DFF_X1 port map( D => mux_out_5_15_port, CK => CLOCK, 
                           Q => pipe1_1_15_port, QN => n_1331);
   addends_reg_5_15_inst : DFF_X1 port map( D => pipe1_1_15_port, CK => CLOCK, 
                           Q => addends_5_15_port, QN => n_1332);
   pipe1_reg_1_14_inst : DFF_X1 port map( D => mux_out_5_14_port, CK => CLOCK, 
                           Q => pipe1_1_14_port, QN => n_1333);
   addends_reg_5_14_inst : DFF_X1 port map( D => pipe1_1_14_port, CK => CLOCK, 
                           Q => addends_5_14_port, QN => n_1334);
   pipe1_reg_1_13_inst : DFF_X1 port map( D => mux_out_5_13_port, CK => CLOCK, 
                           Q => pipe1_1_13_port, QN => n_1335);
   addends_reg_5_13_inst : DFF_X1 port map( D => pipe1_1_13_port, CK => CLOCK, 
                           Q => addends_5_13_port, QN => n_1336);
   pipe1_reg_1_12_inst : DFF_X1 port map( D => mux_out_5_12_port, CK => CLOCK, 
                           Q => pipe1_1_12_port, QN => n_1337);
   addends_reg_5_12_inst : DFF_X1 port map( D => pipe1_1_12_port, CK => CLOCK, 
                           Q => addends_5_12_port, QN => n_1338);
   pipe1_reg_1_11_inst : DFF_X1 port map( D => mux_out_5_11_port, CK => CLOCK, 
                           Q => pipe1_1_11_port, QN => n_1339);
   addends_reg_5_11_inst : DFF_X1 port map( D => pipe1_1_11_port, CK => CLOCK, 
                           Q => addends_5_11_port, QN => n_1340);
   pipe1_reg_1_10_inst : DFF_X1 port map( D => mux_out_5_10_port, CK => CLOCK, 
                           Q => pipe1_1_10_port, QN => n_1341);
   addends_reg_5_10_inst : DFF_X1 port map( D => pipe1_1_10_port, CK => CLOCK, 
                           Q => addends_5_10_port, QN => n_1342);
   pipe1_reg_1_9_inst : DFF_X1 port map( D => mux_out_5_9_port, CK => CLOCK, Q 
                           => pipe1_1_9_port, QN => n_1343);
   addends_reg_5_9_inst : DFF_X1 port map( D => pipe1_1_9_port, CK => CLOCK, Q 
                           => addends_5_9_port, QN => n_1344);
   pipe1_reg_1_8_inst : DFF_X1 port map( D => mux_out_5_8_port, CK => CLOCK, Q 
                           => pipe1_1_8_port, QN => n_1345);
   addends_reg_5_8_inst : DFF_X1 port map( D => pipe1_1_8_port, CK => CLOCK, Q 
                           => addends_5_8_port, QN => n_1346);
   pipe1_reg_1_7_inst : DFF_X1 port map( D => mux_out_5_7_port, CK => CLOCK, Q 
                           => pipe1_1_7_port, QN => n_1347);
   addends_reg_5_7_inst : DFF_X1 port map( D => pipe1_1_7_port, CK => CLOCK, Q 
                           => addends_5_7_port, QN => n_1348);
   pipe1_reg_1_6_inst : DFF_X1 port map( D => mux_out_5_6_port, CK => CLOCK, Q 
                           => pipe1_1_6_port, QN => n_1349);
   addends_reg_5_6_inst : DFF_X1 port map( D => pipe1_1_6_port, CK => CLOCK, Q 
                           => addends_5_6_port, QN => n_1350);
   pipe1_reg_1_5_inst : DFF_X1 port map( D => mux_out_5_5_port, CK => CLOCK, Q 
                           => pipe1_1_5_port, QN => n_1351);
   addends_reg_5_5_inst : DFF_X1 port map( D => pipe1_1_5_port, CK => CLOCK, Q 
                           => addends_5_5_port, QN => n_1352);
   pipe1_reg_1_4_inst : DFF_X1 port map( D => mux_out_5_4_port, CK => CLOCK, Q 
                           => pipe1_1_4_port, QN => n_1353);
   addends_reg_5_4_inst : DFF_X1 port map( D => pipe1_1_4_port, CK => CLOCK, Q 
                           => addends_5_4_port, QN => n_1354);
   pipe1_reg_1_3_inst : DFF_X1 port map( D => mux_out_5_3_port, CK => CLOCK, Q 
                           => pipe1_1_3_port, QN => n_1355);
   addends_reg_5_3_inst : DFF_X1 port map( D => pipe1_1_3_port, CK => CLOCK, Q 
                           => addends_5_3_port, QN => n_1356);
   pipe1_reg_1_2_inst : DFF_X1 port map( D => mux_out_5_2_port, CK => CLOCK, Q 
                           => pipe1_1_2_port, QN => n_1357);
   addends_reg_5_2_inst : DFF_X1 port map( D => pipe1_1_2_port, CK => CLOCK, Q 
                           => addends_5_2_port, QN => n_1358);
   pipe1_reg_1_1_inst : DFF_X1 port map( D => mux_out_5_1_port, CK => CLOCK, Q 
                           => pipe1_1_1_port, QN => n_1359);
   addends_reg_5_1_inst : DFF_X1 port map( D => pipe1_1_1_port, CK => CLOCK, Q 
                           => addends_5_1_port, QN => n_1360);
   pipe1_reg_1_0_inst : DFF_X1 port map( D => mux_out_5_0_port, CK => CLOCK, Q 
                           => pipe1_1_0_port, QN => n_1361);
   addends_reg_5_0_inst : DFF_X1 port map( D => pipe1_1_0_port, CK => CLOCK, Q 
                           => addends_5_0_port, QN => n_1362);
   pipe1_reg_0_31_inst : DFF_X1 port map( D => mux_out_4_31_port, CK => CLOCK, 
                           Q => pipe1_0_31_port, QN => n_1363);
   addends_reg_4_31_inst : DFF_X1 port map( D => pipe1_0_31_port, CK => CLOCK, 
                           Q => addends_4_31_port, QN => n_1364);
   pipe1_reg_0_30_inst : DFF_X1 port map( D => mux_out_4_30_port, CK => CLOCK, 
                           Q => pipe1_0_30_port, QN => n_1365);
   addends_reg_4_30_inst : DFF_X1 port map( D => pipe1_0_30_port, CK => CLOCK, 
                           Q => addends_4_30_port, QN => n_1366);
   pipe1_reg_0_29_inst : DFF_X1 port map( D => mux_out_4_29_port, CK => CLOCK, 
                           Q => pipe1_0_29_port, QN => n_1367);
   addends_reg_4_29_inst : DFF_X1 port map( D => pipe1_0_29_port, CK => CLOCK, 
                           Q => addends_4_29_port, QN => n_1368);
   pipe1_reg_0_28_inst : DFF_X1 port map( D => mux_out_4_28_port, CK => CLOCK, 
                           Q => pipe1_0_28_port, QN => n_1369);
   addends_reg_4_28_inst : DFF_X1 port map( D => pipe1_0_28_port, CK => CLOCK, 
                           Q => addends_4_28_port, QN => n_1370);
   pipe1_reg_0_27_inst : DFF_X1 port map( D => mux_out_4_27_port, CK => CLOCK, 
                           Q => pipe1_0_27_port, QN => n_1371);
   addends_reg_4_27_inst : DFF_X1 port map( D => pipe1_0_27_port, CK => CLOCK, 
                           Q => addends_4_27_port, QN => n_1372);
   pipe1_reg_0_26_inst : DFF_X1 port map( D => mux_out_4_26_port, CK => CLOCK, 
                           Q => pipe1_0_26_port, QN => n_1373);
   addends_reg_4_26_inst : DFF_X1 port map( D => pipe1_0_26_port, CK => CLOCK, 
                           Q => addends_4_26_port, QN => n_1374);
   pipe1_reg_0_25_inst : DFF_X1 port map( D => mux_out_4_25_port, CK => CLOCK, 
                           Q => pipe1_0_25_port, QN => n_1375);
   addends_reg_4_25_inst : DFF_X1 port map( D => pipe1_0_25_port, CK => CLOCK, 
                           Q => addends_4_25_port, QN => n_1376);
   pipe1_reg_0_24_inst : DFF_X1 port map( D => mux_out_4_24_port, CK => CLOCK, 
                           Q => pipe1_0_24_port, QN => n_1377);
   addends_reg_4_24_inst : DFF_X1 port map( D => pipe1_0_24_port, CK => CLOCK, 
                           Q => addends_4_24_port, QN => n_1378);
   pipe1_reg_0_23_inst : DFF_X1 port map( D => mux_out_4_23_port, CK => CLOCK, 
                           Q => pipe1_0_23_port, QN => n_1379);
   addends_reg_4_23_inst : DFF_X1 port map( D => pipe1_0_23_port, CK => CLOCK, 
                           Q => addends_4_23_port, QN => n_1380);
   pipe1_reg_0_22_inst : DFF_X1 port map( D => mux_out_4_22_port, CK => CLOCK, 
                           Q => pipe1_0_22_port, QN => n_1381);
   addends_reg_4_22_inst : DFF_X1 port map( D => pipe1_0_22_port, CK => CLOCK, 
                           Q => addends_4_22_port, QN => n_1382);
   pipe1_reg_0_21_inst : DFF_X1 port map( D => mux_out_4_21_port, CK => CLOCK, 
                           Q => pipe1_0_21_port, QN => n_1383);
   addends_reg_4_21_inst : DFF_X1 port map( D => pipe1_0_21_port, CK => CLOCK, 
                           Q => addends_4_21_port, QN => n_1384);
   pipe1_reg_0_20_inst : DFF_X1 port map( D => mux_out_4_20_port, CK => CLOCK, 
                           Q => pipe1_0_20_port, QN => n_1385);
   addends_reg_4_20_inst : DFF_X1 port map( D => pipe1_0_20_port, CK => CLOCK, 
                           Q => addends_4_20_port, QN => n_1386);
   pipe1_reg_0_19_inst : DFF_X1 port map( D => mux_out_4_19_port, CK => CLOCK, 
                           Q => pipe1_0_19_port, QN => n_1387);
   addends_reg_4_19_inst : DFF_X1 port map( D => pipe1_0_19_port, CK => CLOCK, 
                           Q => addends_4_19_port, QN => n_1388);
   pipe1_reg_0_18_inst : DFF_X1 port map( D => mux_out_4_18_port, CK => CLOCK, 
                           Q => pipe1_0_18_port, QN => n_1389);
   addends_reg_4_18_inst : DFF_X1 port map( D => pipe1_0_18_port, CK => CLOCK, 
                           Q => addends_4_18_port, QN => n_1390);
   pipe1_reg_0_17_inst : DFF_X1 port map( D => mux_out_4_17_port, CK => CLOCK, 
                           Q => pipe1_0_17_port, QN => n_1391);
   addends_reg_4_17_inst : DFF_X1 port map( D => pipe1_0_17_port, CK => CLOCK, 
                           Q => addends_4_17_port, QN => n_1392);
   pipe1_reg_0_16_inst : DFF_X1 port map( D => mux_out_4_16_port, CK => CLOCK, 
                           Q => pipe1_0_16_port, QN => n_1393);
   addends_reg_4_16_inst : DFF_X1 port map( D => pipe1_0_16_port, CK => CLOCK, 
                           Q => addends_4_16_port, QN => n_1394);
   pipe1_reg_0_15_inst : DFF_X1 port map( D => mux_out_4_15_port, CK => CLOCK, 
                           Q => pipe1_0_15_port, QN => n_1395);
   addends_reg_4_15_inst : DFF_X1 port map( D => pipe1_0_15_port, CK => CLOCK, 
                           Q => addends_4_15_port, QN => n_1396);
   pipe1_reg_0_14_inst : DFF_X1 port map( D => mux_out_4_14_port, CK => CLOCK, 
                           Q => pipe1_0_14_port, QN => n_1397);
   addends_reg_4_14_inst : DFF_X1 port map( D => pipe1_0_14_port, CK => CLOCK, 
                           Q => addends_4_14_port, QN => n_1398);
   pipe1_reg_0_13_inst : DFF_X1 port map( D => mux_out_4_13_port, CK => CLOCK, 
                           Q => pipe1_0_13_port, QN => n_1399);
   addends_reg_4_13_inst : DFF_X1 port map( D => pipe1_0_13_port, CK => CLOCK, 
                           Q => addends_4_13_port, QN => n_1400);
   pipe1_reg_0_12_inst : DFF_X1 port map( D => mux_out_4_12_port, CK => CLOCK, 
                           Q => pipe1_0_12_port, QN => n_1401);
   addends_reg_4_12_inst : DFF_X1 port map( D => pipe1_0_12_port, CK => CLOCK, 
                           Q => addends_4_12_port, QN => n_1402);
   pipe1_reg_0_11_inst : DFF_X1 port map( D => mux_out_4_11_port, CK => CLOCK, 
                           Q => pipe1_0_11_port, QN => n_1403);
   addends_reg_4_11_inst : DFF_X1 port map( D => pipe1_0_11_port, CK => CLOCK, 
                           Q => addends_4_11_port, QN => n_1404);
   pipe1_reg_0_10_inst : DFF_X1 port map( D => mux_out_4_10_port, CK => CLOCK, 
                           Q => pipe1_0_10_port, QN => n_1405);
   addends_reg_4_10_inst : DFF_X1 port map( D => pipe1_0_10_port, CK => CLOCK, 
                           Q => addends_4_10_port, QN => n_1406);
   pipe1_reg_0_9_inst : DFF_X1 port map( D => mux_out_4_9_port, CK => CLOCK, Q 
                           => pipe1_0_9_port, QN => n_1407);
   addends_reg_4_9_inst : DFF_X1 port map( D => pipe1_0_9_port, CK => CLOCK, Q 
                           => addends_4_9_port, QN => n_1408);
   pipe1_reg_0_8_inst : DFF_X1 port map( D => mux_out_4_8_port, CK => CLOCK, Q 
                           => pipe1_0_8_port, QN => n_1409);
   addends_reg_4_8_inst : DFF_X1 port map( D => pipe1_0_8_port, CK => CLOCK, Q 
                           => addends_4_8_port, QN => n_1410);
   pipe1_reg_0_7_inst : DFF_X1 port map( D => mux_out_4_7_port, CK => CLOCK, Q 
                           => pipe1_0_7_port, QN => n_1411);
   addends_reg_4_7_inst : DFF_X1 port map( D => pipe1_0_7_port, CK => CLOCK, Q 
                           => addends_4_7_port, QN => n_1412);
   pipe1_reg_0_6_inst : DFF_X1 port map( D => mux_out_4_6_port, CK => CLOCK, Q 
                           => pipe1_0_6_port, QN => n_1413);
   addends_reg_4_6_inst : DFF_X1 port map( D => pipe1_0_6_port, CK => CLOCK, Q 
                           => addends_4_6_port, QN => n_1414);
   pipe1_reg_0_5_inst : DFF_X1 port map( D => mux_out_4_5_port, CK => CLOCK, Q 
                           => pipe1_0_5_port, QN => n_1415);
   addends_reg_4_5_inst : DFF_X1 port map( D => pipe1_0_5_port, CK => CLOCK, Q 
                           => addends_4_5_port, QN => n_1416);
   pipe1_reg_0_4_inst : DFF_X1 port map( D => mux_out_4_4_port, CK => CLOCK, Q 
                           => pipe1_0_4_port, QN => n_1417);
   addends_reg_4_4_inst : DFF_X1 port map( D => pipe1_0_4_port, CK => CLOCK, Q 
                           => addends_4_4_port, QN => n_1418);
   pipe1_reg_0_3_inst : DFF_X1 port map( D => mux_out_4_3_port, CK => CLOCK, Q 
                           => pipe1_0_3_port, QN => n_1419);
   addends_reg_4_3_inst : DFF_X1 port map( D => pipe1_0_3_port, CK => CLOCK, Q 
                           => addends_4_3_port, QN => n_1420);
   pipe1_reg_0_2_inst : DFF_X1 port map( D => mux_out_4_2_port, CK => CLOCK, Q 
                           => pipe1_0_2_port, QN => n_1421);
   addends_reg_4_2_inst : DFF_X1 port map( D => pipe1_0_2_port, CK => CLOCK, Q 
                           => addends_4_2_port, QN => n_1422);
   pipe1_reg_0_1_inst : DFF_X1 port map( D => mux_out_4_1_port, CK => CLOCK, Q 
                           => pipe1_0_1_port, QN => n_1423);
   addends_reg_4_1_inst : DFF_X1 port map( D => pipe1_0_1_port, CK => CLOCK, Q 
                           => addends_4_1_port, QN => n_1424);
   pipe1_reg_0_0_inst : DFF_X1 port map( D => mux_out_4_0_port, CK => CLOCK, Q 
                           => pipe1_0_0_port, QN => n_1425);
   pipe2_reg_1_31_inst : DFF_X1 port map( D => pipe1_3_31_port, CK => CLOCK, Q 
                           => pipe2_1_31_port, QN => n_1426);
   addends_reg_7_31_inst : DFF_X1 port map( D => pipe2_1_31_port, CK => CLOCK, 
                           Q => addends_7_31_port, QN => n_1427);
   pipe2_reg_1_30_inst : DFF_X1 port map( D => pipe1_3_30_port, CK => CLOCK, Q 
                           => pipe2_1_30_port, QN => n_1428);
   addends_reg_7_30_inst : DFF_X1 port map( D => pipe2_1_30_port, CK => CLOCK, 
                           Q => addends_7_30_port, QN => n_1429);
   pipe2_reg_1_29_inst : DFF_X1 port map( D => pipe1_3_29_port, CK => CLOCK, Q 
                           => pipe2_1_29_port, QN => n_1430);
   addends_reg_7_29_inst : DFF_X1 port map( D => pipe2_1_29_port, CK => CLOCK, 
                           Q => addends_7_29_port, QN => n_1431);
   pipe2_reg_1_28_inst : DFF_X1 port map( D => pipe1_3_28_port, CK => CLOCK, Q 
                           => pipe2_1_28_port, QN => n_1432);
   addends_reg_7_28_inst : DFF_X1 port map( D => pipe2_1_28_port, CK => CLOCK, 
                           Q => addends_7_28_port, QN => n_1433);
   pipe2_reg_1_27_inst : DFF_X1 port map( D => pipe1_3_27_port, CK => CLOCK, Q 
                           => pipe2_1_27_port, QN => n_1434);
   addends_reg_7_27_inst : DFF_X1 port map( D => pipe2_1_27_port, CK => CLOCK, 
                           Q => addends_7_27_port, QN => n_1435);
   pipe2_reg_1_26_inst : DFF_X1 port map( D => pipe1_3_26_port, CK => CLOCK, Q 
                           => pipe2_1_26_port, QN => n_1436);
   addends_reg_7_26_inst : DFF_X1 port map( D => pipe2_1_26_port, CK => CLOCK, 
                           Q => addends_7_26_port, QN => n_1437);
   pipe2_reg_1_25_inst : DFF_X1 port map( D => pipe1_3_25_port, CK => CLOCK, Q 
                           => pipe2_1_25_port, QN => n_1438);
   addends_reg_7_25_inst : DFF_X1 port map( D => pipe2_1_25_port, CK => CLOCK, 
                           Q => addends_7_25_port, QN => n_1439);
   pipe2_reg_1_24_inst : DFF_X1 port map( D => pipe1_3_24_port, CK => CLOCK, Q 
                           => pipe2_1_24_port, QN => n_1440);
   addends_reg_7_24_inst : DFF_X1 port map( D => pipe2_1_24_port, CK => CLOCK, 
                           Q => addends_7_24_port, QN => n_1441);
   pipe2_reg_1_23_inst : DFF_X1 port map( D => pipe1_3_23_port, CK => CLOCK, Q 
                           => pipe2_1_23_port, QN => n_1442);
   addends_reg_7_23_inst : DFF_X1 port map( D => pipe2_1_23_port, CK => CLOCK, 
                           Q => addends_7_23_port, QN => n_1443);
   pipe2_reg_1_22_inst : DFF_X1 port map( D => pipe1_3_22_port, CK => CLOCK, Q 
                           => pipe2_1_22_port, QN => n_1444);
   addends_reg_7_22_inst : DFF_X1 port map( D => pipe2_1_22_port, CK => CLOCK, 
                           Q => addends_7_22_port, QN => n_1445);
   pipe2_reg_1_21_inst : DFF_X1 port map( D => pipe1_3_21_port, CK => CLOCK, Q 
                           => pipe2_1_21_port, QN => n_1446);
   addends_reg_7_21_inst : DFF_X1 port map( D => pipe2_1_21_port, CK => CLOCK, 
                           Q => addends_7_21_port, QN => n_1447);
   pipe2_reg_1_20_inst : DFF_X1 port map( D => pipe1_3_20_port, CK => CLOCK, Q 
                           => pipe2_1_20_port, QN => n_1448);
   addends_reg_7_20_inst : DFF_X1 port map( D => pipe2_1_20_port, CK => CLOCK, 
                           Q => addends_7_20_port, QN => n_1449);
   pipe2_reg_1_19_inst : DFF_X1 port map( D => pipe1_3_19_port, CK => CLOCK, Q 
                           => pipe2_1_19_port, QN => n_1450);
   addends_reg_7_19_inst : DFF_X1 port map( D => pipe2_1_19_port, CK => CLOCK, 
                           Q => addends_7_19_port, QN => n_1451);
   pipe2_reg_1_18_inst : DFF_X1 port map( D => pipe1_3_18_port, CK => CLOCK, Q 
                           => pipe2_1_18_port, QN => n_1452);
   addends_reg_7_18_inst : DFF_X1 port map( D => pipe2_1_18_port, CK => CLOCK, 
                           Q => addends_7_18_port, QN => n_1453);
   pipe2_reg_1_17_inst : DFF_X1 port map( D => pipe1_3_17_port, CK => CLOCK, Q 
                           => pipe2_1_17_port, QN => n_1454);
   addends_reg_7_17_inst : DFF_X1 port map( D => pipe2_1_17_port, CK => CLOCK, 
                           Q => addends_7_17_port, QN => n_1455);
   pipe2_reg_1_16_inst : DFF_X1 port map( D => pipe1_3_16_port, CK => CLOCK, Q 
                           => pipe2_1_16_port, QN => n_1456);
   addends_reg_7_16_inst : DFF_X1 port map( D => pipe2_1_16_port, CK => CLOCK, 
                           Q => addends_7_16_port, QN => n_1457);
   pipe2_reg_1_15_inst : DFF_X1 port map( D => pipe1_3_15_port, CK => CLOCK, Q 
                           => pipe2_1_15_port, QN => n_1458);
   addends_reg_7_15_inst : DFF_X1 port map( D => pipe2_1_15_port, CK => CLOCK, 
                           Q => addends_7_15_port, QN => n_1459);
   pipe2_reg_1_14_inst : DFF_X1 port map( D => pipe1_3_14_port, CK => CLOCK, Q 
                           => pipe2_1_14_port, QN => n_1460);
   addends_reg_7_14_inst : DFF_X1 port map( D => pipe2_1_14_port, CK => CLOCK, 
                           Q => addends_7_14_port, QN => n_1461);
   pipe2_reg_1_13_inst : DFF_X1 port map( D => pipe1_3_13_port, CK => CLOCK, Q 
                           => pipe2_1_13_port, QN => n_1462);
   addends_reg_7_13_inst : DFF_X1 port map( D => pipe2_1_13_port, CK => CLOCK, 
                           Q => addends_7_13_port, QN => n_1463);
   pipe2_reg_1_12_inst : DFF_X1 port map( D => pipe1_3_12_port, CK => CLOCK, Q 
                           => pipe2_1_12_port, QN => n_1464);
   addends_reg_7_12_inst : DFF_X1 port map( D => pipe2_1_12_port, CK => CLOCK, 
                           Q => addends_7_12_port, QN => n_1465);
   pipe2_reg_1_11_inst : DFF_X1 port map( D => pipe1_3_11_port, CK => CLOCK, Q 
                           => pipe2_1_11_port, QN => n_1466);
   addends_reg_7_11_inst : DFF_X1 port map( D => pipe2_1_11_port, CK => CLOCK, 
                           Q => addends_7_11_port, QN => n_1467);
   pipe2_reg_1_10_inst : DFF_X1 port map( D => pipe1_3_10_port, CK => CLOCK, Q 
                           => pipe2_1_10_port, QN => n_1468);
   addends_reg_7_10_inst : DFF_X1 port map( D => pipe2_1_10_port, CK => CLOCK, 
                           Q => addends_7_10_port, QN => n_1469);
   pipe2_reg_1_9_inst : DFF_X1 port map( D => pipe1_3_9_port, CK => CLOCK, Q =>
                           pipe2_1_9_port, QN => n_1470);
   addends_reg_7_9_inst : DFF_X1 port map( D => pipe2_1_9_port, CK => CLOCK, Q 
                           => addends_7_9_port, QN => n_1471);
   pipe2_reg_1_8_inst : DFF_X1 port map( D => pipe1_3_8_port, CK => CLOCK, Q =>
                           pipe2_1_8_port, QN => n_1472);
   addends_reg_7_8_inst : DFF_X1 port map( D => pipe2_1_8_port, CK => CLOCK, Q 
                           => addends_7_8_port, QN => n_1473);
   pipe2_reg_1_7_inst : DFF_X1 port map( D => pipe1_3_7_port, CK => CLOCK, Q =>
                           pipe2_1_7_port, QN => n_1474);
   addends_reg_7_7_inst : DFF_X1 port map( D => pipe2_1_7_port, CK => CLOCK, Q 
                           => addends_7_7_port, QN => n_1475);
   pipe2_reg_1_6_inst : DFF_X1 port map( D => pipe1_3_6_port, CK => CLOCK, Q =>
                           pipe2_1_6_port, QN => n_1476);
   addends_reg_7_6_inst : DFF_X1 port map( D => pipe2_1_6_port, CK => CLOCK, Q 
                           => addends_7_6_port, QN => n_1477);
   pipe2_reg_1_5_inst : DFF_X1 port map( D => pipe1_3_5_port, CK => CLOCK, Q =>
                           pipe2_1_5_port, QN => n_1478);
   addends_reg_7_5_inst : DFF_X1 port map( D => pipe2_1_5_port, CK => CLOCK, Q 
                           => addends_7_5_port, QN => n_1479);
   pipe2_reg_1_4_inst : DFF_X1 port map( D => pipe1_3_4_port, CK => CLOCK, Q =>
                           pipe2_1_4_port, QN => n_1480);
   addends_reg_7_4_inst : DFF_X1 port map( D => pipe2_1_4_port, CK => CLOCK, Q 
                           => addends_7_4_port, QN => n_1481);
   pipe2_reg_1_3_inst : DFF_X1 port map( D => pipe1_3_3_port, CK => CLOCK, Q =>
                           pipe2_1_3_port, QN => n_1482);
   addends_reg_7_3_inst : DFF_X1 port map( D => pipe2_1_3_port, CK => CLOCK, Q 
                           => addends_7_3_port, QN => n_1483);
   pipe2_reg_1_2_inst : DFF_X1 port map( D => pipe1_3_2_port, CK => CLOCK, Q =>
                           pipe2_1_2_port, QN => n_1484);
   addends_reg_7_2_inst : DFF_X1 port map( D => pipe2_1_2_port, CK => CLOCK, Q 
                           => addends_7_2_port, QN => n_1485);
   pipe2_reg_1_1_inst : DFF_X1 port map( D => pipe1_3_1_port, CK => CLOCK, Q =>
                           pipe2_1_1_port, QN => n_1486);
   addends_reg_7_1_inst : DFF_X1 port map( D => pipe2_1_1_port, CK => CLOCK, Q 
                           => addends_7_1_port, QN => n_1487);
   pipe2_reg_1_0_inst : DFF_X1 port map( D => pipe1_3_0_port, CK => CLOCK, Q =>
                           pipe2_1_0_port, QN => n_1488);
   addends_reg_7_0_inst : DFF_X1 port map( D => pipe2_1_0_port, CK => CLOCK, Q 
                           => addends_7_0_port, QN => n_1489);
   pipe2_reg_0_31_inst : DFF_X1 port map( D => pipe1_2_31_port, CK => CLOCK, Q 
                           => pipe2_0_31_port, QN => n_1490);
   addends_reg_6_31_inst : DFF_X1 port map( D => pipe2_0_31_port, CK => CLOCK, 
                           Q => addends_6_31_port, QN => n_1491);
   pipe2_reg_0_30_inst : DFF_X1 port map( D => pipe1_2_30_port, CK => CLOCK, Q 
                           => pipe2_0_30_port, QN => n_1492);
   addends_reg_6_30_inst : DFF_X1 port map( D => pipe2_0_30_port, CK => CLOCK, 
                           Q => addends_6_30_port, QN => n_1493);
   pipe2_reg_0_29_inst : DFF_X1 port map( D => pipe1_2_29_port, CK => CLOCK, Q 
                           => pipe2_0_29_port, QN => n_1494);
   addends_reg_6_29_inst : DFF_X1 port map( D => pipe2_0_29_port, CK => CLOCK, 
                           Q => addends_6_29_port, QN => n_1495);
   pipe2_reg_0_28_inst : DFF_X1 port map( D => pipe1_2_28_port, CK => CLOCK, Q 
                           => pipe2_0_28_port, QN => n_1496);
   addends_reg_6_28_inst : DFF_X1 port map( D => pipe2_0_28_port, CK => CLOCK, 
                           Q => addends_6_28_port, QN => n_1497);
   pipe2_reg_0_27_inst : DFF_X1 port map( D => pipe1_2_27_port, CK => CLOCK, Q 
                           => pipe2_0_27_port, QN => n_1498);
   addends_reg_6_27_inst : DFF_X1 port map( D => pipe2_0_27_port, CK => CLOCK, 
                           Q => addends_6_27_port, QN => n_1499);
   pipe2_reg_0_26_inst : DFF_X1 port map( D => pipe1_2_26_port, CK => CLOCK, Q 
                           => pipe2_0_26_port, QN => n_1500);
   addends_reg_6_26_inst : DFF_X1 port map( D => pipe2_0_26_port, CK => CLOCK, 
                           Q => addends_6_26_port, QN => n_1501);
   pipe2_reg_0_25_inst : DFF_X1 port map( D => pipe1_2_25_port, CK => CLOCK, Q 
                           => pipe2_0_25_port, QN => n_1502);
   addends_reg_6_25_inst : DFF_X1 port map( D => pipe2_0_25_port, CK => CLOCK, 
                           Q => addends_6_25_port, QN => n_1503);
   pipe2_reg_0_24_inst : DFF_X1 port map( D => pipe1_2_24_port, CK => CLOCK, Q 
                           => pipe2_0_24_port, QN => n_1504);
   addends_reg_6_24_inst : DFF_X1 port map( D => pipe2_0_24_port, CK => CLOCK, 
                           Q => addends_6_24_port, QN => n_1505);
   pipe2_reg_0_23_inst : DFF_X1 port map( D => pipe1_2_23_port, CK => CLOCK, Q 
                           => pipe2_0_23_port, QN => n_1506);
   addends_reg_6_23_inst : DFF_X1 port map( D => pipe2_0_23_port, CK => CLOCK, 
                           Q => addends_6_23_port, QN => n_1507);
   pipe2_reg_0_22_inst : DFF_X1 port map( D => pipe1_2_22_port, CK => CLOCK, Q 
                           => pipe2_0_22_port, QN => n_1508);
   addends_reg_6_22_inst : DFF_X1 port map( D => pipe2_0_22_port, CK => CLOCK, 
                           Q => addends_6_22_port, QN => n_1509);
   pipe2_reg_0_21_inst : DFF_X1 port map( D => pipe1_2_21_port, CK => CLOCK, Q 
                           => pipe2_0_21_port, QN => n_1510);
   addends_reg_6_21_inst : DFF_X1 port map( D => pipe2_0_21_port, CK => CLOCK, 
                           Q => addends_6_21_port, QN => n_1511);
   pipe2_reg_0_20_inst : DFF_X1 port map( D => pipe1_2_20_port, CK => CLOCK, Q 
                           => pipe2_0_20_port, QN => n_1512);
   addends_reg_6_20_inst : DFF_X1 port map( D => pipe2_0_20_port, CK => CLOCK, 
                           Q => addends_6_20_port, QN => n_1513);
   pipe2_reg_0_19_inst : DFF_X1 port map( D => pipe1_2_19_port, CK => CLOCK, Q 
                           => pipe2_0_19_port, QN => n_1514);
   addends_reg_6_19_inst : DFF_X1 port map( D => pipe2_0_19_port, CK => CLOCK, 
                           Q => addends_6_19_port, QN => n_1515);
   pipe2_reg_0_18_inst : DFF_X1 port map( D => pipe1_2_18_port, CK => CLOCK, Q 
                           => pipe2_0_18_port, QN => n_1516);
   addends_reg_6_18_inst : DFF_X1 port map( D => pipe2_0_18_port, CK => CLOCK, 
                           Q => addends_6_18_port, QN => n_1517);
   pipe2_reg_0_17_inst : DFF_X1 port map( D => pipe1_2_17_port, CK => CLOCK, Q 
                           => pipe2_0_17_port, QN => n_1518);
   addends_reg_6_17_inst : DFF_X1 port map( D => pipe2_0_17_port, CK => CLOCK, 
                           Q => addends_6_17_port, QN => n_1519);
   pipe2_reg_0_16_inst : DFF_X1 port map( D => pipe1_2_16_port, CK => CLOCK, Q 
                           => pipe2_0_16_port, QN => n_1520);
   addends_reg_6_16_inst : DFF_X1 port map( D => pipe2_0_16_port, CK => CLOCK, 
                           Q => addends_6_16_port, QN => n_1521);
   pipe2_reg_0_15_inst : DFF_X1 port map( D => pipe1_2_15_port, CK => CLOCK, Q 
                           => pipe2_0_15_port, QN => n_1522);
   addends_reg_6_15_inst : DFF_X1 port map( D => pipe2_0_15_port, CK => CLOCK, 
                           Q => addends_6_15_port, QN => n_1523);
   pipe2_reg_0_14_inst : DFF_X1 port map( D => pipe1_2_14_port, CK => CLOCK, Q 
                           => pipe2_0_14_port, QN => n_1524);
   addends_reg_6_14_inst : DFF_X1 port map( D => pipe2_0_14_port, CK => CLOCK, 
                           Q => addends_6_14_port, QN => n_1525);
   pipe2_reg_0_13_inst : DFF_X1 port map( D => pipe1_2_13_port, CK => CLOCK, Q 
                           => pipe2_0_13_port, QN => n_1526);
   addends_reg_6_13_inst : DFF_X1 port map( D => pipe2_0_13_port, CK => CLOCK, 
                           Q => addends_6_13_port, QN => n_1527);
   pipe2_reg_0_12_inst : DFF_X1 port map( D => pipe1_2_12_port, CK => CLOCK, Q 
                           => pipe2_0_12_port, QN => n_1528);
   addends_reg_6_12_inst : DFF_X1 port map( D => pipe2_0_12_port, CK => CLOCK, 
                           Q => addends_6_12_port, QN => n_1529);
   pipe2_reg_0_11_inst : DFF_X1 port map( D => pipe1_2_11_port, CK => CLOCK, Q 
                           => pipe2_0_11_port, QN => n_1530);
   addends_reg_6_11_inst : DFF_X1 port map( D => pipe2_0_11_port, CK => CLOCK, 
                           Q => addends_6_11_port, QN => n_1531);
   pipe2_reg_0_10_inst : DFF_X1 port map( D => pipe1_2_10_port, CK => CLOCK, Q 
                           => pipe2_0_10_port, QN => n_1532);
   addends_reg_6_10_inst : DFF_X1 port map( D => pipe2_0_10_port, CK => CLOCK, 
                           Q => addends_6_10_port, QN => n_1533);
   pipe2_reg_0_9_inst : DFF_X1 port map( D => pipe1_2_9_port, CK => CLOCK, Q =>
                           pipe2_0_9_port, QN => n_1534);
   addends_reg_6_9_inst : DFF_X1 port map( D => pipe2_0_9_port, CK => CLOCK, Q 
                           => addends_6_9_port, QN => n_1535);
   pipe2_reg_0_8_inst : DFF_X1 port map( D => pipe1_2_8_port, CK => CLOCK, Q =>
                           pipe2_0_8_port, QN => n_1536);
   addends_reg_6_8_inst : DFF_X1 port map( D => pipe2_0_8_port, CK => CLOCK, Q 
                           => addends_6_8_port, QN => n_1537);
   pipe2_reg_0_7_inst : DFF_X1 port map( D => pipe1_2_7_port, CK => CLOCK, Q =>
                           pipe2_0_7_port, QN => n_1538);
   addends_reg_6_7_inst : DFF_X1 port map( D => pipe2_0_7_port, CK => CLOCK, Q 
                           => addends_6_7_port, QN => n_1539);
   pipe2_reg_0_6_inst : DFF_X1 port map( D => pipe1_2_6_port, CK => CLOCK, Q =>
                           pipe2_0_6_port, QN => n_1540);
   addends_reg_6_6_inst : DFF_X1 port map( D => pipe2_0_6_port, CK => CLOCK, Q 
                           => addends_6_6_port, QN => n_1541);
   pipe2_reg_0_5_inst : DFF_X1 port map( D => pipe1_2_5_port, CK => CLOCK, Q =>
                           pipe2_0_5_port, QN => n_1542);
   addends_reg_6_5_inst : DFF_X1 port map( D => pipe2_0_5_port, CK => CLOCK, Q 
                           => addends_6_5_port, QN => n_1543);
   pipe2_reg_0_4_inst : DFF_X1 port map( D => pipe1_2_4_port, CK => CLOCK, Q =>
                           pipe2_0_4_port, QN => n_1544);
   addends_reg_6_4_inst : DFF_X1 port map( D => pipe2_0_4_port, CK => CLOCK, Q 
                           => addends_6_4_port, QN => n_1545);
   pipe2_reg_0_3_inst : DFF_X1 port map( D => pipe1_2_3_port, CK => CLOCK, Q =>
                           pipe2_0_3_port, QN => n_1546);
   pipe2_reg_0_2_inst : DFF_X1 port map( D => pipe1_2_2_port, CK => CLOCK, Q =>
                           pipe2_0_2_port, QN => n_1547);
   pipe2_reg_0_1_inst : DFF_X1 port map( D => pipe1_2_1_port, CK => CLOCK, Q =>
                           pipe2_0_1_port, QN => n_1548);
   pipe2_reg_0_0_inst : DFF_X1 port map( D => pipe1_2_0_port, CK => CLOCK, Q =>
                           pipe2_0_0_port, QN => n_1549);
   enc_1 : ENCODER_0 port map( INPUT(2) => B(1), INPUT(1) => B(0), INPUT(0) => 
                           X_Logic0_port, OUTPUT(2) => selector_2_port, 
                           OUTPUT(1) => selector_1_port, OUTPUT(0) => 
                           selector_0_port);
   enc_2 : ENCODER_7 port map( INPUT(2) => B(3), INPUT(1) => B(2), INPUT(0) => 
                           B(1), OUTPUT(2) => selector_5_port, OUTPUT(1) => 
                           selector_4_port, OUTPUT(0) => selector_3_port);
   enc_3 : ENCODER_6 port map( INPUT(2) => B(5), INPUT(1) => B(4), INPUT(0) => 
                           B(3), OUTPUT(2) => selector_8_port, OUTPUT(1) => 
                           selector_7_port, OUTPUT(0) => selector_6_port);
   enc_4 : ENCODER_5 port map( INPUT(2) => B(7), INPUT(1) => B(6), INPUT(0) => 
                           B(5), OUTPUT(2) => selector_11_port, OUTPUT(1) => 
                           selector_10_port, OUTPUT(0) => selector_9_port);
   enc_5 : ENCODER_4 port map( INPUT(2) => B(9), INPUT(1) => B(8), INPUT(0) => 
                           B(7), OUTPUT(2) => selector_14_port, OUTPUT(1) => 
                           selector_13_port, OUTPUT(0) => selector_12_port);
   enc_6 : ENCODER_3 port map( INPUT(2) => B(11), INPUT(1) => B(10), INPUT(0) 
                           => B(9), OUTPUT(2) => selector_17_port, OUTPUT(1) =>
                           selector_16_port, OUTPUT(0) => selector_15_port);
   enc_7 : ENCODER_2 port map( INPUT(2) => B(13), INPUT(1) => B(12), INPUT(0) 
                           => B(11), OUTPUT(2) => selector_20_port, OUTPUT(1) 
                           => selector_19_port, OUTPUT(0) => selector_18_port);
   enc_8 : ENCODER_1 port map( INPUT(2) => B(15), INPUT(1) => B(14), INPUT(0) 
                           => B(13), OUTPUT(2) => selector_23_port, OUTPUT(1) 
                           => selector_22_port, OUTPUT(0) => selector_21_port);
   MUX_I_0 : MUX5to1_NBIT32_8 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => A(15), B(14) => A(14), B(13)
                           => A(13), B(12) => A(12), B(11) => A(11), B(10) => 
                           A(10), B(9) => A(9), B(8) => A(8), B(7) => A(7), 
                           B(6) => A(6), B(5) => A(5), B(4) => A(4), B(3) => 
                           A(3), B(2) => A(2), B(1) => A(1), B(0) => n20, C(31)
                           => n6, C(30) => n6, C(29) => n6, C(28) => n6, C(27) 
                           => n6, C(26) => n6, C(25) => n6, C(24) => n6, C(23) 
                           => n6, C(22) => n6, C(21) => n6, C(20) => n6, C(19) 
                           => n6, C(18) => n6, C(17) => n6, C(16) => n6, C(15) 
                           => A_neg_0_15_port, C(14) => A_neg_0_14_port, C(13) 
                           => A_neg_0_13_port, C(12) => A_neg_0_12_port, C(11) 
                           => A_neg_0_11_port, C(10) => A_neg_0_10_port, C(9) 
                           => A_neg_0_9_port, C(8) => A_neg_0_8_port, C(7) => 
                           A_neg_0_7_port, C(6) => A_neg_0_6_port, C(5) => 
                           A_neg_0_5_port, C(4) => A_neg_0_4_port, C(3) => 
                           A_neg_0_3_port, C(2) => A_neg_0_2_port, C(1) => 
                           A_neg_0_1_port, C(0) => n20, D(31) => X_Logic0_port,
                           D(30) => X_Logic0_port, D(29) => X_Logic0_port, 
                           D(28) => X_Logic0_port, D(27) => X_Logic0_port, 
                           D(26) => X_Logic0_port, D(25) => X_Logic0_port, 
                           D(24) => X_Logic0_port, D(23) => X_Logic0_port, 
                           D(22) => X_Logic0_port, D(21) => X_Logic0_port, 
                           D(20) => X_Logic0_port, D(19) => X_Logic0_port, 
                           D(18) => X_Logic0_port, D(17) => X_Logic0_port, 
                           D(16) => A(15), D(15) => A(14), D(14) => A(13), 
                           D(13) => A(12), D(12) => A(11), D(11) => A(10), 
                           D(10) => A(9), D(9) => A(8), D(8) => A(7), D(7) => 
                           A(6), D(6) => A(5), D(5) => A(4), D(4) => A(3), D(3)
                           => A(2), D(2) => A(1), D(1) => A(0), D(0) => 
                           X_Logic0_port, E(31) => n8, E(30) => n8, E(29) => n8
                           , E(28) => n8, E(27) => n8, E(26) => n8, E(25) => n8
                           , E(24) => n8, E(23) => n8, E(22) => n8, E(21) => n8
                           , E(20) => n8, E(19) => n8, E(18) => n8, E(17) => n8
                           , E(16) => A_neg_1_16_port, E(15) => A_neg_1_15_port
                           , E(14) => A_neg_1_14_port, E(13) => A_neg_1_13_port
                           , E(12) => A_neg_1_12_port, E(11) => A_neg_1_11_port
                           , E(10) => A_neg_1_10_port, E(9) => A_neg_1_9_port, 
                           E(8) => A_neg_1_8_port, E(7) => A_neg_1_7_port, E(6)
                           => A_neg_1_6_port, E(5) => A_neg_1_5_port, E(4) => 
                           A_neg_1_4_port, E(3) => A_neg_1_3_port, E(2) => 
                           A_neg_1_2_port, E(1) => A(0), E(0) => n69, SEL(2) =>
                           selector_2_port, SEL(1) => selector_1_port, SEL(0) 
                           => selector_0_port, Y(31) => addends_0_31_port, 
                           Y(30) => addends_0_30_port, Y(29) => 
                           addends_0_29_port, Y(28) => addends_0_28_port, Y(27)
                           => addends_0_27_port, Y(26) => addends_0_26_port, 
                           Y(25) => addends_0_25_port, Y(24) => 
                           addends_0_24_port, Y(23) => addends_0_23_port, Y(22)
                           => addends_0_22_port, Y(21) => addends_0_21_port, 
                           Y(20) => addends_0_20_port, Y(19) => 
                           addends_0_19_port, Y(18) => addends_0_18_port, Y(17)
                           => addends_0_17_port, Y(16) => addends_0_16_port, 
                           Y(15) => addends_0_15_port, Y(14) => 
                           addends_0_14_port, Y(13) => addends_0_13_port, Y(12)
                           => addends_0_12_port, Y(11) => addends_0_11_port, 
                           Y(10) => addends_0_10_port, Y(9) => addends_0_9_port
                           , Y(8) => addends_0_8_port, Y(7) => addends_0_7_port
                           , Y(6) => addends_0_6_port, Y(5) => addends_0_5_port
                           , Y(4) => addends_0_4_port, Y(3) => addends_0_3_port
                           , Y(2) => addends_0_2_port, Y(1) => addends_0_1_port
                           , Y(0) => addends_0_0_port);
   MUX_I_1 : MUX5to1_NBIT32_7 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => A(15), B(16) => A(14), B(15)
                           => A(13), B(14) => A(12), B(13) => A(11), B(12) => 
                           A(10), B(11) => A(9), B(10) => A(8), B(9) => A(7), 
                           B(8) => A(6), B(7) => A(5), B(6) => A(4), B(5) => 
                           A(3), B(4) => A(2), B(3) => A(1), B(2) => A(0), B(1)
                           => X_Logic0_port, B(0) => X_Logic0_port, C(31) => n9
                           , C(30) => n9, C(29) => n9, C(28) => n9, C(27) => n9
                           , C(26) => n9, C(25) => n9, C(24) => n9, C(23) => n9
                           , C(22) => n9, C(21) => n9, C(20) => n9, C(19) => n9
                           , C(18) => n9, C(17) => A_neg_2_17_port, C(16) => 
                           A_neg_2_16_port, C(15) => A_neg_2_15_port, C(14) => 
                           A_neg_2_14_port, C(13) => A_neg_2_13_port, C(12) => 
                           A_neg_2_12_port, C(11) => A_neg_2_11_port, C(10) => 
                           A_neg_2_10_port, C(9) => A_neg_2_9_port, C(8) => 
                           A_neg_2_8_port, C(7) => A_neg_2_7_port, C(6) => 
                           A_neg_2_6_port, C(5) => A_neg_2_5_port, C(4) => 
                           A_neg_2_4_port, C(3) => A_neg_2_3_port, C(2) => n20,
                           C(1) => n69, C(0) => n69, D(31) => X_Logic0_port, 
                           D(30) => X_Logic0_port, D(29) => X_Logic0_port, 
                           D(28) => X_Logic0_port, D(27) => X_Logic0_port, 
                           D(26) => X_Logic0_port, D(25) => X_Logic0_port, 
                           D(24) => X_Logic0_port, D(23) => X_Logic0_port, 
                           D(22) => X_Logic0_port, D(21) => X_Logic0_port, 
                           D(20) => X_Logic0_port, D(19) => X_Logic0_port, 
                           D(18) => A(15), D(17) => A(14), D(16) => A(13), 
                           D(15) => A(12), D(14) => A(11), D(13) => A(10), 
                           D(12) => A(9), D(11) => A(8), D(10) => A(7), D(9) =>
                           A(6), D(8) => A(5), D(7) => A(4), D(6) => A(3), D(5)
                           => A(2), D(4) => A(1), D(3) => A(0), D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n11, E(30) => n11, E(29) => 
                           n11, E(28) => n11, E(27) => n11, E(26) => n11, E(25)
                           => n11, E(24) => n11, E(23) => n11, E(22) => n11, 
                           E(21) => n11, E(20) => n11, E(19) => n11, E(18) => 
                           A_neg_3_18_port, E(17) => A_neg_3_17_port, E(16) => 
                           A_neg_3_16_port, E(15) => A_neg_3_15_port, E(14) => 
                           A_neg_3_14_port, E(13) => A_neg_3_13_port, E(12) => 
                           A_neg_3_12_port, E(11) => A_neg_3_11_port, E(10) => 
                           A_neg_3_10_port, E(9) => A_neg_3_9_port, E(8) => 
                           A_neg_3_8_port, E(7) => A_neg_3_7_port, E(6) => 
                           A_neg_3_6_port, E(5) => A_neg_3_5_port, E(4) => 
                           A_neg_3_4_port, E(3) => A(0), E(2) => n69, E(1) => 
                           n69, E(0) => n69, SEL(2) => selector_5_port, SEL(1) 
                           => selector_4_port, SEL(0) => selector_3_port, Y(31)
                           => addends_1_31_port, Y(30) => addends_1_30_port, 
                           Y(29) => addends_1_29_port, Y(28) => 
                           addends_1_28_port, Y(27) => addends_1_27_port, Y(26)
                           => addends_1_26_port, Y(25) => addends_1_25_port, 
                           Y(24) => addends_1_24_port, Y(23) => 
                           addends_1_23_port, Y(22) => addends_1_22_port, Y(21)
                           => addends_1_21_port, Y(20) => addends_1_20_port, 
                           Y(19) => addends_1_19_port, Y(18) => 
                           addends_1_18_port, Y(17) => addends_1_17_port, Y(16)
                           => addends_1_16_port, Y(15) => addends_1_15_port, 
                           Y(14) => addends_1_14_port, Y(13) => 
                           addends_1_13_port, Y(12) => addends_1_12_port, Y(11)
                           => addends_1_11_port, Y(10) => addends_1_10_port, 
                           Y(9) => addends_1_9_port, Y(8) => addends_1_8_port, 
                           Y(7) => addends_1_7_port, Y(6) => addends_1_6_port, 
                           Y(5) => addends_1_5_port, Y(4) => addends_1_4_port, 
                           Y(3) => addends_1_3_port, Y(2) => addends_1_2_port, 
                           Y(1) => addends_1_1_port, Y(0) => addends_1_0_port);
   MUX_I_2 : MUX5to1_NBIT32_6 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => A(15), B(18) => A(14), B(17)
                           => A(13), B(16) => A(12), B(15) => A(11), B(14) => 
                           A(10), B(13) => A(9), B(12) => A(8), B(11) => A(7), 
                           B(10) => A(6), B(9) => A(5), B(8) => A(4), B(7) => 
                           A(3), B(6) => A(2), B(5) => A(1), B(4) => A(0), B(3)
                           => X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n2, 
                           C(30) => n2, C(29) => n2, C(28) => n2, C(27) => n2, 
                           C(26) => n2, C(25) => n2, C(24) => n2, C(23) => n2, 
                           C(22) => n2, C(21) => n2, C(20) => n2, C(19) => 
                           A_neg_4_19_port, C(18) => A_neg_4_18_port, C(17) => 
                           A_neg_4_17_port, C(16) => A_neg_4_16_port, C(15) => 
                           A_neg_4_15_port, C(14) => A_neg_4_14_port, C(13) => 
                           A_neg_4_13_port, C(12) => A_neg_4_12_port, C(11) => 
                           A_neg_4_11_port, C(10) => A_neg_4_10_port, C(9) => 
                           A_neg_4_9_port, C(8) => A_neg_4_8_port, C(7) => 
                           A_neg_4_7_port, C(6) => A_neg_4_6_port, C(5) => 
                           A_neg_4_5_port, C(4) => n20, C(3) => n69, C(2) => 
                           n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => A(15), D(19) => A(14), D(18)
                           => A(13), D(17) => A(12), D(16) => A(11), D(15) => 
                           A(10), D(14) => A(9), D(13) => A(8), D(12) => A(7), 
                           D(11) => A(6), D(10) => A(5), D(9) => A(4), D(8) => 
                           A(3), D(7) => A(2), D(6) => A(1), D(5) => A(0), D(4)
                           => X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n3, E(30) => n3, E(29) => n3
                           , E(28) => n3, E(27) => n3, E(26) => n3, E(25) => n3
                           , E(24) => n3, E(23) => n3, E(22) => n3, E(21) => n3
                           , E(20) => A_neg_5_20_port, E(19) => A_neg_5_19_port
                           , E(18) => A_neg_5_18_port, E(17) => A_neg_5_17_port
                           , E(16) => A_neg_5_16_port, E(15) => A_neg_5_15_port
                           , E(14) => A_neg_5_14_port, E(13) => A_neg_5_13_port
                           , E(12) => A_neg_5_12_port, E(11) => A_neg_5_11_port
                           , E(10) => A_neg_5_10_port, E(9) => A_neg_5_9_port, 
                           E(8) => A_neg_5_8_port, E(7) => A_neg_5_7_port, E(6)
                           => A_neg_5_6_port, E(5) => A(0), E(4) => n69, E(3) 
                           => n69, E(2) => n69, E(1) => n69, E(0) => n69, 
                           SEL(2) => selector_8_port, SEL(1) => selector_7_port
                           , SEL(0) => selector_6_port, Y(31) => 
                           mux_out_2_31_port, Y(30) => mux_out_2_30_port, Y(29)
                           => mux_out_2_29_port, Y(28) => mux_out_2_28_port, 
                           Y(27) => mux_out_2_27_port, Y(26) => 
                           mux_out_2_26_port, Y(25) => mux_out_2_25_port, Y(24)
                           => mux_out_2_24_port, Y(23) => mux_out_2_23_port, 
                           Y(22) => mux_out_2_22_port, Y(21) => 
                           mux_out_2_21_port, Y(20) => mux_out_2_20_port, Y(19)
                           => mux_out_2_19_port, Y(18) => mux_out_2_18_port, 
                           Y(17) => mux_out_2_17_port, Y(16) => 
                           mux_out_2_16_port, Y(15) => mux_out_2_15_port, Y(14)
                           => mux_out_2_14_port, Y(13) => mux_out_2_13_port, 
                           Y(12) => mux_out_2_12_port, Y(11) => 
                           mux_out_2_11_port, Y(10) => mux_out_2_10_port, Y(9) 
                           => mux_out_2_9_port, Y(8) => mux_out_2_8_port, Y(7) 
                           => mux_out_2_7_port, Y(6) => mux_out_2_6_port, Y(5) 
                           => mux_out_2_5_port, Y(4) => mux_out_2_4_port, Y(3) 
                           => mux_out_2_3_port, Y(2) => mux_out_2_2_port, Y(1) 
                           => mux_out_2_1_port, Y(0) => mux_out_2_0_port);
   MUX_I_3 : MUX5to1_NBIT32_5 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => A(15), B(20) => A(14), B(19)
                           => A(13), B(18) => A(12), B(17) => A(11), B(16) => 
                           A(10), B(15) => A(9), B(14) => A(8), B(13) => A(7), 
                           B(12) => A(6), B(11) => A(5), B(10) => A(4), B(9) =>
                           A(3), B(8) => A(2), B(7) => A(1), B(6) => n20, B(5) 
                           => X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n4, 
                           C(30) => n4, C(29) => n4, C(28) => n4, C(27) => n4, 
                           C(26) => n4, C(25) => n4, C(24) => n4, C(23) => n4, 
                           C(22) => n4, C(21) => A_neg_6_21_port, C(20) => 
                           A_neg_6_20_port, C(19) => A_neg_6_19_port, C(18) => 
                           A_neg_6_18_port, C(17) => A_neg_6_17_port, C(16) => 
                           A_neg_6_16_port, C(15) => A_neg_6_15_port, C(14) => 
                           A_neg_6_14_port, C(13) => A_neg_6_13_port, C(12) => 
                           A_neg_6_12_port, C(11) => A_neg_6_11_port, C(10) => 
                           A_neg_6_10_port, C(9) => A_neg_6_9_port, C(8) => 
                           A_neg_6_8_port, C(7) => A_neg_6_7_port, C(6) => n20,
                           C(5) => n69, C(4) => n69, C(3) => n69, C(2) => n69, 
                           C(1) => n69, C(0) => n69, D(31) => X_Logic0_port, 
                           D(30) => X_Logic0_port, D(29) => X_Logic0_port, 
                           D(28) => X_Logic0_port, D(27) => X_Logic0_port, 
                           D(26) => X_Logic0_port, D(25) => X_Logic0_port, 
                           D(24) => X_Logic0_port, D(23) => X_Logic0_port, 
                           D(22) => A(15), D(21) => A(14), D(20) => A(13), 
                           D(19) => A(12), D(18) => A(11), D(17) => A(10), 
                           D(16) => A(9), D(15) => A(8), D(14) => A(7), D(13) 
                           => A(6), D(12) => A(5), D(11) => A(4), D(10) => A(3)
                           , D(9) => A(2), D(8) => A(1), D(7) => A(0), D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n5, E(30) => n5, E(29) => n5
                           , E(28) => n5, E(27) => n5, E(26) => n5, E(25) => n5
                           , E(24) => n5, E(23) => n5, E(22) => A_neg_7_22_port
                           , E(21) => A_neg_7_21_port, E(20) => A_neg_7_20_port
                           , E(19) => A_neg_7_19_port, E(18) => A_neg_7_18_port
                           , E(17) => A_neg_7_17_port, E(16) => A_neg_7_16_port
                           , E(15) => A_neg_7_15_port, E(14) => A_neg_7_14_port
                           , E(13) => A_neg_7_13_port, E(12) => A_neg_7_12_port
                           , E(11) => A_neg_7_11_port, E(10) => A_neg_7_10_port
                           , E(9) => A_neg_7_9_port, E(8) => A_neg_7_8_port, 
                           E(7) => A(0), E(6) => n69, E(5) => n69, E(4) => n69,
                           E(3) => n69, E(2) => n69, E(1) => n69, E(0) => n69, 
                           SEL(2) => selector_11_port, SEL(1) => 
                           selector_10_port, SEL(0) => selector_9_port, Y(31) 
                           => mux_out_3_31_port, Y(30) => mux_out_3_30_port, 
                           Y(29) => mux_out_3_29_port, Y(28) => 
                           mux_out_3_28_port, Y(27) => mux_out_3_27_port, Y(26)
                           => mux_out_3_26_port, Y(25) => mux_out_3_25_port, 
                           Y(24) => mux_out_3_24_port, Y(23) => 
                           mux_out_3_23_port, Y(22) => mux_out_3_22_port, Y(21)
                           => mux_out_3_21_port, Y(20) => mux_out_3_20_port, 
                           Y(19) => mux_out_3_19_port, Y(18) => 
                           mux_out_3_18_port, Y(17) => mux_out_3_17_port, Y(16)
                           => mux_out_3_16_port, Y(15) => mux_out_3_15_port, 
                           Y(14) => mux_out_3_14_port, Y(13) => 
                           mux_out_3_13_port, Y(12) => mux_out_3_12_port, Y(11)
                           => mux_out_3_11_port, Y(10) => mux_out_3_10_port, 
                           Y(9) => mux_out_3_9_port, Y(8) => mux_out_3_8_port, 
                           Y(7) => mux_out_3_7_port, Y(6) => mux_out_3_6_port, 
                           Y(5) => mux_out_3_5_port, Y(4) => mux_out_3_4_port, 
                           Y(3) => mux_out_3_3_port, Y(2) => mux_out_3_2_port, 
                           Y(1) => mux_out_3_1_port, Y(0) => mux_out_3_0_port);
   MUX_I_4 : MUX5to1_NBIT32_4 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => A(15), B(22) => A(14), B(21)
                           => A(13), B(20) => A(12), B(19) => A(11), B(18) => 
                           A(10), B(17) => A(9), B(16) => A(8), B(15) => A(7), 
                           B(14) => A(6), B(13) => A(5), B(12) => A(4), B(11) 
                           => A(3), B(10) => A(2), B(9) => A(1), B(8) => n20, 
                           B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) 
                           => X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n7, 
                           C(30) => n7, C(29) => n7, C(28) => n7, C(27) => n7, 
                           C(26) => n7, C(25) => n7, C(24) => n7, C(23) => 
                           A_neg_8_23_port, C(22) => A_neg_8_22_port, C(21) => 
                           A_neg_8_21_port, C(20) => A_neg_8_20_port, C(19) => 
                           A_neg_8_19_port, C(18) => A_neg_8_18_port, C(17) => 
                           A_neg_8_17_port, C(16) => A_neg_8_16_port, C(15) => 
                           A_neg_8_15_port, C(14) => A_neg_8_14_port, C(13) => 
                           A_neg_8_13_port, C(12) => A_neg_8_12_port, C(11) => 
                           A_neg_8_11_port, C(10) => A_neg_8_10_port, C(9) => 
                           A_neg_8_9_port, C(8) => n20, C(7) => n69, C(6) => 
                           n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) => 
                           n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => A(15), D(23) => A(14), D(22)
                           => A(13), D(21) => A(12), D(20) => A(11), D(19) => 
                           A(10), D(18) => A(9), D(17) => A(8), D(16) => A(7), 
                           D(15) => A(6), D(14) => A(5), D(13) => A(4), D(12) 
                           => A(3), D(11) => A(2), D(10) => A(1), D(9) => A(0),
                           D(8) => X_Logic0_port, D(7) => X_Logic0_port, D(6) 
                           => X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n10, E(30) => n10, E(29) => 
                           n10, E(28) => n10, E(27) => n10, E(26) => n10, E(25)
                           => n10, E(24) => A_neg_9_24_port, E(23) => 
                           A_neg_9_23_port, E(22) => A_neg_9_22_port, E(21) => 
                           A_neg_9_21_port, E(20) => A_neg_9_20_port, E(19) => 
                           A_neg_9_19_port, E(18) => A_neg_9_18_port, E(17) => 
                           A_neg_9_17_port, E(16) => A_neg_9_16_port, E(15) => 
                           A_neg_9_15_port, E(14) => A_neg_9_14_port, E(13) => 
                           A_neg_9_13_port, E(12) => A_neg_9_12_port, E(11) => 
                           A_neg_9_11_port, E(10) => A_neg_9_10_port, E(9) => 
                           A(0), E(8) => n69, E(7) => n69, E(6) => n69, E(5) =>
                           n69, E(4) => n69, E(3) => n69, E(2) => n69, E(1) => 
                           n69, E(0) => n69, SEL(2) => selector_14_port, SEL(1)
                           => selector_13_port, SEL(0) => selector_12_port, 
                           Y(31) => mux_out_4_31_port, Y(30) => 
                           mux_out_4_30_port, Y(29) => mux_out_4_29_port, Y(28)
                           => mux_out_4_28_port, Y(27) => mux_out_4_27_port, 
                           Y(26) => mux_out_4_26_port, Y(25) => 
                           mux_out_4_25_port, Y(24) => mux_out_4_24_port, Y(23)
                           => mux_out_4_23_port, Y(22) => mux_out_4_22_port, 
                           Y(21) => mux_out_4_21_port, Y(20) => 
                           mux_out_4_20_port, Y(19) => mux_out_4_19_port, Y(18)
                           => mux_out_4_18_port, Y(17) => mux_out_4_17_port, 
                           Y(16) => mux_out_4_16_port, Y(15) => 
                           mux_out_4_15_port, Y(14) => mux_out_4_14_port, Y(13)
                           => mux_out_4_13_port, Y(12) => mux_out_4_12_port, 
                           Y(11) => mux_out_4_11_port, Y(10) => 
                           mux_out_4_10_port, Y(9) => mux_out_4_9_port, Y(8) =>
                           mux_out_4_8_port, Y(7) => mux_out_4_7_port, Y(6) => 
                           mux_out_4_6_port, Y(5) => mux_out_4_5_port, Y(4) => 
                           mux_out_4_4_port, Y(3) => mux_out_4_3_port, Y(2) => 
                           mux_out_4_2_port, Y(1) => mux_out_4_1_port, Y(0) => 
                           mux_out_4_0_port);
   MUX_I_5 : MUX5to1_NBIT32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => A(15), B(24) => A(14), B(23)
                           => A(13), B(22) => A(12), B(21) => A(11), B(20) => 
                           A(10), B(19) => A(9), B(18) => A(8), B(17) => A(7), 
                           B(16) => A(6), B(15) => A(5), B(14) => A(4), B(13) 
                           => A(3), B(12) => A(2), B(11) => A(1), B(10) => n20,
                           B(9) => X_Logic0_port, B(8) => X_Logic0_port, B(7) 
                           => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n12, 
                           C(30) => n12, C(29) => n12, C(28) => n12, C(27) => 
                           n12, C(26) => n12, C(25) => A_neg_10_25_port, C(24) 
                           => A_neg_10_24_port, C(23) => A_neg_10_23_port, 
                           C(22) => A_neg_10_22_port, C(21) => A_neg_10_21_port
                           , C(20) => A_neg_10_20_port, C(19) => 
                           A_neg_10_19_port, C(18) => A_neg_10_18_port, C(17) 
                           => A_neg_10_17_port, C(16) => A_neg_10_16_port, 
                           C(15) => A_neg_10_15_port, C(14) => A_neg_10_14_port
                           , C(13) => A_neg_10_13_port, C(12) => 
                           A_neg_10_12_port, C(11) => A_neg_10_11_port, C(10) 
                           => n20, C(9) => n69, C(8) => n69, C(7) => n69, C(6) 
                           => n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) 
                           => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => A(15), D(25) => A(14), D(24)
                           => A(13), D(23) => A(12), D(22) => A(11), D(21) => 
                           A(10), D(20) => A(9), D(19) => A(8), D(18) => A(7), 
                           D(17) => A(6), D(16) => A(5), D(15) => A(4), D(14) 
                           => A(3), D(13) => A(2), D(12) => A(1), D(11) => A(0)
                           , D(10) => X_Logic0_port, D(9) => X_Logic0_port, 
                           D(8) => X_Logic0_port, D(7) => X_Logic0_port, D(6) 
                           => X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n13, E(30) => n13, E(29) => 
                           n13, E(28) => n13, E(27) => n13, E(26) => 
                           A_neg_11_26_port, E(25) => A_neg_11_25_port, E(24) 
                           => A_neg_11_24_port, E(23) => A_neg_11_23_port, 
                           E(22) => A_neg_11_22_port, E(21) => A_neg_11_21_port
                           , E(20) => A_neg_11_20_port, E(19) => 
                           A_neg_11_19_port, E(18) => A_neg_11_18_port, E(17) 
                           => A_neg_11_17_port, E(16) => A_neg_11_16_port, 
                           E(15) => A_neg_11_15_port, E(14) => A_neg_11_14_port
                           , E(13) => A_neg_11_13_port, E(12) => 
                           A_neg_11_12_port, E(11) => A(0), E(10) => n69, E(9) 
                           => n69, E(8) => n69, E(7) => n69, E(6) => n69, E(5) 
                           => n69, E(4) => n69, E(3) => n69, E(2) => n69, E(1) 
                           => n69, E(0) => n69, SEL(2) => selector_17_port, 
                           SEL(1) => selector_16_port, SEL(0) => 
                           selector_15_port, Y(31) => mux_out_5_31_port, Y(30) 
                           => mux_out_5_30_port, Y(29) => mux_out_5_29_port, 
                           Y(28) => mux_out_5_28_port, Y(27) => 
                           mux_out_5_27_port, Y(26) => mux_out_5_26_port, Y(25)
                           => mux_out_5_25_port, Y(24) => mux_out_5_24_port, 
                           Y(23) => mux_out_5_23_port, Y(22) => 
                           mux_out_5_22_port, Y(21) => mux_out_5_21_port, Y(20)
                           => mux_out_5_20_port, Y(19) => mux_out_5_19_port, 
                           Y(18) => mux_out_5_18_port, Y(17) => 
                           mux_out_5_17_port, Y(16) => mux_out_5_16_port, Y(15)
                           => mux_out_5_15_port, Y(14) => mux_out_5_14_port, 
                           Y(13) => mux_out_5_13_port, Y(12) => 
                           mux_out_5_12_port, Y(11) => mux_out_5_11_port, Y(10)
                           => mux_out_5_10_port, Y(9) => mux_out_5_9_port, Y(8)
                           => mux_out_5_8_port, Y(7) => mux_out_5_7_port, Y(6) 
                           => mux_out_5_6_port, Y(5) => mux_out_5_5_port, Y(4) 
                           => mux_out_5_4_port, Y(3) => mux_out_5_3_port, Y(2) 
                           => mux_out_5_2_port, Y(1) => mux_out_5_1_port, Y(0) 
                           => mux_out_5_0_port);
   MUX_I_6 : MUX5to1_NBIT32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => A(15), B(26) => A(14), B(25)
                           => A(13), B(24) => A(12), B(23) => A(11), B(22) => 
                           A(10), B(21) => A(9), B(20) => A(8), B(19) => A(7), 
                           B(18) => A(6), B(17) => A(5), B(16) => A(4), B(15) 
                           => A(3), B(14) => A(2), B(13) => A(1), B(12) => n20,
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n14, 
                           C(30) => n14, C(29) => n14, C(28) => n14, C(27) => 
                           A_neg_12_27_port, C(26) => A_neg_12_26_port, C(25) 
                           => A_neg_12_25_port, C(24) => A_neg_12_24_port, 
                           C(23) => A_neg_12_23_port, C(22) => A_neg_12_22_port
                           , C(21) => A_neg_12_21_port, C(20) => 
                           A_neg_12_20_port, C(19) => A_neg_12_19_port, C(18) 
                           => A_neg_12_18_port, C(17) => A_neg_12_17_port, 
                           C(16) => A_neg_12_16_port, C(15) => A_neg_12_15_port
                           , C(14) => A_neg_12_14_port, C(13) => 
                           A_neg_12_13_port, C(12) => n20, C(11) => n69, C(10) 
                           => n69, C(9) => n69, C(8) => n69, C(7) => n69, C(6) 
                           => n69, C(5) => n69, C(4) => n69, C(3) => n69, C(2) 
                           => n69, C(1) => n69, C(0) => n69, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => A(15), D(27) => A(14), D(26)
                           => A(13), D(25) => A(12), D(24) => A(11), D(23) => 
                           A(10), D(22) => A(9), D(21) => A(8), D(20) => A(7), 
                           D(19) => A(6), D(18) => A(5), D(17) => A(4), D(16) 
                           => A(3), D(15) => A(2), D(14) => A(1), D(13) => A(0)
                           , D(12) => X_Logic0_port, D(11) => X_Logic0_port, 
                           D(10) => X_Logic0_port, D(9) => X_Logic0_port, D(8) 
                           => X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n15, E(30) => n15, E(29) => 
                           n15, E(28) => A_neg_13_28_port, E(27) => 
                           A_neg_13_27_port, E(26) => A_neg_13_26_port, E(25) 
                           => A_neg_13_25_port, E(24) => A_neg_13_24_port, 
                           E(23) => A_neg_13_23_port, E(22) => A_neg_13_22_port
                           , E(21) => A_neg_13_21_port, E(20) => 
                           A_neg_13_20_port, E(19) => A_neg_13_19_port, E(18) 
                           => A_neg_13_18_port, E(17) => A_neg_13_17_port, 
                           E(16) => A_neg_13_16_port, E(15) => A_neg_13_15_port
                           , E(14) => A_neg_13_14_port, E(13) => n20, E(12) => 
                           n69, E(11) => n69, E(10) => n69, E(9) => n69, E(8) 
                           => n69, E(7) => n69, E(6) => n69, E(5) => n69, E(4) 
                           => n69, E(3) => n69, E(2) => n69, E(1) => n69, E(0) 
                           => n69, SEL(2) => selector_20_port, SEL(1) => 
                           selector_19_port, SEL(0) => selector_18_port, Y(31) 
                           => mux_out_6_31_port, Y(30) => mux_out_6_30_port, 
                           Y(29) => mux_out_6_29_port, Y(28) => 
                           mux_out_6_28_port, Y(27) => mux_out_6_27_port, Y(26)
                           => mux_out_6_26_port, Y(25) => mux_out_6_25_port, 
                           Y(24) => mux_out_6_24_port, Y(23) => 
                           mux_out_6_23_port, Y(22) => mux_out_6_22_port, Y(21)
                           => mux_out_6_21_port, Y(20) => mux_out_6_20_port, 
                           Y(19) => mux_out_6_19_port, Y(18) => 
                           mux_out_6_18_port, Y(17) => mux_out_6_17_port, Y(16)
                           => mux_out_6_16_port, Y(15) => mux_out_6_15_port, 
                           Y(14) => mux_out_6_14_port, Y(13) => 
                           mux_out_6_13_port, Y(12) => mux_out_6_12_port, Y(11)
                           => mux_out_6_11_port, Y(10) => mux_out_6_10_port, 
                           Y(9) => mux_out_6_9_port, Y(8) => mux_out_6_8_port, 
                           Y(7) => mux_out_6_7_port, Y(6) => mux_out_6_6_port, 
                           Y(5) => mux_out_6_5_port, Y(4) => mux_out_6_4_port, 
                           Y(3) => mux_out_6_3_port, Y(2) => mux_out_6_2_port, 
                           Y(1) => mux_out_6_1_port, Y(0) => mux_out_6_0_port);
   MUX_I_7 : MUX5to1_NBIT32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => A(15), B(28) => A(14), B(27)
                           => A(13), B(26) => A(12), B(25) => A(11), B(24) => 
                           A(10), B(23) => A(9), B(22) => A(8), B(21) => A(7), 
                           B(20) => A(6), B(19) => A(5), B(18) => A(4), B(17) 
                           => A(3), B(16) => A(2), B(15) => A(1), B(14) => n20,
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => n16, 
                           C(30) => n16, C(29) => A_neg_14_29_port, C(28) => 
                           A_neg_14_28_port, C(27) => A_neg_14_27_port, C(26) 
                           => A_neg_14_26_port, C(25) => A_neg_14_25_port, 
                           C(24) => A_neg_14_24_port, C(23) => A_neg_14_23_port
                           , C(22) => A_neg_14_22_port, C(21) => 
                           A_neg_14_21_port, C(20) => A_neg_14_20_port, C(19) 
                           => A_neg_14_19_port, C(18) => A_neg_14_18_port, 
                           C(17) => A_neg_14_17_port, C(16) => A_neg_14_16_port
                           , C(15) => A_neg_14_15_port, C(14) => n20, C(13) => 
                           n69, C(12) => n69, C(11) => n69, C(10) => n69, C(9) 
                           => n69, C(8) => n69, C(7) => n69, C(6) => n69, C(5) 
                           => n69, C(4) => n69, C(3) => n69, C(2) => n69, C(1) 
                           => n69, C(0) => n69, D(31) => X_Logic0_port, D(30) 
                           => A(15), D(29) => A(14), D(28) => A(13), D(27) => 
                           A(12), D(26) => A(11), D(25) => A(10), D(24) => A(9)
                           , D(23) => A(8), D(22) => A(7), D(21) => A(6), D(20)
                           => A(5), D(19) => A(4), D(18) => A(3), D(17) => A(2)
                           , D(16) => A(1), D(15) => A(0), D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => n1, E(30) => 
                           A_neg_15_30_port, E(29) => A_neg_15_29_port, E(28) 
                           => A_neg_15_28_port, E(27) => A_neg_15_27_port, 
                           E(26) => A_neg_15_26_port, E(25) => A_neg_15_25_port
                           , E(24) => A_neg_15_24_port, E(23) => 
                           A_neg_15_23_port, E(22) => A_neg_15_22_port, E(21) 
                           => A_neg_15_21_port, E(20) => A_neg_15_20_port, 
                           E(19) => A_neg_15_19_port, E(18) => A_neg_15_18_port
                           , E(17) => A_neg_15_17_port, E(16) => 
                           A_neg_15_16_port, E(15) => n20, E(14) => n69, E(13) 
                           => n69, E(12) => n69, E(11) => n69, E(10) => n69, 
                           E(9) => n69, E(8) => n69, E(7) => n69, E(6) => n69, 
                           E(5) => n69, E(4) => n69, E(3) => n69, E(2) => n69, 
                           E(1) => n69, E(0) => n69, SEL(2) => selector_23_port
                           , SEL(1) => selector_22_port, SEL(0) => 
                           selector_21_port, Y(31) => mux_out_7_31_port, Y(30) 
                           => mux_out_7_30_port, Y(29) => mux_out_7_29_port, 
                           Y(28) => mux_out_7_28_port, Y(27) => 
                           mux_out_7_27_port, Y(26) => mux_out_7_26_port, Y(25)
                           => mux_out_7_25_port, Y(24) => mux_out_7_24_port, 
                           Y(23) => mux_out_7_23_port, Y(22) => 
                           mux_out_7_22_port, Y(21) => mux_out_7_21_port, Y(20)
                           => mux_out_7_20_port, Y(19) => mux_out_7_19_port, 
                           Y(18) => mux_out_7_18_port, Y(17) => 
                           mux_out_7_17_port, Y(16) => mux_out_7_16_port, Y(15)
                           => mux_out_7_15_port, Y(14) => mux_out_7_14_port, 
                           Y(13) => mux_out_7_13_port, Y(12) => 
                           mux_out_7_12_port, Y(11) => mux_out_7_11_port, Y(10)
                           => mux_out_7_10_port, Y(9) => mux_out_7_9_port, Y(8)
                           => mux_out_7_8_port, Y(7) => mux_out_7_7_port, Y(6) 
                           => mux_out_7_6_port, Y(5) => mux_out_7_5_port, Y(4) 
                           => mux_out_7_4_port, Y(3) => mux_out_7_3_port, Y(2) 
                           => mux_out_7_2_port, Y(1) => mux_out_7_1_port, Y(0) 
                           => mux_out_7_0_port);
   ADD0 : ADDER_NBIT32_NBIT_PER_BLOCK4_7 port map( A(31) => addends_0_31_port, 
                           A(30) => addends_0_30_port, A(29) => 
                           addends_0_29_port, A(28) => addends_0_28_port, A(27)
                           => addends_0_27_port, A(26) => addends_0_26_port, 
                           A(25) => addends_0_25_port, A(24) => 
                           addends_0_24_port, A(23) => addends_0_23_port, A(22)
                           => addends_0_22_port, A(21) => addends_0_21_port, 
                           A(20) => addends_0_20_port, A(19) => 
                           addends_0_19_port, A(18) => addends_0_18_port, A(17)
                           => addends_0_17_port, A(16) => addends_0_16_port, 
                           A(15) => addends_0_15_port, A(14) => 
                           addends_0_14_port, A(13) => addends_0_13_port, A(12)
                           => addends_0_12_port, A(11) => addends_0_11_port, 
                           A(10) => addends_0_10_port, A(9) => addends_0_9_port
                           , A(8) => addends_0_8_port, A(7) => addends_0_7_port
                           , A(6) => addends_0_6_port, A(5) => addends_0_5_port
                           , A(4) => addends_0_4_port, A(3) => addends_0_3_port
                           , A(2) => addends_0_2_port, A(1) => addends_0_1_port
                           , A(0) => addends_0_0_port, B(31) => 
                           addends_1_31_port, B(30) => addends_1_30_port, B(29)
                           => addends_1_29_port, B(28) => addends_1_28_port, 
                           B(27) => addends_1_27_port, B(26) => 
                           addends_1_26_port, B(25) => addends_1_25_port, B(24)
                           => addends_1_24_port, B(23) => addends_1_23_port, 
                           B(22) => addends_1_22_port, B(21) => 
                           addends_1_21_port, B(20) => addends_1_20_port, B(19)
                           => addends_1_19_port, B(18) => addends_1_18_port, 
                           B(17) => addends_1_17_port, B(16) => 
                           addends_1_16_port, B(15) => addends_1_15_port, B(14)
                           => addends_1_14_port, B(13) => addends_1_13_port, 
                           B(12) => addends_1_12_port, B(11) => 
                           addends_1_11_port, B(10) => addends_1_10_port, B(9) 
                           => addends_1_9_port, B(8) => addends_1_8_port, B(7) 
                           => addends_1_7_port, B(6) => addends_1_6_port, B(5) 
                           => addends_1_5_port, B(4) => addends_1_4_port, B(3) 
                           => addends_1_3_port, B(2) => addends_1_2_port, B(1) 
                           => addends_1_1_port, B(0) => addends_1_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_0_31_port, S(30) => reg_in_0_30_port
                           , S(29) => reg_in_0_29_port, S(28) => 
                           reg_in_0_28_port, S(27) => reg_in_0_27_port, S(26) 
                           => reg_in_0_26_port, S(25) => reg_in_0_25_port, 
                           S(24) => reg_in_0_24_port, S(23) => reg_in_0_23_port
                           , S(22) => reg_in_0_22_port, S(21) => 
                           reg_in_0_21_port, S(20) => reg_in_0_20_port, S(19) 
                           => reg_in_0_19_port, S(18) => reg_in_0_18_port, 
                           S(17) => reg_in_0_17_port, S(16) => reg_in_0_16_port
                           , S(15) => reg_in_0_15_port, S(14) => 
                           reg_in_0_14_port, S(13) => reg_in_0_13_port, S(12) 
                           => reg_in_0_12_port, S(11) => reg_in_0_11_port, 
                           S(10) => reg_in_0_10_port, S(9) => reg_in_0_9_port, 
                           S(8) => reg_in_0_8_port, S(7) => reg_in_0_7_port, 
                           S(6) => reg_in_0_6_port, S(5) => reg_in_0_5_port, 
                           S(4) => reg_in_0_4_port, S(3) => reg_in_0_3_port, 
                           S(2) => reg_in_0_2_port, S(1) => reg_in_0_1_port, 
                           S(0) => reg_in_0_0_port, Cout => n_1550);
   REG0 : REG_NBIT32_3 port map( clk => CLOCK, reset => X_Logic0_port, enable 
                           => X_Logic1_port, data_in(31) => reg_in_0_31_port, 
                           data_in(30) => reg_in_0_30_port, data_in(29) => 
                           reg_in_0_29_port, data_in(28) => reg_in_0_28_port, 
                           data_in(27) => reg_in_0_27_port, data_in(26) => 
                           reg_in_0_26_port, data_in(25) => reg_in_0_25_port, 
                           data_in(24) => reg_in_0_24_port, data_in(23) => 
                           reg_in_0_23_port, data_in(22) => reg_in_0_22_port, 
                           data_in(21) => reg_in_0_21_port, data_in(20) => 
                           reg_in_0_20_port, data_in(19) => reg_in_0_19_port, 
                           data_in(18) => reg_in_0_18_port, data_in(17) => 
                           reg_in_0_17_port, data_in(16) => reg_in_0_16_port, 
                           data_in(15) => reg_in_0_15_port, data_in(14) => 
                           reg_in_0_14_port, data_in(13) => reg_in_0_13_port, 
                           data_in(12) => reg_in_0_12_port, data_in(11) => 
                           reg_in_0_11_port, data_in(10) => reg_in_0_10_port, 
                           data_in(9) => reg_in_0_9_port, data_in(8) => 
                           reg_in_0_8_port, data_in(7) => reg_in_0_7_port, 
                           data_in(6) => reg_in_0_6_port, data_in(5) => 
                           reg_in_0_5_port, data_in(4) => reg_in_0_4_port, 
                           data_in(3) => reg_in_0_3_port, data_in(2) => 
                           reg_in_0_2_port, data_in(1) => reg_in_0_1_port, 
                           data_in(0) => reg_in_0_0_port, data_out(31) => 
                           reg_out_0_31_port, data_out(30) => reg_out_0_30_port
                           , data_out(29) => reg_out_0_29_port, data_out(28) =>
                           reg_out_0_28_port, data_out(27) => reg_out_0_27_port
                           , data_out(26) => reg_out_0_26_port, data_out(25) =>
                           reg_out_0_25_port, data_out(24) => reg_out_0_24_port
                           , data_out(23) => reg_out_0_23_port, data_out(22) =>
                           reg_out_0_22_port, data_out(21) => reg_out_0_21_port
                           , data_out(20) => reg_out_0_20_port, data_out(19) =>
                           reg_out_0_19_port, data_out(18) => reg_out_0_18_port
                           , data_out(17) => reg_out_0_17_port, data_out(16) =>
                           reg_out_0_16_port, data_out(15) => reg_out_0_15_port
                           , data_out(14) => reg_out_0_14_port, data_out(13) =>
                           reg_out_0_13_port, data_out(12) => reg_out_0_12_port
                           , data_out(11) => reg_out_0_11_port, data_out(10) =>
                           reg_out_0_10_port, data_out(9) => reg_out_0_9_port, 
                           data_out(8) => reg_out_0_8_port, data_out(7) => 
                           reg_out_0_7_port, data_out(6) => reg_out_0_6_port, 
                           data_out(5) => reg_out_0_5_port, data_out(4) => 
                           reg_out_0_4_port, data_out(3) => reg_out_0_3_port, 
                           data_out(2) => reg_out_0_2_port, data_out(1) => 
                           reg_out_0_1_port, data_out(0) => reg_out_0_0_port);
   ADD_0i_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_6 port map( A(31) => 
                           reg_out_0_31_port, A(30) => reg_out_0_30_port, A(29)
                           => reg_out_0_29_port, A(28) => reg_out_0_28_port, 
                           A(27) => reg_out_0_27_port, A(26) => 
                           reg_out_0_26_port, A(25) => reg_out_0_25_port, A(24)
                           => reg_out_0_24_port, A(23) => reg_out_0_23_port, 
                           A(22) => reg_out_0_22_port, A(21) => 
                           reg_out_0_21_port, A(20) => reg_out_0_20_port, A(19)
                           => reg_out_0_19_port, A(18) => reg_out_0_18_port, 
                           A(17) => reg_out_0_17_port, A(16) => 
                           reg_out_0_16_port, A(15) => reg_out_0_15_port, A(14)
                           => reg_out_0_14_port, A(13) => reg_out_0_13_port, 
                           A(12) => reg_out_0_12_port, A(11) => 
                           reg_out_0_11_port, A(10) => reg_out_0_10_port, A(9) 
                           => reg_out_0_9_port, A(8) => reg_out_0_8_port, A(7) 
                           => reg_out_0_7_port, A(6) => reg_out_0_6_port, A(5) 
                           => reg_out_0_5_port, A(4) => reg_out_0_4_port, A(3) 
                           => reg_out_0_3_port, A(2) => reg_out_0_2_port, A(1) 
                           => reg_out_0_1_port, A(0) => reg_out_0_0_port, B(31)
                           => addends_2_31_port, B(30) => addends_2_30_port, 
                           B(29) => addends_2_29_port, B(28) => 
                           addends_2_28_port, B(27) => addends_2_27_port, B(26)
                           => addends_2_26_port, B(25) => addends_2_25_port, 
                           B(24) => addends_2_24_port, B(23) => 
                           addends_2_23_port, B(22) => addends_2_22_port, B(21)
                           => addends_2_21_port, B(20) => addends_2_20_port, 
                           B(19) => addends_2_19_port, B(18) => 
                           addends_2_18_port, B(17) => addends_2_17_port, B(16)
                           => addends_2_16_port, B(15) => addends_2_15_port, 
                           B(14) => addends_2_14_port, B(13) => 
                           addends_2_13_port, B(12) => addends_2_12_port, B(11)
                           => addends_2_11_port, B(10) => addends_2_10_port, 
                           B(9) => addends_2_9_port, B(8) => addends_2_8_port, 
                           B(7) => addends_2_7_port, B(6) => addends_2_6_port, 
                           B(5) => addends_2_5_port, B(4) => addends_2_4_port, 
                           B(3) => addends_2_3_port, B(2) => addends_2_2_port, 
                           B(1) => addends_2_1_port, B(0) => addends_2_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_0_31_port, S(30) => 
                           add_out_0_30_port, S(29) => add_out_0_29_port, S(28)
                           => add_out_0_28_port, S(27) => add_out_0_27_port, 
                           S(26) => add_out_0_26_port, S(25) => 
                           add_out_0_25_port, S(24) => add_out_0_24_port, S(23)
                           => add_out_0_23_port, S(22) => add_out_0_22_port, 
                           S(21) => add_out_0_21_port, S(20) => 
                           add_out_0_20_port, S(19) => add_out_0_19_port, S(18)
                           => add_out_0_18_port, S(17) => add_out_0_17_port, 
                           S(16) => add_out_0_16_port, S(15) => 
                           add_out_0_15_port, S(14) => add_out_0_14_port, S(13)
                           => add_out_0_13_port, S(12) => add_out_0_12_port, 
                           S(11) => add_out_0_11_port, S(10) => 
                           add_out_0_10_port, S(9) => add_out_0_9_port, S(8) =>
                           add_out_0_8_port, S(7) => add_out_0_7_port, S(6) => 
                           add_out_0_6_port, S(5) => add_out_0_5_port, S(4) => 
                           add_out_0_4_port, S(3) => add_out_0_3_port, S(2) => 
                           add_out_0_2_port, S(1) => add_out_0_1_port, S(0) => 
                           add_out_0_0_port, Cout => n_1551);
   ADD_1i_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_5 port map( A(31) => 
                           add_out_0_31_port, A(30) => add_out_0_30_port, A(29)
                           => add_out_0_29_port, A(28) => add_out_0_28_port, 
                           A(27) => add_out_0_27_port, A(26) => 
                           add_out_0_26_port, A(25) => add_out_0_25_port, A(24)
                           => add_out_0_24_port, A(23) => add_out_0_23_port, 
                           A(22) => add_out_0_22_port, A(21) => 
                           add_out_0_21_port, A(20) => add_out_0_20_port, A(19)
                           => add_out_0_19_port, A(18) => add_out_0_18_port, 
                           A(17) => add_out_0_17_port, A(16) => 
                           add_out_0_16_port, A(15) => add_out_0_15_port, A(14)
                           => add_out_0_14_port, A(13) => add_out_0_13_port, 
                           A(12) => add_out_0_12_port, A(11) => 
                           add_out_0_11_port, A(10) => add_out_0_10_port, A(9) 
                           => add_out_0_9_port, A(8) => add_out_0_8_port, A(7) 
                           => add_out_0_7_port, A(6) => add_out_0_6_port, A(5) 
                           => add_out_0_5_port, A(4) => add_out_0_4_port, A(3) 
                           => add_out_0_3_port, A(2) => add_out_0_2_port, A(1) 
                           => add_out_0_1_port, A(0) => add_out_0_0_port, B(31)
                           => addends_3_31_port, B(30) => addends_3_30_port, 
                           B(29) => addends_3_29_port, B(28) => 
                           addends_3_28_port, B(27) => addends_3_27_port, B(26)
                           => addends_3_26_port, B(25) => addends_3_25_port, 
                           B(24) => addends_3_24_port, B(23) => 
                           addends_3_23_port, B(22) => addends_3_22_port, B(21)
                           => addends_3_21_port, B(20) => addends_3_20_port, 
                           B(19) => addends_3_19_port, B(18) => 
                           addends_3_18_port, B(17) => addends_3_17_port, B(16)
                           => addends_3_16_port, B(15) => addends_3_15_port, 
                           B(14) => addends_3_14_port, B(13) => 
                           addends_3_13_port, B(12) => addends_3_12_port, B(11)
                           => addends_3_11_port, B(10) => addends_3_10_port, 
                           B(9) => addends_3_9_port, B(8) => addends_3_8_port, 
                           B(7) => addends_3_7_port, B(6) => addends_3_6_port, 
                           B(5) => addends_3_5_port, B(4) => addends_3_4_port, 
                           B(3) => addends_3_3_port, B(2) => addends_3_2_port, 
                           B(1) => addends_3_1_port, B(0) => addends_3_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_1_31_port, S(30) => reg_in_1_30_port
                           , S(29) => reg_in_1_29_port, S(28) => 
                           reg_in_1_28_port, S(27) => reg_in_1_27_port, S(26) 
                           => reg_in_1_26_port, S(25) => reg_in_1_25_port, 
                           S(24) => reg_in_1_24_port, S(23) => reg_in_1_23_port
                           , S(22) => reg_in_1_22_port, S(21) => 
                           reg_in_1_21_port, S(20) => reg_in_1_20_port, S(19) 
                           => reg_in_1_19_port, S(18) => reg_in_1_18_port, 
                           S(17) => reg_in_1_17_port, S(16) => reg_in_1_16_port
                           , S(15) => reg_in_1_15_port, S(14) => 
                           reg_in_1_14_port, S(13) => reg_in_1_13_port, S(12) 
                           => reg_in_1_12_port, S(11) => reg_in_1_11_port, 
                           S(10) => reg_in_1_10_port, S(9) => reg_in_1_9_port, 
                           S(8) => reg_in_1_8_port, S(7) => reg_in_1_7_port, 
                           S(6) => reg_in_1_6_port, S(5) => reg_in_1_5_port, 
                           S(4) => reg_in_1_4_port, S(3) => reg_in_1_3_port, 
                           S(2) => reg_in_1_2_port, S(1) => reg_in_1_1_port, 
                           S(0) => reg_in_1_0_port, Cout => n_1552);
   REG_i_1 : REG_NBIT32_2 port map( clk => CLOCK, reset => X_Logic0_port, 
                           enable => X_Logic1_port, data_in(31) => 
                           reg_in_1_31_port, data_in(30) => reg_in_1_30_port, 
                           data_in(29) => reg_in_1_29_port, data_in(28) => 
                           reg_in_1_28_port, data_in(27) => reg_in_1_27_port, 
                           data_in(26) => reg_in_1_26_port, data_in(25) => 
                           reg_in_1_25_port, data_in(24) => reg_in_1_24_port, 
                           data_in(23) => reg_in_1_23_port, data_in(22) => 
                           reg_in_1_22_port, data_in(21) => reg_in_1_21_port, 
                           data_in(20) => reg_in_1_20_port, data_in(19) => 
                           reg_in_1_19_port, data_in(18) => reg_in_1_18_port, 
                           data_in(17) => reg_in_1_17_port, data_in(16) => 
                           reg_in_1_16_port, data_in(15) => reg_in_1_15_port, 
                           data_in(14) => reg_in_1_14_port, data_in(13) => 
                           reg_in_1_13_port, data_in(12) => reg_in_1_12_port, 
                           data_in(11) => reg_in_1_11_port, data_in(10) => 
                           reg_in_1_10_port, data_in(9) => reg_in_1_9_port, 
                           data_in(8) => reg_in_1_8_port, data_in(7) => 
                           reg_in_1_7_port, data_in(6) => reg_in_1_6_port, 
                           data_in(5) => reg_in_1_5_port, data_in(4) => 
                           reg_in_1_4_port, data_in(3) => reg_in_1_3_port, 
                           data_in(2) => reg_in_1_2_port, data_in(1) => 
                           reg_in_1_1_port, data_in(0) => reg_in_1_0_port, 
                           data_out(31) => reg_out_1_31_port, data_out(30) => 
                           reg_out_1_30_port, data_out(29) => reg_out_1_29_port
                           , data_out(28) => reg_out_1_28_port, data_out(27) =>
                           reg_out_1_27_port, data_out(26) => reg_out_1_26_port
                           , data_out(25) => reg_out_1_25_port, data_out(24) =>
                           reg_out_1_24_port, data_out(23) => reg_out_1_23_port
                           , data_out(22) => reg_out_1_22_port, data_out(21) =>
                           reg_out_1_21_port, data_out(20) => reg_out_1_20_port
                           , data_out(19) => reg_out_1_19_port, data_out(18) =>
                           reg_out_1_18_port, data_out(17) => reg_out_1_17_port
                           , data_out(16) => reg_out_1_16_port, data_out(15) =>
                           reg_out_1_15_port, data_out(14) => reg_out_1_14_port
                           , data_out(13) => reg_out_1_13_port, data_out(12) =>
                           reg_out_1_12_port, data_out(11) => reg_out_1_11_port
                           , data_out(10) => reg_out_1_10_port, data_out(9) => 
                           reg_out_1_9_port, data_out(8) => reg_out_1_8_port, 
                           data_out(7) => reg_out_1_7_port, data_out(6) => 
                           reg_out_1_6_port, data_out(5) => reg_out_1_5_port, 
                           data_out(4) => reg_out_1_4_port, data_out(3) => 
                           reg_out_1_3_port, data_out(2) => reg_out_1_2_port, 
                           data_out(1) => reg_out_1_1_port, data_out(0) => 
                           reg_out_1_0_port);
   ADD_0i_2 : ADDER_NBIT32_NBIT_PER_BLOCK4_4 port map( A(31) => 
                           reg_out_1_31_port, A(30) => reg_out_1_30_port, A(29)
                           => reg_out_1_29_port, A(28) => reg_out_1_28_port, 
                           A(27) => reg_out_1_27_port, A(26) => 
                           reg_out_1_26_port, A(25) => reg_out_1_25_port, A(24)
                           => reg_out_1_24_port, A(23) => reg_out_1_23_port, 
                           A(22) => reg_out_1_22_port, A(21) => 
                           reg_out_1_21_port, A(20) => reg_out_1_20_port, A(19)
                           => reg_out_1_19_port, A(18) => reg_out_1_18_port, 
                           A(17) => reg_out_1_17_port, A(16) => 
                           reg_out_1_16_port, A(15) => reg_out_1_15_port, A(14)
                           => reg_out_1_14_port, A(13) => reg_out_1_13_port, 
                           A(12) => reg_out_1_12_port, A(11) => 
                           reg_out_1_11_port, A(10) => reg_out_1_10_port, A(9) 
                           => reg_out_1_9_port, A(8) => reg_out_1_8_port, A(7) 
                           => reg_out_1_7_port, A(6) => reg_out_1_6_port, A(5) 
                           => reg_out_1_5_port, A(4) => reg_out_1_4_port, A(3) 
                           => reg_out_1_3_port, A(2) => reg_out_1_2_port, A(1) 
                           => reg_out_1_1_port, A(0) => reg_out_1_0_port, B(31)
                           => addends_4_31_port, B(30) => addends_4_30_port, 
                           B(29) => addends_4_29_port, B(28) => 
                           addends_4_28_port, B(27) => addends_4_27_port, B(26)
                           => addends_4_26_port, B(25) => addends_4_25_port, 
                           B(24) => addends_4_24_port, B(23) => 
                           addends_4_23_port, B(22) => addends_4_22_port, B(21)
                           => addends_4_21_port, B(20) => addends_4_20_port, 
                           B(19) => addends_4_19_port, B(18) => 
                           addends_4_18_port, B(17) => addends_4_17_port, B(16)
                           => addends_4_16_port, B(15) => addends_4_15_port, 
                           B(14) => addends_4_14_port, B(13) => 
                           addends_4_13_port, B(12) => addends_4_12_port, B(11)
                           => addends_4_11_port, B(10) => addends_4_10_port, 
                           B(9) => addends_4_9_port, B(8) => addends_4_8_port, 
                           B(7) => addends_4_7_port, B(6) => addends_4_6_port, 
                           B(5) => addends_4_5_port, B(4) => addends_4_4_port, 
                           B(3) => addends_4_3_port, B(2) => addends_4_2_port, 
                           B(1) => addends_4_1_port, B(0) => addends_4_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_1_31_port, S(30) => 
                           add_out_1_30_port, S(29) => add_out_1_29_port, S(28)
                           => add_out_1_28_port, S(27) => add_out_1_27_port, 
                           S(26) => add_out_1_26_port, S(25) => 
                           add_out_1_25_port, S(24) => add_out_1_24_port, S(23)
                           => add_out_1_23_port, S(22) => add_out_1_22_port, 
                           S(21) => add_out_1_21_port, S(20) => 
                           add_out_1_20_port, S(19) => add_out_1_19_port, S(18)
                           => add_out_1_18_port, S(17) => add_out_1_17_port, 
                           S(16) => add_out_1_16_port, S(15) => 
                           add_out_1_15_port, S(14) => add_out_1_14_port, S(13)
                           => add_out_1_13_port, S(12) => add_out_1_12_port, 
                           S(11) => add_out_1_11_port, S(10) => 
                           add_out_1_10_port, S(9) => add_out_1_9_port, S(8) =>
                           add_out_1_8_port, S(7) => add_out_1_7_port, S(6) => 
                           add_out_1_6_port, S(5) => add_out_1_5_port, S(4) => 
                           add_out_1_4_port, S(3) => add_out_1_3_port, S(2) => 
                           add_out_1_2_port, S(1) => add_out_1_1_port, S(0) => 
                           add_out_1_0_port, Cout => n_1553);
   ADD_1i_2 : ADDER_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => 
                           add_out_1_31_port, A(30) => add_out_1_30_port, A(29)
                           => add_out_1_29_port, A(28) => add_out_1_28_port, 
                           A(27) => add_out_1_27_port, A(26) => 
                           add_out_1_26_port, A(25) => add_out_1_25_port, A(24)
                           => add_out_1_24_port, A(23) => add_out_1_23_port, 
                           A(22) => add_out_1_22_port, A(21) => 
                           add_out_1_21_port, A(20) => add_out_1_20_port, A(19)
                           => add_out_1_19_port, A(18) => add_out_1_18_port, 
                           A(17) => add_out_1_17_port, A(16) => 
                           add_out_1_16_port, A(15) => add_out_1_15_port, A(14)
                           => add_out_1_14_port, A(13) => add_out_1_13_port, 
                           A(12) => add_out_1_12_port, A(11) => 
                           add_out_1_11_port, A(10) => add_out_1_10_port, A(9) 
                           => add_out_1_9_port, A(8) => add_out_1_8_port, A(7) 
                           => add_out_1_7_port, A(6) => add_out_1_6_port, A(5) 
                           => add_out_1_5_port, A(4) => add_out_1_4_port, A(3) 
                           => add_out_1_3_port, A(2) => add_out_1_2_port, A(1) 
                           => add_out_1_1_port, A(0) => add_out_1_0_port, B(31)
                           => addends_5_31_port, B(30) => addends_5_30_port, 
                           B(29) => addends_5_29_port, B(28) => 
                           addends_5_28_port, B(27) => addends_5_27_port, B(26)
                           => addends_5_26_port, B(25) => addends_5_25_port, 
                           B(24) => addends_5_24_port, B(23) => 
                           addends_5_23_port, B(22) => addends_5_22_port, B(21)
                           => addends_5_21_port, B(20) => addends_5_20_port, 
                           B(19) => addends_5_19_port, B(18) => 
                           addends_5_18_port, B(17) => addends_5_17_port, B(16)
                           => addends_5_16_port, B(15) => addends_5_15_port, 
                           B(14) => addends_5_14_port, B(13) => 
                           addends_5_13_port, B(12) => addends_5_12_port, B(11)
                           => addends_5_11_port, B(10) => addends_5_10_port, 
                           B(9) => addends_5_9_port, B(8) => addends_5_8_port, 
                           B(7) => addends_5_7_port, B(6) => addends_5_6_port, 
                           B(5) => addends_5_5_port, B(4) => addends_5_4_port, 
                           B(3) => addends_5_3_port, B(2) => addends_5_2_port, 
                           B(1) => addends_5_1_port, B(0) => addends_5_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => reg_in_2_31_port, S(30) => reg_in_2_30_port
                           , S(29) => reg_in_2_29_port, S(28) => 
                           reg_in_2_28_port, S(27) => reg_in_2_27_port, S(26) 
                           => reg_in_2_26_port, S(25) => reg_in_2_25_port, 
                           S(24) => reg_in_2_24_port, S(23) => reg_in_2_23_port
                           , S(22) => reg_in_2_22_port, S(21) => 
                           reg_in_2_21_port, S(20) => reg_in_2_20_port, S(19) 
                           => reg_in_2_19_port, S(18) => reg_in_2_18_port, 
                           S(17) => reg_in_2_17_port, S(16) => reg_in_2_16_port
                           , S(15) => reg_in_2_15_port, S(14) => 
                           reg_in_2_14_port, S(13) => reg_in_2_13_port, S(12) 
                           => reg_in_2_12_port, S(11) => reg_in_2_11_port, 
                           S(10) => reg_in_2_10_port, S(9) => reg_in_2_9_port, 
                           S(8) => reg_in_2_8_port, S(7) => reg_in_2_7_port, 
                           S(6) => reg_in_2_6_port, S(5) => reg_in_2_5_port, 
                           S(4) => reg_in_2_4_port, S(3) => reg_in_2_3_port, 
                           S(2) => reg_in_2_2_port, S(1) => reg_in_2_1_port, 
                           S(0) => reg_in_2_0_port, Cout => n_1554);
   REG_i_2 : REG_NBIT32_1 port map( clk => CLOCK, reset => X_Logic0_port, 
                           enable => X_Logic1_port, data_in(31) => 
                           reg_in_2_31_port, data_in(30) => reg_in_2_30_port, 
                           data_in(29) => reg_in_2_29_port, data_in(28) => 
                           reg_in_2_28_port, data_in(27) => reg_in_2_27_port, 
                           data_in(26) => reg_in_2_26_port, data_in(25) => 
                           reg_in_2_25_port, data_in(24) => reg_in_2_24_port, 
                           data_in(23) => reg_in_2_23_port, data_in(22) => 
                           reg_in_2_22_port, data_in(21) => reg_in_2_21_port, 
                           data_in(20) => reg_in_2_20_port, data_in(19) => 
                           reg_in_2_19_port, data_in(18) => reg_in_2_18_port, 
                           data_in(17) => reg_in_2_17_port, data_in(16) => 
                           reg_in_2_16_port, data_in(15) => reg_in_2_15_port, 
                           data_in(14) => reg_in_2_14_port, data_in(13) => 
                           reg_in_2_13_port, data_in(12) => reg_in_2_12_port, 
                           data_in(11) => reg_in_2_11_port, data_in(10) => 
                           reg_in_2_10_port, data_in(9) => reg_in_2_9_port, 
                           data_in(8) => reg_in_2_8_port, data_in(7) => 
                           reg_in_2_7_port, data_in(6) => reg_in_2_6_port, 
                           data_in(5) => reg_in_2_5_port, data_in(4) => 
                           reg_in_2_4_port, data_in(3) => reg_in_2_3_port, 
                           data_in(2) => reg_in_2_2_port, data_in(1) => 
                           reg_in_2_1_port, data_in(0) => reg_in_2_0_port, 
                           data_out(31) => reg_out_2_31_port, data_out(30) => 
                           reg_out_2_30_port, data_out(29) => reg_out_2_29_port
                           , data_out(28) => reg_out_2_28_port, data_out(27) =>
                           reg_out_2_27_port, data_out(26) => reg_out_2_26_port
                           , data_out(25) => reg_out_2_25_port, data_out(24) =>
                           reg_out_2_24_port, data_out(23) => reg_out_2_23_port
                           , data_out(22) => reg_out_2_22_port, data_out(21) =>
                           reg_out_2_21_port, data_out(20) => reg_out_2_20_port
                           , data_out(19) => reg_out_2_19_port, data_out(18) =>
                           reg_out_2_18_port, data_out(17) => reg_out_2_17_port
                           , data_out(16) => reg_out_2_16_port, data_out(15) =>
                           reg_out_2_15_port, data_out(14) => reg_out_2_14_port
                           , data_out(13) => reg_out_2_13_port, data_out(12) =>
                           reg_out_2_12_port, data_out(11) => reg_out_2_11_port
                           , data_out(10) => reg_out_2_10_port, data_out(9) => 
                           reg_out_2_9_port, data_out(8) => reg_out_2_8_port, 
                           data_out(7) => reg_out_2_7_port, data_out(6) => 
                           reg_out_2_6_port, data_out(5) => reg_out_2_5_port, 
                           data_out(4) => reg_out_2_4_port, data_out(3) => 
                           reg_out_2_3_port, data_out(2) => reg_out_2_2_port, 
                           data_out(1) => reg_out_2_1_port, data_out(0) => 
                           reg_out_2_0_port);
   ADD_N_1 : ADDER_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => 
                           reg_out_2_31_port, A(30) => reg_out_2_30_port, A(29)
                           => reg_out_2_29_port, A(28) => reg_out_2_28_port, 
                           A(27) => reg_out_2_27_port, A(26) => 
                           reg_out_2_26_port, A(25) => reg_out_2_25_port, A(24)
                           => reg_out_2_24_port, A(23) => reg_out_2_23_port, 
                           A(22) => reg_out_2_22_port, A(21) => 
                           reg_out_2_21_port, A(20) => reg_out_2_20_port, A(19)
                           => reg_out_2_19_port, A(18) => reg_out_2_18_port, 
                           A(17) => reg_out_2_17_port, A(16) => 
                           reg_out_2_16_port, A(15) => reg_out_2_15_port, A(14)
                           => reg_out_2_14_port, A(13) => reg_out_2_13_port, 
                           A(12) => reg_out_2_12_port, A(11) => 
                           reg_out_2_11_port, A(10) => reg_out_2_10_port, A(9) 
                           => reg_out_2_9_port, A(8) => reg_out_2_8_port, A(7) 
                           => reg_out_2_7_port, A(6) => reg_out_2_6_port, A(5) 
                           => reg_out_2_5_port, A(4) => reg_out_2_4_port, A(3) 
                           => reg_out_2_3_port, A(2) => reg_out_2_2_port, A(1) 
                           => reg_out_2_1_port, A(0) => reg_out_2_0_port, B(31)
                           => addends_6_31_port, B(30) => addends_6_30_port, 
                           B(29) => addends_6_29_port, B(28) => 
                           addends_6_28_port, B(27) => addends_6_27_port, B(26)
                           => addends_6_26_port, B(25) => addends_6_25_port, 
                           B(24) => addends_6_24_port, B(23) => 
                           addends_6_23_port, B(22) => addends_6_22_port, B(21)
                           => addends_6_21_port, B(20) => addends_6_20_port, 
                           B(19) => addends_6_19_port, B(18) => 
                           addends_6_18_port, B(17) => addends_6_17_port, B(16)
                           => addends_6_16_port, B(15) => addends_6_15_port, 
                           B(14) => addends_6_14_port, B(13) => 
                           addends_6_13_port, B(12) => addends_6_12_port, B(11)
                           => addends_6_11_port, B(10) => addends_6_10_port, 
                           B(9) => addends_6_9_port, B(8) => addends_6_8_port, 
                           B(7) => addends_6_7_port, B(6) => addends_6_6_port, 
                           B(5) => addends_6_5_port, B(4) => addends_6_4_port, 
                           B(3) => addends_6_3_port, B(2) => addends_6_2_port, 
                           B(1) => addends_6_1_port, B(0) => addends_6_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => add_out_2_31_port, S(30) => 
                           add_out_2_30_port, S(29) => add_out_2_29_port, S(28)
                           => add_out_2_28_port, S(27) => add_out_2_27_port, 
                           S(26) => add_out_2_26_port, S(25) => 
                           add_out_2_25_port, S(24) => add_out_2_24_port, S(23)
                           => add_out_2_23_port, S(22) => add_out_2_22_port, 
                           S(21) => add_out_2_21_port, S(20) => 
                           add_out_2_20_port, S(19) => add_out_2_19_port, S(18)
                           => add_out_2_18_port, S(17) => add_out_2_17_port, 
                           S(16) => add_out_2_16_port, S(15) => 
                           add_out_2_15_port, S(14) => add_out_2_14_port, S(13)
                           => add_out_2_13_port, S(12) => add_out_2_12_port, 
                           S(11) => add_out_2_11_port, S(10) => 
                           add_out_2_10_port, S(9) => add_out_2_9_port, S(8) =>
                           add_out_2_8_port, S(7) => add_out_2_7_port, S(6) => 
                           add_out_2_6_port, S(5) => add_out_2_5_port, S(4) => 
                           add_out_2_4_port, S(3) => add_out_2_3_port, S(2) => 
                           add_out_2_2_port, S(1) => add_out_2_1_port, S(0) => 
                           add_out_2_0_port, Cout => n_1555);
   ADD_N : ADDER_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => add_out_2_31_port,
                           A(30) => add_out_2_30_port, A(29) => 
                           add_out_2_29_port, A(28) => add_out_2_28_port, A(27)
                           => add_out_2_27_port, A(26) => add_out_2_26_port, 
                           A(25) => add_out_2_25_port, A(24) => 
                           add_out_2_24_port, A(23) => add_out_2_23_port, A(22)
                           => add_out_2_22_port, A(21) => add_out_2_21_port, 
                           A(20) => add_out_2_20_port, A(19) => 
                           add_out_2_19_port, A(18) => add_out_2_18_port, A(17)
                           => add_out_2_17_port, A(16) => add_out_2_16_port, 
                           A(15) => add_out_2_15_port, A(14) => 
                           add_out_2_14_port, A(13) => add_out_2_13_port, A(12)
                           => add_out_2_12_port, A(11) => add_out_2_11_port, 
                           A(10) => add_out_2_10_port, A(9) => add_out_2_9_port
                           , A(8) => add_out_2_8_port, A(7) => add_out_2_7_port
                           , A(6) => add_out_2_6_port, A(5) => add_out_2_5_port
                           , A(4) => add_out_2_4_port, A(3) => add_out_2_3_port
                           , A(2) => add_out_2_2_port, A(1) => add_out_2_1_port
                           , A(0) => add_out_2_0_port, B(31) => 
                           addends_7_31_port, B(30) => addends_7_30_port, B(29)
                           => addends_7_29_port, B(28) => addends_7_28_port, 
                           B(27) => addends_7_27_port, B(26) => 
                           addends_7_26_port, B(25) => addends_7_25_port, B(24)
                           => addends_7_24_port, B(23) => addends_7_23_port, 
                           B(22) => addends_7_22_port, B(21) => 
                           addends_7_21_port, B(20) => addends_7_20_port, B(19)
                           => addends_7_19_port, B(18) => addends_7_18_port, 
                           B(17) => addends_7_17_port, B(16) => 
                           addends_7_16_port, B(15) => addends_7_15_port, B(14)
                           => addends_7_14_port, B(13) => addends_7_13_port, 
                           B(12) => addends_7_12_port, B(11) => 
                           addends_7_11_port, B(10) => addends_7_10_port, B(9) 
                           => addends_7_9_port, B(8) => addends_7_8_port, B(7) 
                           => addends_7_7_port, B(6) => addends_7_6_port, B(5) 
                           => addends_7_5_port, B(4) => addends_7_4_port, B(3) 
                           => addends_7_3_port, B(2) => addends_7_2_port, B(1) 
                           => addends_7_1_port, B(0) => addends_7_0_port, 
                           ADD_SUB => X_Logic0_port, Cin => X_Logic0_port, 
                           S(31) => Y(31), S(30) => Y(30), S(29) => Y(29), 
                           S(28) => Y(28), S(27) => Y(27), S(26) => Y(26), 
                           S(25) => Y(25), S(24) => Y(24), S(23) => Y(23), 
                           S(22) => Y(22), S(21) => Y(21), S(20) => Y(20), 
                           S(19) => Y(19), S(18) => Y(18), S(17) => Y(17), 
                           S(16) => Y(16), S(15) => Y(15), S(14) => Y(14), 
                           S(13) => Y(13), S(12) => Y(12), S(11) => Y(11), 
                           S(10) => Y(10), S(9) => Y(9), S(8) => Y(8), S(7) => 
                           Y(7), S(6) => Y(6), S(5) => Y(5), S(4) => Y(4), S(3)
                           => Y(3), S(2) => Y(2), S(1) => Y(1), S(0) => Y(0), 
                           Cout => n_1556);
   addends_reg_6_2_inst : DFF_X1 port map( D => pipe2_0_2_port, CK => CLOCK, Q 
                           => addends_6_2_port, QN => n_1557);
   addends_reg_6_1_inst : DFF_X1 port map( D => pipe2_0_1_port, CK => CLOCK, Q 
                           => addends_6_1_port, QN => n_1558);
   addends_reg_4_0_inst : DFF_X1 port map( D => pipe1_0_0_port, CK => CLOCK, Q 
                           => addends_4_0_port, QN => n_1559);
   addends_reg_6_0_inst : DFF_X1 port map( D => pipe2_0_0_port, CK => CLOCK, Q 
                           => addends_6_0_port, QN => n_1560);
   addends_reg_6_3_inst : DFF_X1 port map( D => pipe2_0_3_port, CK => CLOCK, Q 
                           => addends_6_3_port, QN => n_1561);
   U3 : NAND2_X1 port map( A1 => sub_126_G16_carry_30_port, A2 => n67, ZN => n1
                           );
   U4 : BUF_X1 port map( A => n68, Z => n66);
   U5 : BUF_X1 port map( A => n26, Z => n24);
   U6 : BUF_X1 port map( A => n29, Z => n27);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n35, Z => n33);
   U9 : BUF_X1 port map( A => n38, Z => n36);
   U10 : BUF_X1 port map( A => n41, Z => n39);
   U11 : BUF_X1 port map( A => n44, Z => n42);
   U12 : BUF_X1 port map( A => n47, Z => n45);
   U13 : BUF_X1 port map( A => n50, Z => n48);
   U14 : BUF_X1 port map( A => n53, Z => n51);
   U15 : BUF_X1 port map( A => n56, Z => n54);
   U16 : BUF_X1 port map( A => n59, Z => n57);
   U17 : BUF_X1 port map( A => n62, Z => n60);
   U18 : BUF_X1 port map( A => n65, Z => n63);
   U19 : BUF_X1 port map( A => n23, Z => n21);
   U20 : BUF_X1 port map( A => n23, Z => n22);
   U21 : NAND2_X1 port map( A1 => sub_126_G5_carry_19_port, A2 => n67, ZN => n2
                           );
   U22 : NAND2_X1 port map( A1 => sub_126_G6_carry_20_port, A2 => n67, ZN => n3
                           );
   U23 : NAND2_X1 port map( A1 => sub_126_G7_carry_21_port, A2 => n67, ZN => n4
                           );
   U24 : NAND2_X1 port map( A1 => sub_126_G8_carry_22_port, A2 => n67, ZN => n5
                           );
   U25 : NAND2_X1 port map( A1 => sub_126_carry_15_port, A2 => n66, ZN => n6);
   U26 : NAND2_X1 port map( A1 => sub_126_G9_carry_23_port, A2 => n67, ZN => n7
                           );
   U27 : NAND2_X1 port map( A1 => sub_126_G2_carry_16_port, A2 => n67, ZN => n8
                           );
   U28 : NAND2_X1 port map( A1 => sub_126_G3_carry_17_port, A2 => n67, ZN => n9
                           );
   U29 : NAND2_X1 port map( A1 => sub_126_G10_carry_24_port, A2 => n67, ZN => 
                           n10);
   U30 : NAND2_X1 port map( A1 => sub_126_G4_carry_18_port, A2 => n67, ZN => 
                           n11);
   U31 : NAND2_X1 port map( A1 => sub_126_G11_carry_25_port, A2 => n67, ZN => 
                           n12);
   U32 : NAND2_X1 port map( A1 => sub_126_G12_carry_26_port, A2 => n67, ZN => 
                           n13);
   U33 : NAND2_X1 port map( A1 => sub_126_G13_carry_27_port, A2 => n67, ZN => 
                           n14);
   U34 : NAND2_X1 port map( A1 => sub_126_G14_carry_28_port, A2 => n67, ZN => 
                           n15);
   U35 : NAND2_X1 port map( A1 => sub_126_G15_carry_29_port, A2 => n67, ZN => 
                           n16);
   U36 : INV_X1 port map( A => n21, ZN => n20);
   U37 : BUF_X1 port map( A => n22, Z => n18);
   U38 : BUF_X1 port map( A => n22, Z => n17);
   U39 : BUF_X1 port map( A => n22, Z => n19);
   U40 : BUF_X1 port map( A => n26, Z => n25);
   U41 : BUF_X1 port map( A => n29, Z => n28);
   U42 : BUF_X1 port map( A => n32, Z => n31);
   U43 : BUF_X1 port map( A => n35, Z => n34);
   U44 : BUF_X1 port map( A => n38, Z => n37);
   U45 : BUF_X1 port map( A => n41, Z => n40);
   U46 : BUF_X1 port map( A => n44, Z => n43);
   U47 : BUF_X1 port map( A => n47, Z => n46);
   U48 : BUF_X1 port map( A => n50, Z => n49);
   U49 : BUF_X1 port map( A => n53, Z => n52);
   U50 : BUF_X1 port map( A => n56, Z => n55);
   U51 : BUF_X1 port map( A => n59, Z => n58);
   U52 : BUF_X1 port map( A => n62, Z => n61);
   U53 : BUF_X1 port map( A => n65, Z => n64);
   U54 : BUF_X1 port map( A => n68, Z => n67);
   U55 : INV_X1 port map( A => A(0), ZN => n23);
   U56 : INV_X1 port map( A => A(1), ZN => n26);
   U57 : INV_X1 port map( A => A(2), ZN => n29);
   U58 : INV_X1 port map( A => A(3), ZN => n32);
   U59 : INV_X1 port map( A => A(4), ZN => n35);
   U60 : INV_X1 port map( A => A(5), ZN => n38);
   U61 : INV_X1 port map( A => A(6), ZN => n41);
   U62 : INV_X1 port map( A => A(7), ZN => n44);
   U63 : INV_X1 port map( A => A(8), ZN => n47);
   U64 : INV_X1 port map( A => A(9), ZN => n50);
   U65 : INV_X1 port map( A => A(10), ZN => n53);
   U66 : INV_X1 port map( A => A(11), ZN => n56);
   U67 : INV_X1 port map( A => A(12), ZN => n59);
   U68 : INV_X1 port map( A => A(13), ZN => n62);
   U69 : INV_X1 port map( A => A(14), ZN => n65);
   U70 : INV_X1 port map( A => A(15), ZN => n68);
   U71 : XOR2_X1 port map( A => n66, B => sub_126_G2_carry_16_port, Z => 
                           A_neg_1_16_port);
   U72 : AND2_X1 port map( A1 => sub_126_G2_carry_15_port, A2 => n64, ZN => 
                           sub_126_G2_carry_16_port);
   U73 : XOR2_X1 port map( A => n63, B => sub_126_G2_carry_15_port, Z => 
                           A_neg_1_15_port);
   U74 : AND2_X1 port map( A1 => sub_126_G2_carry_14_port, A2 => n61, ZN => 
                           sub_126_G2_carry_15_port);
   U75 : XOR2_X1 port map( A => n60, B => sub_126_G2_carry_14_port, Z => 
                           A_neg_1_14_port);
   U76 : AND2_X1 port map( A1 => sub_126_G2_carry_13_port, A2 => n58, ZN => 
                           sub_126_G2_carry_14_port);
   U77 : XOR2_X1 port map( A => n57, B => sub_126_G2_carry_13_port, Z => 
                           A_neg_1_13_port);
   U78 : AND2_X1 port map( A1 => sub_126_G2_carry_12_port, A2 => n55, ZN => 
                           sub_126_G2_carry_13_port);
   U79 : XOR2_X1 port map( A => n54, B => sub_126_G2_carry_12_port, Z => 
                           A_neg_1_12_port);
   U80 : AND2_X1 port map( A1 => sub_126_G2_carry_11_port, A2 => n52, ZN => 
                           sub_126_G2_carry_12_port);
   U81 : XOR2_X1 port map( A => n51, B => sub_126_G2_carry_11_port, Z => 
                           A_neg_1_11_port);
   U82 : AND2_X1 port map( A1 => sub_126_G2_carry_10_port, A2 => n49, ZN => 
                           sub_126_G2_carry_11_port);
   U83 : XOR2_X1 port map( A => n48, B => sub_126_G2_carry_10_port, Z => 
                           A_neg_1_10_port);
   U84 : AND2_X1 port map( A1 => sub_126_G2_carry_9_port, A2 => n46, ZN => 
                           sub_126_G2_carry_10_port);
   U85 : XOR2_X1 port map( A => n45, B => sub_126_G2_carry_9_port, Z => 
                           A_neg_1_9_port);
   U86 : AND2_X1 port map( A1 => sub_126_G2_carry_8_port, A2 => n43, ZN => 
                           sub_126_G2_carry_9_port);
   U87 : XOR2_X1 port map( A => n42, B => sub_126_G2_carry_8_port, Z => 
                           A_neg_1_8_port);
   U88 : AND2_X1 port map( A1 => sub_126_G2_carry_7_port, A2 => n40, ZN => 
                           sub_126_G2_carry_8_port);
   U89 : XOR2_X1 port map( A => n39, B => sub_126_G2_carry_7_port, Z => 
                           A_neg_1_7_port);
   U90 : AND2_X1 port map( A1 => sub_126_G2_carry_6_port, A2 => n37, ZN => 
                           sub_126_G2_carry_7_port);
   U91 : XOR2_X1 port map( A => n36, B => sub_126_G2_carry_6_port, Z => 
                           A_neg_1_6_port);
   U92 : AND2_X1 port map( A1 => sub_126_G2_carry_5_port, A2 => n34, ZN => 
                           sub_126_G2_carry_6_port);
   U93 : XOR2_X1 port map( A => n33, B => sub_126_G2_carry_5_port, Z => 
                           A_neg_1_5_port);
   U94 : AND2_X1 port map( A1 => sub_126_G2_carry_4_port, A2 => n31, ZN => 
                           sub_126_G2_carry_5_port);
   U95 : XOR2_X1 port map( A => n30, B => sub_126_G2_carry_4_port, Z => 
                           A_neg_1_4_port);
   U96 : AND2_X1 port map( A1 => sub_126_G2_carry_3_port, A2 => n28, ZN => 
                           sub_126_G2_carry_4_port);
   U97 : XOR2_X1 port map( A => n27, B => sub_126_G2_carry_3_port, Z => 
                           A_neg_1_3_port);
   U98 : AND2_X1 port map( A1 => n19, A2 => n25, ZN => sub_126_G2_carry_3_port)
                           ;
   U99 : XOR2_X1 port map( A => n24, B => n18, Z => A_neg_1_2_port);
   U100 : XOR2_X1 port map( A => n66, B => sub_126_carry_15_port, Z => 
                           A_neg_0_15_port);
   U101 : AND2_X1 port map( A1 => sub_126_carry_14_port, A2 => n63, ZN => 
                           sub_126_carry_15_port);
   U102 : XOR2_X1 port map( A => n63, B => sub_126_carry_14_port, Z => 
                           A_neg_0_14_port);
   U103 : AND2_X1 port map( A1 => sub_126_carry_13_port, A2 => n60, ZN => 
                           sub_126_carry_14_port);
   U104 : XOR2_X1 port map( A => n60, B => sub_126_carry_13_port, Z => 
                           A_neg_0_13_port);
   U105 : AND2_X1 port map( A1 => sub_126_carry_12_port, A2 => n57, ZN => 
                           sub_126_carry_13_port);
   U106 : XOR2_X1 port map( A => n57, B => sub_126_carry_12_port, Z => 
                           A_neg_0_12_port);
   U107 : AND2_X1 port map( A1 => sub_126_carry_11_port, A2 => n54, ZN => 
                           sub_126_carry_12_port);
   U108 : XOR2_X1 port map( A => n54, B => sub_126_carry_11_port, Z => 
                           A_neg_0_11_port);
   U109 : AND2_X1 port map( A1 => sub_126_carry_10_port, A2 => n51, ZN => 
                           sub_126_carry_11_port);
   U110 : XOR2_X1 port map( A => n51, B => sub_126_carry_10_port, Z => 
                           A_neg_0_10_port);
   U111 : AND2_X1 port map( A1 => sub_126_carry_9_port, A2 => n48, ZN => 
                           sub_126_carry_10_port);
   U112 : XOR2_X1 port map( A => n48, B => sub_126_carry_9_port, Z => 
                           A_neg_0_9_port);
   U113 : AND2_X1 port map( A1 => sub_126_carry_8_port, A2 => n45, ZN => 
                           sub_126_carry_9_port);
   U114 : XOR2_X1 port map( A => n45, B => sub_126_carry_8_port, Z => 
                           A_neg_0_8_port);
   U115 : AND2_X1 port map( A1 => sub_126_carry_7_port, A2 => n42, ZN => 
                           sub_126_carry_8_port);
   U116 : XOR2_X1 port map( A => n42, B => sub_126_carry_7_port, Z => 
                           A_neg_0_7_port);
   U117 : AND2_X1 port map( A1 => sub_126_carry_6_port, A2 => n39, ZN => 
                           sub_126_carry_7_port);
   U118 : XOR2_X1 port map( A => n39, B => sub_126_carry_6_port, Z => 
                           A_neg_0_6_port);
   U119 : AND2_X1 port map( A1 => sub_126_carry_5_port, A2 => n36, ZN => 
                           sub_126_carry_6_port);
   U120 : XOR2_X1 port map( A => n36, B => sub_126_carry_5_port, Z => 
                           A_neg_0_5_port);
   U121 : AND2_X1 port map( A1 => sub_126_carry_4_port, A2 => n33, ZN => 
                           sub_126_carry_5_port);
   U122 : XOR2_X1 port map( A => n33, B => sub_126_carry_4_port, Z => 
                           A_neg_0_4_port);
   U123 : AND2_X1 port map( A1 => sub_126_carry_3_port, A2 => n30, ZN => 
                           sub_126_carry_4_port);
   U124 : XOR2_X1 port map( A => n30, B => sub_126_carry_3_port, Z => 
                           A_neg_0_3_port);
   U125 : AND2_X1 port map( A1 => sub_126_carry_2_port, A2 => n27, ZN => 
                           sub_126_carry_3_port);
   U126 : XOR2_X1 port map( A => n27, B => sub_126_carry_2_port, Z => 
                           A_neg_0_2_port);
   U127 : AND2_X1 port map( A1 => n19, A2 => n24, ZN => sub_126_carry_2_port);
   U128 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_0_1_port);
   U129 : XOR2_X1 port map( A => n66, B => sub_126_G4_carry_18_port, Z => 
                           A_neg_3_18_port);
   U130 : AND2_X1 port map( A1 => sub_126_G4_carry_17_port, A2 => n64, ZN => 
                           sub_126_G4_carry_18_port);
   U131 : XOR2_X1 port map( A => n63, B => sub_126_G4_carry_17_port, Z => 
                           A_neg_3_17_port);
   U132 : AND2_X1 port map( A1 => sub_126_G4_carry_16_port, A2 => n61, ZN => 
                           sub_126_G4_carry_17_port);
   U133 : XOR2_X1 port map( A => n60, B => sub_126_G4_carry_16_port, Z => 
                           A_neg_3_16_port);
   U134 : AND2_X1 port map( A1 => sub_126_G4_carry_15_port, A2 => n58, ZN => 
                           sub_126_G4_carry_16_port);
   U135 : XOR2_X1 port map( A => n57, B => sub_126_G4_carry_15_port, Z => 
                           A_neg_3_15_port);
   U136 : AND2_X1 port map( A1 => sub_126_G4_carry_14_port, A2 => n55, ZN => 
                           sub_126_G4_carry_15_port);
   U137 : XOR2_X1 port map( A => n54, B => sub_126_G4_carry_14_port, Z => 
                           A_neg_3_14_port);
   U138 : AND2_X1 port map( A1 => sub_126_G4_carry_13_port, A2 => n52, ZN => 
                           sub_126_G4_carry_14_port);
   U139 : XOR2_X1 port map( A => n51, B => sub_126_G4_carry_13_port, Z => 
                           A_neg_3_13_port);
   U140 : AND2_X1 port map( A1 => sub_126_G4_carry_12_port, A2 => n49, ZN => 
                           sub_126_G4_carry_13_port);
   U141 : XOR2_X1 port map( A => n48, B => sub_126_G4_carry_12_port, Z => 
                           A_neg_3_12_port);
   U142 : AND2_X1 port map( A1 => sub_126_G4_carry_11_port, A2 => n46, ZN => 
                           sub_126_G4_carry_12_port);
   U143 : XOR2_X1 port map( A => n45, B => sub_126_G4_carry_11_port, Z => 
                           A_neg_3_11_port);
   U144 : AND2_X1 port map( A1 => sub_126_G4_carry_10_port, A2 => n43, ZN => 
                           sub_126_G4_carry_11_port);
   U145 : XOR2_X1 port map( A => n42, B => sub_126_G4_carry_10_port, Z => 
                           A_neg_3_10_port);
   U146 : AND2_X1 port map( A1 => sub_126_G4_carry_9_port, A2 => n40, ZN => 
                           sub_126_G4_carry_10_port);
   U147 : XOR2_X1 port map( A => n39, B => sub_126_G4_carry_9_port, Z => 
                           A_neg_3_9_port);
   U148 : AND2_X1 port map( A1 => sub_126_G4_carry_8_port, A2 => n37, ZN => 
                           sub_126_G4_carry_9_port);
   U149 : XOR2_X1 port map( A => n36, B => sub_126_G4_carry_8_port, Z => 
                           A_neg_3_8_port);
   U150 : AND2_X1 port map( A1 => sub_126_G4_carry_7_port, A2 => n34, ZN => 
                           sub_126_G4_carry_8_port);
   U151 : XOR2_X1 port map( A => n33, B => sub_126_G4_carry_7_port, Z => 
                           A_neg_3_7_port);
   U152 : AND2_X1 port map( A1 => sub_126_G4_carry_6_port, A2 => n31, ZN => 
                           sub_126_G4_carry_7_port);
   U153 : XOR2_X1 port map( A => n30, B => sub_126_G4_carry_6_port, Z => 
                           A_neg_3_6_port);
   U154 : AND2_X1 port map( A1 => sub_126_G4_carry_5_port, A2 => n28, ZN => 
                           sub_126_G4_carry_6_port);
   U155 : XOR2_X1 port map( A => n27, B => sub_126_G4_carry_5_port, Z => 
                           A_neg_3_5_port);
   U156 : AND2_X1 port map( A1 => n19, A2 => n25, ZN => sub_126_G4_carry_5_port
                           );
   U157 : XOR2_X1 port map( A => n24, B => n18, Z => A_neg_3_4_port);
   U158 : XOR2_X1 port map( A => n66, B => sub_126_G3_carry_17_port, Z => 
                           A_neg_2_17_port);
   U159 : AND2_X1 port map( A1 => sub_126_G3_carry_16_port, A2 => n64, ZN => 
                           sub_126_G3_carry_17_port);
   U160 : XOR2_X1 port map( A => n63, B => sub_126_G3_carry_16_port, Z => 
                           A_neg_2_16_port);
   U161 : AND2_X1 port map( A1 => sub_126_G3_carry_15_port, A2 => n61, ZN => 
                           sub_126_G3_carry_16_port);
   U162 : XOR2_X1 port map( A => n60, B => sub_126_G3_carry_15_port, Z => 
                           A_neg_2_15_port);
   U163 : AND2_X1 port map( A1 => sub_126_G3_carry_14_port, A2 => n58, ZN => 
                           sub_126_G3_carry_15_port);
   U164 : XOR2_X1 port map( A => n57, B => sub_126_G3_carry_14_port, Z => 
                           A_neg_2_14_port);
   U165 : AND2_X1 port map( A1 => sub_126_G3_carry_13_port, A2 => n55, ZN => 
                           sub_126_G3_carry_14_port);
   U166 : XOR2_X1 port map( A => n54, B => sub_126_G3_carry_13_port, Z => 
                           A_neg_2_13_port);
   U167 : AND2_X1 port map( A1 => sub_126_G3_carry_12_port, A2 => n52, ZN => 
                           sub_126_G3_carry_13_port);
   U168 : XOR2_X1 port map( A => n51, B => sub_126_G3_carry_12_port, Z => 
                           A_neg_2_12_port);
   U169 : AND2_X1 port map( A1 => sub_126_G3_carry_11_port, A2 => n49, ZN => 
                           sub_126_G3_carry_12_port);
   U170 : XOR2_X1 port map( A => n48, B => sub_126_G3_carry_11_port, Z => 
                           A_neg_2_11_port);
   U171 : AND2_X1 port map( A1 => sub_126_G3_carry_10_port, A2 => n46, ZN => 
                           sub_126_G3_carry_11_port);
   U172 : XOR2_X1 port map( A => n45, B => sub_126_G3_carry_10_port, Z => 
                           A_neg_2_10_port);
   U173 : AND2_X1 port map( A1 => sub_126_G3_carry_9_port, A2 => n43, ZN => 
                           sub_126_G3_carry_10_port);
   U174 : XOR2_X1 port map( A => n42, B => sub_126_G3_carry_9_port, Z => 
                           A_neg_2_9_port);
   U175 : AND2_X1 port map( A1 => sub_126_G3_carry_8_port, A2 => n40, ZN => 
                           sub_126_G3_carry_9_port);
   U176 : XOR2_X1 port map( A => n39, B => sub_126_G3_carry_8_port, Z => 
                           A_neg_2_8_port);
   U177 : AND2_X1 port map( A1 => sub_126_G3_carry_7_port, A2 => n37, ZN => 
                           sub_126_G3_carry_8_port);
   U178 : XOR2_X1 port map( A => n36, B => sub_126_G3_carry_7_port, Z => 
                           A_neg_2_7_port);
   U179 : AND2_X1 port map( A1 => sub_126_G3_carry_6_port, A2 => n34, ZN => 
                           sub_126_G3_carry_7_port);
   U180 : XOR2_X1 port map( A => n33, B => sub_126_G3_carry_6_port, Z => 
                           A_neg_2_6_port);
   U181 : AND2_X1 port map( A1 => sub_126_G3_carry_5_port, A2 => n31, ZN => 
                           sub_126_G3_carry_6_port);
   U182 : XOR2_X1 port map( A => n30, B => sub_126_G3_carry_5_port, Z => 
                           A_neg_2_5_port);
   U183 : AND2_X1 port map( A1 => sub_126_G3_carry_4_port, A2 => n28, ZN => 
                           sub_126_G3_carry_5_port);
   U184 : XOR2_X1 port map( A => n27, B => sub_126_G3_carry_4_port, Z => 
                           A_neg_2_4_port);
   U185 : AND2_X1 port map( A1 => n19, A2 => n25, ZN => sub_126_G3_carry_4_port
                           );
   U186 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_2_3_port);
   U187 : XOR2_X1 port map( A => n66, B => sub_126_G6_carry_20_port, Z => 
                           A_neg_5_20_port);
   U188 : AND2_X1 port map( A1 => sub_126_G6_carry_19_port, A2 => n64, ZN => 
                           sub_126_G6_carry_20_port);
   U189 : XOR2_X1 port map( A => n63, B => sub_126_G6_carry_19_port, Z => 
                           A_neg_5_19_port);
   U190 : AND2_X1 port map( A1 => sub_126_G6_carry_18_port, A2 => n61, ZN => 
                           sub_126_G6_carry_19_port);
   U191 : XOR2_X1 port map( A => n60, B => sub_126_G6_carry_18_port, Z => 
                           A_neg_5_18_port);
   U192 : AND2_X1 port map( A1 => sub_126_G6_carry_17_port, A2 => n58, ZN => 
                           sub_126_G6_carry_18_port);
   U193 : XOR2_X1 port map( A => n57, B => sub_126_G6_carry_17_port, Z => 
                           A_neg_5_17_port);
   U194 : AND2_X1 port map( A1 => sub_126_G6_carry_16_port, A2 => n55, ZN => 
                           sub_126_G6_carry_17_port);
   U195 : XOR2_X1 port map( A => n54, B => sub_126_G6_carry_16_port, Z => 
                           A_neg_5_16_port);
   U196 : AND2_X1 port map( A1 => sub_126_G6_carry_15_port, A2 => n52, ZN => 
                           sub_126_G6_carry_16_port);
   U197 : XOR2_X1 port map( A => n51, B => sub_126_G6_carry_15_port, Z => 
                           A_neg_5_15_port);
   U198 : AND2_X1 port map( A1 => sub_126_G6_carry_14_port, A2 => n49, ZN => 
                           sub_126_G6_carry_15_port);
   U199 : XOR2_X1 port map( A => n48, B => sub_126_G6_carry_14_port, Z => 
                           A_neg_5_14_port);
   U200 : AND2_X1 port map( A1 => sub_126_G6_carry_13_port, A2 => n46, ZN => 
                           sub_126_G6_carry_14_port);
   U201 : XOR2_X1 port map( A => n45, B => sub_126_G6_carry_13_port, Z => 
                           A_neg_5_13_port);
   U202 : AND2_X1 port map( A1 => sub_126_G6_carry_12_port, A2 => n43, ZN => 
                           sub_126_G6_carry_13_port);
   U203 : XOR2_X1 port map( A => n42, B => sub_126_G6_carry_12_port, Z => 
                           A_neg_5_12_port);
   U204 : AND2_X1 port map( A1 => sub_126_G6_carry_11_port, A2 => n40, ZN => 
                           sub_126_G6_carry_12_port);
   U205 : XOR2_X1 port map( A => n39, B => sub_126_G6_carry_11_port, Z => 
                           A_neg_5_11_port);
   U206 : AND2_X1 port map( A1 => sub_126_G6_carry_10_port, A2 => n37, ZN => 
                           sub_126_G6_carry_11_port);
   U207 : XOR2_X1 port map( A => n36, B => sub_126_G6_carry_10_port, Z => 
                           A_neg_5_10_port);
   U208 : AND2_X1 port map( A1 => sub_126_G6_carry_9_port, A2 => n34, ZN => 
                           sub_126_G6_carry_10_port);
   U209 : XOR2_X1 port map( A => n33, B => sub_126_G6_carry_9_port, Z => 
                           A_neg_5_9_port);
   U210 : AND2_X1 port map( A1 => sub_126_G6_carry_8_port, A2 => n31, ZN => 
                           sub_126_G6_carry_9_port);
   U211 : XOR2_X1 port map( A => n30, B => sub_126_G6_carry_8_port, Z => 
                           A_neg_5_8_port);
   U212 : AND2_X1 port map( A1 => sub_126_G6_carry_7_port, A2 => n28, ZN => 
                           sub_126_G6_carry_8_port);
   U213 : XOR2_X1 port map( A => n27, B => sub_126_G6_carry_7_port, Z => 
                           A_neg_5_7_port);
   U214 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => sub_126_G6_carry_7_port
                           );
   U215 : XOR2_X1 port map( A => n24, B => n18, Z => A_neg_5_6_port);
   U216 : XOR2_X1 port map( A => n66, B => sub_126_G5_carry_19_port, Z => 
                           A_neg_4_19_port);
   U217 : AND2_X1 port map( A1 => sub_126_G5_carry_18_port, A2 => n64, ZN => 
                           sub_126_G5_carry_19_port);
   U218 : XOR2_X1 port map( A => n63, B => sub_126_G5_carry_18_port, Z => 
                           A_neg_4_18_port);
   U219 : AND2_X1 port map( A1 => sub_126_G5_carry_17_port, A2 => n61, ZN => 
                           sub_126_G5_carry_18_port);
   U220 : XOR2_X1 port map( A => n60, B => sub_126_G5_carry_17_port, Z => 
                           A_neg_4_17_port);
   U221 : AND2_X1 port map( A1 => sub_126_G5_carry_16_port, A2 => n58, ZN => 
                           sub_126_G5_carry_17_port);
   U222 : XOR2_X1 port map( A => n57, B => sub_126_G5_carry_16_port, Z => 
                           A_neg_4_16_port);
   U223 : AND2_X1 port map( A1 => sub_126_G5_carry_15_port, A2 => n55, ZN => 
                           sub_126_G5_carry_16_port);
   U224 : XOR2_X1 port map( A => n54, B => sub_126_G5_carry_15_port, Z => 
                           A_neg_4_15_port);
   U225 : AND2_X1 port map( A1 => sub_126_G5_carry_14_port, A2 => n52, ZN => 
                           sub_126_G5_carry_15_port);
   U226 : XOR2_X1 port map( A => n51, B => sub_126_G5_carry_14_port, Z => 
                           A_neg_4_14_port);
   U227 : AND2_X1 port map( A1 => sub_126_G5_carry_13_port, A2 => n49, ZN => 
                           sub_126_G5_carry_14_port);
   U228 : XOR2_X1 port map( A => n48, B => sub_126_G5_carry_13_port, Z => 
                           A_neg_4_13_port);
   U229 : AND2_X1 port map( A1 => sub_126_G5_carry_12_port, A2 => n46, ZN => 
                           sub_126_G5_carry_13_port);
   U230 : XOR2_X1 port map( A => n45, B => sub_126_G5_carry_12_port, Z => 
                           A_neg_4_12_port);
   U231 : AND2_X1 port map( A1 => sub_126_G5_carry_11_port, A2 => n43, ZN => 
                           sub_126_G5_carry_12_port);
   U232 : XOR2_X1 port map( A => n42, B => sub_126_G5_carry_11_port, Z => 
                           A_neg_4_11_port);
   U233 : AND2_X1 port map( A1 => sub_126_G5_carry_10_port, A2 => n40, ZN => 
                           sub_126_G5_carry_11_port);
   U234 : XOR2_X1 port map( A => n39, B => sub_126_G5_carry_10_port, Z => 
                           A_neg_4_10_port);
   U235 : AND2_X1 port map( A1 => sub_126_G5_carry_9_port, A2 => n37, ZN => 
                           sub_126_G5_carry_10_port);
   U236 : XOR2_X1 port map( A => n36, B => sub_126_G5_carry_9_port, Z => 
                           A_neg_4_9_port);
   U237 : AND2_X1 port map( A1 => sub_126_G5_carry_8_port, A2 => n34, ZN => 
                           sub_126_G5_carry_9_port);
   U238 : XOR2_X1 port map( A => n33, B => sub_126_G5_carry_8_port, Z => 
                           A_neg_4_8_port);
   U239 : AND2_X1 port map( A1 => sub_126_G5_carry_7_port, A2 => n31, ZN => 
                           sub_126_G5_carry_8_port);
   U240 : XOR2_X1 port map( A => n30, B => sub_126_G5_carry_7_port, Z => 
                           A_neg_4_7_port);
   U241 : AND2_X1 port map( A1 => sub_126_G5_carry_6_port, A2 => n28, ZN => 
                           sub_126_G5_carry_7_port);
   U242 : XOR2_X1 port map( A => n27, B => sub_126_G5_carry_6_port, Z => 
                           A_neg_4_6_port);
   U243 : AND2_X1 port map( A1 => n19, A2 => n25, ZN => sub_126_G5_carry_6_port
                           );
   U244 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_4_5_port);
   U245 : XOR2_X1 port map( A => n66, B => sub_126_G8_carry_22_port, Z => 
                           A_neg_7_22_port);
   U246 : AND2_X1 port map( A1 => sub_126_G8_carry_21_port, A2 => n64, ZN => 
                           sub_126_G8_carry_22_port);
   U247 : XOR2_X1 port map( A => n63, B => sub_126_G8_carry_21_port, Z => 
                           A_neg_7_21_port);
   U248 : AND2_X1 port map( A1 => sub_126_G8_carry_20_port, A2 => n61, ZN => 
                           sub_126_G8_carry_21_port);
   U249 : XOR2_X1 port map( A => n60, B => sub_126_G8_carry_20_port, Z => 
                           A_neg_7_20_port);
   U250 : AND2_X1 port map( A1 => sub_126_G8_carry_19_port, A2 => n58, ZN => 
                           sub_126_G8_carry_20_port);
   U251 : XOR2_X1 port map( A => n57, B => sub_126_G8_carry_19_port, Z => 
                           A_neg_7_19_port);
   U252 : AND2_X1 port map( A1 => sub_126_G8_carry_18_port, A2 => n55, ZN => 
                           sub_126_G8_carry_19_port);
   U253 : XOR2_X1 port map( A => n54, B => sub_126_G8_carry_18_port, Z => 
                           A_neg_7_18_port);
   U254 : AND2_X1 port map( A1 => sub_126_G8_carry_17_port, A2 => n52, ZN => 
                           sub_126_G8_carry_18_port);
   U255 : XOR2_X1 port map( A => n51, B => sub_126_G8_carry_17_port, Z => 
                           A_neg_7_17_port);
   U256 : AND2_X1 port map( A1 => sub_126_G8_carry_16_port, A2 => n49, ZN => 
                           sub_126_G8_carry_17_port);
   U257 : XOR2_X1 port map( A => n48, B => sub_126_G8_carry_16_port, Z => 
                           A_neg_7_16_port);
   U258 : AND2_X1 port map( A1 => sub_126_G8_carry_15_port, A2 => n46, ZN => 
                           sub_126_G8_carry_16_port);
   U259 : XOR2_X1 port map( A => n45, B => sub_126_G8_carry_15_port, Z => 
                           A_neg_7_15_port);
   U260 : AND2_X1 port map( A1 => sub_126_G8_carry_14_port, A2 => n43, ZN => 
                           sub_126_G8_carry_15_port);
   U261 : XOR2_X1 port map( A => n42, B => sub_126_G8_carry_14_port, Z => 
                           A_neg_7_14_port);
   U262 : AND2_X1 port map( A1 => sub_126_G8_carry_13_port, A2 => n40, ZN => 
                           sub_126_G8_carry_14_port);
   U263 : XOR2_X1 port map( A => n39, B => sub_126_G8_carry_13_port, Z => 
                           A_neg_7_13_port);
   U264 : AND2_X1 port map( A1 => sub_126_G8_carry_12_port, A2 => n37, ZN => 
                           sub_126_G8_carry_13_port);
   U265 : XOR2_X1 port map( A => n36, B => sub_126_G8_carry_12_port, Z => 
                           A_neg_7_12_port);
   U266 : AND2_X1 port map( A1 => sub_126_G8_carry_11_port, A2 => n34, ZN => 
                           sub_126_G8_carry_12_port);
   U267 : XOR2_X1 port map( A => n33, B => sub_126_G8_carry_11_port, Z => 
                           A_neg_7_11_port);
   U268 : AND2_X1 port map( A1 => sub_126_G8_carry_10_port, A2 => n31, ZN => 
                           sub_126_G8_carry_11_port);
   U269 : XOR2_X1 port map( A => n30, B => sub_126_G8_carry_10_port, Z => 
                           A_neg_7_10_port);
   U270 : AND2_X1 port map( A1 => sub_126_G8_carry_9_port, A2 => n28, ZN => 
                           sub_126_G8_carry_10_port);
   U271 : XOR2_X1 port map( A => n27, B => sub_126_G8_carry_9_port, Z => 
                           A_neg_7_9_port);
   U272 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => sub_126_G8_carry_9_port
                           );
   U273 : XOR2_X1 port map( A => n24, B => n18, Z => A_neg_7_8_port);
   U274 : XOR2_X1 port map( A => n66, B => sub_126_G7_carry_21_port, Z => 
                           A_neg_6_21_port);
   U275 : AND2_X1 port map( A1 => sub_126_G7_carry_20_port, A2 => n64, ZN => 
                           sub_126_G7_carry_21_port);
   U276 : XOR2_X1 port map( A => n63, B => sub_126_G7_carry_20_port, Z => 
                           A_neg_6_20_port);
   U277 : AND2_X1 port map( A1 => sub_126_G7_carry_19_port, A2 => n61, ZN => 
                           sub_126_G7_carry_20_port);
   U278 : XOR2_X1 port map( A => n60, B => sub_126_G7_carry_19_port, Z => 
                           A_neg_6_19_port);
   U279 : AND2_X1 port map( A1 => sub_126_G7_carry_18_port, A2 => n58, ZN => 
                           sub_126_G7_carry_19_port);
   U280 : XOR2_X1 port map( A => n57, B => sub_126_G7_carry_18_port, Z => 
                           A_neg_6_18_port);
   U281 : AND2_X1 port map( A1 => sub_126_G7_carry_17_port, A2 => n55, ZN => 
                           sub_126_G7_carry_18_port);
   U282 : XOR2_X1 port map( A => n54, B => sub_126_G7_carry_17_port, Z => 
                           A_neg_6_17_port);
   U283 : AND2_X1 port map( A1 => sub_126_G7_carry_16_port, A2 => n52, ZN => 
                           sub_126_G7_carry_17_port);
   U284 : XOR2_X1 port map( A => n51, B => sub_126_G7_carry_16_port, Z => 
                           A_neg_6_16_port);
   U285 : AND2_X1 port map( A1 => sub_126_G7_carry_15_port, A2 => n49, ZN => 
                           sub_126_G7_carry_16_port);
   U286 : XOR2_X1 port map( A => n48, B => sub_126_G7_carry_15_port, Z => 
                           A_neg_6_15_port);
   U287 : AND2_X1 port map( A1 => sub_126_G7_carry_14_port, A2 => n46, ZN => 
                           sub_126_G7_carry_15_port);
   U288 : XOR2_X1 port map( A => n45, B => sub_126_G7_carry_14_port, Z => 
                           A_neg_6_14_port);
   U289 : AND2_X1 port map( A1 => sub_126_G7_carry_13_port, A2 => n43, ZN => 
                           sub_126_G7_carry_14_port);
   U290 : XOR2_X1 port map( A => n42, B => sub_126_G7_carry_13_port, Z => 
                           A_neg_6_13_port);
   U291 : AND2_X1 port map( A1 => sub_126_G7_carry_12_port, A2 => n40, ZN => 
                           sub_126_G7_carry_13_port);
   U292 : XOR2_X1 port map( A => n39, B => sub_126_G7_carry_12_port, Z => 
                           A_neg_6_12_port);
   U293 : AND2_X1 port map( A1 => sub_126_G7_carry_11_port, A2 => n37, ZN => 
                           sub_126_G7_carry_12_port);
   U294 : XOR2_X1 port map( A => n36, B => sub_126_G7_carry_11_port, Z => 
                           A_neg_6_11_port);
   U295 : AND2_X1 port map( A1 => sub_126_G7_carry_10_port, A2 => n34, ZN => 
                           sub_126_G7_carry_11_port);
   U296 : XOR2_X1 port map( A => n33, B => sub_126_G7_carry_10_port, Z => 
                           A_neg_6_10_port);
   U297 : AND2_X1 port map( A1 => sub_126_G7_carry_9_port, A2 => n31, ZN => 
                           sub_126_G7_carry_10_port);
   U298 : XOR2_X1 port map( A => n30, B => sub_126_G7_carry_9_port, Z => 
                           A_neg_6_9_port);
   U299 : AND2_X1 port map( A1 => sub_126_G7_carry_8_port, A2 => n28, ZN => 
                           sub_126_G7_carry_9_port);
   U300 : XOR2_X1 port map( A => n27, B => sub_126_G7_carry_8_port, Z => 
                           A_neg_6_8_port);
   U301 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => sub_126_G7_carry_8_port
                           );
   U302 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_6_7_port);
   U303 : XOR2_X1 port map( A => n66, B => sub_126_G10_carry_24_port, Z => 
                           A_neg_9_24_port);
   U304 : AND2_X1 port map( A1 => sub_126_G10_carry_23_port, A2 => n64, ZN => 
                           sub_126_G10_carry_24_port);
   U305 : XOR2_X1 port map( A => n63, B => sub_126_G10_carry_23_port, Z => 
                           A_neg_9_23_port);
   U306 : AND2_X1 port map( A1 => sub_126_G10_carry_22_port, A2 => n61, ZN => 
                           sub_126_G10_carry_23_port);
   U307 : XOR2_X1 port map( A => n60, B => sub_126_G10_carry_22_port, Z => 
                           A_neg_9_22_port);
   U308 : AND2_X1 port map( A1 => sub_126_G10_carry_21_port, A2 => n58, ZN => 
                           sub_126_G10_carry_22_port);
   U309 : XOR2_X1 port map( A => n57, B => sub_126_G10_carry_21_port, Z => 
                           A_neg_9_21_port);
   U310 : AND2_X1 port map( A1 => sub_126_G10_carry_20_port, A2 => n55, ZN => 
                           sub_126_G10_carry_21_port);
   U311 : XOR2_X1 port map( A => n54, B => sub_126_G10_carry_20_port, Z => 
                           A_neg_9_20_port);
   U312 : AND2_X1 port map( A1 => sub_126_G10_carry_19_port, A2 => n52, ZN => 
                           sub_126_G10_carry_20_port);
   U313 : XOR2_X1 port map( A => n51, B => sub_126_G10_carry_19_port, Z => 
                           A_neg_9_19_port);
   U314 : AND2_X1 port map( A1 => sub_126_G10_carry_18_port, A2 => n49, ZN => 
                           sub_126_G10_carry_19_port);
   U315 : XOR2_X1 port map( A => n48, B => sub_126_G10_carry_18_port, Z => 
                           A_neg_9_18_port);
   U316 : AND2_X1 port map( A1 => sub_126_G10_carry_17_port, A2 => n46, ZN => 
                           sub_126_G10_carry_18_port);
   U317 : XOR2_X1 port map( A => n45, B => sub_126_G10_carry_17_port, Z => 
                           A_neg_9_17_port);
   U318 : AND2_X1 port map( A1 => sub_126_G10_carry_16_port, A2 => n43, ZN => 
                           sub_126_G10_carry_17_port);
   U319 : XOR2_X1 port map( A => n42, B => sub_126_G10_carry_16_port, Z => 
                           A_neg_9_16_port);
   U320 : AND2_X1 port map( A1 => sub_126_G10_carry_15_port, A2 => n40, ZN => 
                           sub_126_G10_carry_16_port);
   U321 : XOR2_X1 port map( A => n39, B => sub_126_G10_carry_15_port, Z => 
                           A_neg_9_15_port);
   U322 : AND2_X1 port map( A1 => sub_126_G10_carry_14_port, A2 => n37, ZN => 
                           sub_126_G10_carry_15_port);
   U323 : XOR2_X1 port map( A => n36, B => sub_126_G10_carry_14_port, Z => 
                           A_neg_9_14_port);
   U324 : AND2_X1 port map( A1 => sub_126_G10_carry_13_port, A2 => n34, ZN => 
                           sub_126_G10_carry_14_port);
   U325 : XOR2_X1 port map( A => n33, B => sub_126_G10_carry_13_port, Z => 
                           A_neg_9_13_port);
   U326 : AND2_X1 port map( A1 => sub_126_G10_carry_12_port, A2 => n31, ZN => 
                           sub_126_G10_carry_13_port);
   U327 : XOR2_X1 port map( A => n30, B => sub_126_G10_carry_12_port, Z => 
                           A_neg_9_12_port);
   U328 : AND2_X1 port map( A1 => sub_126_G10_carry_11_port, A2 => n28, ZN => 
                           sub_126_G10_carry_12_port);
   U329 : XOR2_X1 port map( A => n27, B => sub_126_G10_carry_11_port, Z => 
                           A_neg_9_11_port);
   U330 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G10_carry_11_port);
   U331 : XOR2_X1 port map( A => n24, B => n18, Z => A_neg_9_10_port);
   U332 : XOR2_X1 port map( A => n66, B => sub_126_G9_carry_23_port, Z => 
                           A_neg_8_23_port);
   U333 : AND2_X1 port map( A1 => sub_126_G9_carry_22_port, A2 => n64, ZN => 
                           sub_126_G9_carry_23_port);
   U334 : XOR2_X1 port map( A => n63, B => sub_126_G9_carry_22_port, Z => 
                           A_neg_8_22_port);
   U335 : AND2_X1 port map( A1 => sub_126_G9_carry_21_port, A2 => n61, ZN => 
                           sub_126_G9_carry_22_port);
   U336 : XOR2_X1 port map( A => n60, B => sub_126_G9_carry_21_port, Z => 
                           A_neg_8_21_port);
   U337 : AND2_X1 port map( A1 => sub_126_G9_carry_20_port, A2 => n58, ZN => 
                           sub_126_G9_carry_21_port);
   U338 : XOR2_X1 port map( A => n57, B => sub_126_G9_carry_20_port, Z => 
                           A_neg_8_20_port);
   U339 : AND2_X1 port map( A1 => sub_126_G9_carry_19_port, A2 => n55, ZN => 
                           sub_126_G9_carry_20_port);
   U340 : XOR2_X1 port map( A => n54, B => sub_126_G9_carry_19_port, Z => 
                           A_neg_8_19_port);
   U341 : AND2_X1 port map( A1 => sub_126_G9_carry_18_port, A2 => n52, ZN => 
                           sub_126_G9_carry_19_port);
   U342 : XOR2_X1 port map( A => n51, B => sub_126_G9_carry_18_port, Z => 
                           A_neg_8_18_port);
   U343 : AND2_X1 port map( A1 => sub_126_G9_carry_17_port, A2 => n49, ZN => 
                           sub_126_G9_carry_18_port);
   U344 : XOR2_X1 port map( A => n48, B => sub_126_G9_carry_17_port, Z => 
                           A_neg_8_17_port);
   U345 : AND2_X1 port map( A1 => sub_126_G9_carry_16_port, A2 => n46, ZN => 
                           sub_126_G9_carry_17_port);
   U346 : XOR2_X1 port map( A => n45, B => sub_126_G9_carry_16_port, Z => 
                           A_neg_8_16_port);
   U347 : AND2_X1 port map( A1 => sub_126_G9_carry_15_port, A2 => n43, ZN => 
                           sub_126_G9_carry_16_port);
   U348 : XOR2_X1 port map( A => n42, B => sub_126_G9_carry_15_port, Z => 
                           A_neg_8_15_port);
   U349 : AND2_X1 port map( A1 => sub_126_G9_carry_14_port, A2 => n40, ZN => 
                           sub_126_G9_carry_15_port);
   U350 : XOR2_X1 port map( A => n39, B => sub_126_G9_carry_14_port, Z => 
                           A_neg_8_14_port);
   U351 : AND2_X1 port map( A1 => sub_126_G9_carry_13_port, A2 => n37, ZN => 
                           sub_126_G9_carry_14_port);
   U352 : XOR2_X1 port map( A => n36, B => sub_126_G9_carry_13_port, Z => 
                           A_neg_8_13_port);
   U353 : AND2_X1 port map( A1 => sub_126_G9_carry_12_port, A2 => n34, ZN => 
                           sub_126_G9_carry_13_port);
   U354 : XOR2_X1 port map( A => n33, B => sub_126_G9_carry_12_port, Z => 
                           A_neg_8_12_port);
   U355 : AND2_X1 port map( A1 => sub_126_G9_carry_11_port, A2 => n31, ZN => 
                           sub_126_G9_carry_12_port);
   U356 : XOR2_X1 port map( A => n30, B => sub_126_G9_carry_11_port, Z => 
                           A_neg_8_11_port);
   U357 : AND2_X1 port map( A1 => sub_126_G9_carry_10_port, A2 => n28, ZN => 
                           sub_126_G9_carry_11_port);
   U358 : XOR2_X1 port map( A => n27, B => sub_126_G9_carry_10_port, Z => 
                           A_neg_8_10_port);
   U359 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G9_carry_10_port);
   U360 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_8_9_port);
   U361 : XOR2_X1 port map( A => n66, B => sub_126_G12_carry_26_port, Z => 
                           A_neg_11_26_port);
   U362 : AND2_X1 port map( A1 => sub_126_G12_carry_25_port, A2 => n64, ZN => 
                           sub_126_G12_carry_26_port);
   U363 : XOR2_X1 port map( A => n63, B => sub_126_G12_carry_25_port, Z => 
                           A_neg_11_25_port);
   U364 : AND2_X1 port map( A1 => sub_126_G12_carry_24_port, A2 => n61, ZN => 
                           sub_126_G12_carry_25_port);
   U365 : XOR2_X1 port map( A => n60, B => sub_126_G12_carry_24_port, Z => 
                           A_neg_11_24_port);
   U366 : AND2_X1 port map( A1 => sub_126_G12_carry_23_port, A2 => n58, ZN => 
                           sub_126_G12_carry_24_port);
   U367 : XOR2_X1 port map( A => n57, B => sub_126_G12_carry_23_port, Z => 
                           A_neg_11_23_port);
   U368 : AND2_X1 port map( A1 => sub_126_G12_carry_22_port, A2 => n55, ZN => 
                           sub_126_G12_carry_23_port);
   U369 : XOR2_X1 port map( A => n54, B => sub_126_G12_carry_22_port, Z => 
                           A_neg_11_22_port);
   U370 : AND2_X1 port map( A1 => sub_126_G12_carry_21_port, A2 => n52, ZN => 
                           sub_126_G12_carry_22_port);
   U371 : XOR2_X1 port map( A => n51, B => sub_126_G12_carry_21_port, Z => 
                           A_neg_11_21_port);
   U372 : AND2_X1 port map( A1 => sub_126_G12_carry_20_port, A2 => n49, ZN => 
                           sub_126_G12_carry_21_port);
   U373 : XOR2_X1 port map( A => n48, B => sub_126_G12_carry_20_port, Z => 
                           A_neg_11_20_port);
   U374 : AND2_X1 port map( A1 => sub_126_G12_carry_19_port, A2 => n46, ZN => 
                           sub_126_G12_carry_20_port);
   U375 : XOR2_X1 port map( A => n45, B => sub_126_G12_carry_19_port, Z => 
                           A_neg_11_19_port);
   U376 : AND2_X1 port map( A1 => sub_126_G12_carry_18_port, A2 => n43, ZN => 
                           sub_126_G12_carry_19_port);
   U377 : XOR2_X1 port map( A => n42, B => sub_126_G12_carry_18_port, Z => 
                           A_neg_11_18_port);
   U378 : AND2_X1 port map( A1 => sub_126_G12_carry_17_port, A2 => n40, ZN => 
                           sub_126_G12_carry_18_port);
   U379 : XOR2_X1 port map( A => n39, B => sub_126_G12_carry_17_port, Z => 
                           A_neg_11_17_port);
   U380 : AND2_X1 port map( A1 => sub_126_G12_carry_16_port, A2 => n37, ZN => 
                           sub_126_G12_carry_17_port);
   U381 : XOR2_X1 port map( A => n36, B => sub_126_G12_carry_16_port, Z => 
                           A_neg_11_16_port);
   U382 : AND2_X1 port map( A1 => sub_126_G12_carry_15_port, A2 => n34, ZN => 
                           sub_126_G12_carry_16_port);
   U383 : XOR2_X1 port map( A => n33, B => sub_126_G12_carry_15_port, Z => 
                           A_neg_11_15_port);
   U384 : AND2_X1 port map( A1 => sub_126_G12_carry_14_port, A2 => n31, ZN => 
                           sub_126_G12_carry_15_port);
   U385 : XOR2_X1 port map( A => n30, B => sub_126_G12_carry_14_port, Z => 
                           A_neg_11_14_port);
   U386 : AND2_X1 port map( A1 => sub_126_G12_carry_13_port, A2 => n28, ZN => 
                           sub_126_G12_carry_14_port);
   U387 : XOR2_X1 port map( A => n27, B => sub_126_G12_carry_13_port, Z => 
                           A_neg_11_13_port);
   U388 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G12_carry_13_port);
   U389 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_11_12_port);
   U390 : XOR2_X1 port map( A => n66, B => sub_126_G11_carry_25_port, Z => 
                           A_neg_10_25_port);
   U391 : AND2_X1 port map( A1 => sub_126_G11_carry_24_port, A2 => n64, ZN => 
                           sub_126_G11_carry_25_port);
   U392 : XOR2_X1 port map( A => n63, B => sub_126_G11_carry_24_port, Z => 
                           A_neg_10_24_port);
   U393 : AND2_X1 port map( A1 => sub_126_G11_carry_23_port, A2 => n61, ZN => 
                           sub_126_G11_carry_24_port);
   U394 : XOR2_X1 port map( A => n60, B => sub_126_G11_carry_23_port, Z => 
                           A_neg_10_23_port);
   U395 : AND2_X1 port map( A1 => sub_126_G11_carry_22_port, A2 => n58, ZN => 
                           sub_126_G11_carry_23_port);
   U396 : XOR2_X1 port map( A => n57, B => sub_126_G11_carry_22_port, Z => 
                           A_neg_10_22_port);
   U397 : AND2_X1 port map( A1 => sub_126_G11_carry_21_port, A2 => n55, ZN => 
                           sub_126_G11_carry_22_port);
   U398 : XOR2_X1 port map( A => n54, B => sub_126_G11_carry_21_port, Z => 
                           A_neg_10_21_port);
   U399 : AND2_X1 port map( A1 => sub_126_G11_carry_20_port, A2 => n52, ZN => 
                           sub_126_G11_carry_21_port);
   U400 : XOR2_X1 port map( A => n51, B => sub_126_G11_carry_20_port, Z => 
                           A_neg_10_20_port);
   U401 : AND2_X1 port map( A1 => sub_126_G11_carry_19_port, A2 => n49, ZN => 
                           sub_126_G11_carry_20_port);
   U402 : XOR2_X1 port map( A => n48, B => sub_126_G11_carry_19_port, Z => 
                           A_neg_10_19_port);
   U403 : AND2_X1 port map( A1 => sub_126_G11_carry_18_port, A2 => n46, ZN => 
                           sub_126_G11_carry_19_port);
   U404 : XOR2_X1 port map( A => n45, B => sub_126_G11_carry_18_port, Z => 
                           A_neg_10_18_port);
   U405 : AND2_X1 port map( A1 => sub_126_G11_carry_17_port, A2 => n43, ZN => 
                           sub_126_G11_carry_18_port);
   U406 : XOR2_X1 port map( A => n42, B => sub_126_G11_carry_17_port, Z => 
                           A_neg_10_17_port);
   U407 : AND2_X1 port map( A1 => sub_126_G11_carry_16_port, A2 => n40, ZN => 
                           sub_126_G11_carry_17_port);
   U408 : XOR2_X1 port map( A => n39, B => sub_126_G11_carry_16_port, Z => 
                           A_neg_10_16_port);
   U409 : AND2_X1 port map( A1 => sub_126_G11_carry_15_port, A2 => n37, ZN => 
                           sub_126_G11_carry_16_port);
   U410 : XOR2_X1 port map( A => n36, B => sub_126_G11_carry_15_port, Z => 
                           A_neg_10_15_port);
   U411 : AND2_X1 port map( A1 => sub_126_G11_carry_14_port, A2 => n34, ZN => 
                           sub_126_G11_carry_15_port);
   U412 : XOR2_X1 port map( A => n33, B => sub_126_G11_carry_14_port, Z => 
                           A_neg_10_14_port);
   U413 : AND2_X1 port map( A1 => sub_126_G11_carry_13_port, A2 => n31, ZN => 
                           sub_126_G11_carry_14_port);
   U414 : XOR2_X1 port map( A => n30, B => sub_126_G11_carry_13_port, Z => 
                           A_neg_10_13_port);
   U415 : AND2_X1 port map( A1 => sub_126_G11_carry_12_port, A2 => n28, ZN => 
                           sub_126_G11_carry_13_port);
   U416 : XOR2_X1 port map( A => n27, B => sub_126_G11_carry_12_port, Z => 
                           A_neg_10_12_port);
   U417 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G11_carry_12_port);
   U418 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_10_11_port);
   U419 : XOR2_X1 port map( A => n66, B => sub_126_G14_carry_28_port, Z => 
                           A_neg_13_28_port);
   U420 : AND2_X1 port map( A1 => sub_126_G14_carry_27_port, A2 => n64, ZN => 
                           sub_126_G14_carry_28_port);
   U421 : XOR2_X1 port map( A => n63, B => sub_126_G14_carry_27_port, Z => 
                           A_neg_13_27_port);
   U422 : AND2_X1 port map( A1 => sub_126_G14_carry_26_port, A2 => n61, ZN => 
                           sub_126_G14_carry_27_port);
   U423 : XOR2_X1 port map( A => n60, B => sub_126_G14_carry_26_port, Z => 
                           A_neg_13_26_port);
   U424 : AND2_X1 port map( A1 => sub_126_G14_carry_25_port, A2 => n58, ZN => 
                           sub_126_G14_carry_26_port);
   U425 : XOR2_X1 port map( A => n57, B => sub_126_G14_carry_25_port, Z => 
                           A_neg_13_25_port);
   U426 : AND2_X1 port map( A1 => sub_126_G14_carry_24_port, A2 => n55, ZN => 
                           sub_126_G14_carry_25_port);
   U427 : XOR2_X1 port map( A => n54, B => sub_126_G14_carry_24_port, Z => 
                           A_neg_13_24_port);
   U428 : AND2_X1 port map( A1 => sub_126_G14_carry_23_port, A2 => n52, ZN => 
                           sub_126_G14_carry_24_port);
   U429 : XOR2_X1 port map( A => n51, B => sub_126_G14_carry_23_port, Z => 
                           A_neg_13_23_port);
   U430 : AND2_X1 port map( A1 => sub_126_G14_carry_22_port, A2 => n49, ZN => 
                           sub_126_G14_carry_23_port);
   U431 : XOR2_X1 port map( A => n48, B => sub_126_G14_carry_22_port, Z => 
                           A_neg_13_22_port);
   U432 : AND2_X1 port map( A1 => sub_126_G14_carry_21_port, A2 => n46, ZN => 
                           sub_126_G14_carry_22_port);
   U433 : XOR2_X1 port map( A => n45, B => sub_126_G14_carry_21_port, Z => 
                           A_neg_13_21_port);
   U434 : AND2_X1 port map( A1 => sub_126_G14_carry_20_port, A2 => n43, ZN => 
                           sub_126_G14_carry_21_port);
   U435 : XOR2_X1 port map( A => n42, B => sub_126_G14_carry_20_port, Z => 
                           A_neg_13_20_port);
   U436 : AND2_X1 port map( A1 => sub_126_G14_carry_19_port, A2 => n40, ZN => 
                           sub_126_G14_carry_20_port);
   U437 : XOR2_X1 port map( A => n39, B => sub_126_G14_carry_19_port, Z => 
                           A_neg_13_19_port);
   U438 : AND2_X1 port map( A1 => sub_126_G14_carry_18_port, A2 => n37, ZN => 
                           sub_126_G14_carry_19_port);
   U439 : XOR2_X1 port map( A => n36, B => sub_126_G14_carry_18_port, Z => 
                           A_neg_13_18_port);
   U440 : AND2_X1 port map( A1 => sub_126_G14_carry_17_port, A2 => n34, ZN => 
                           sub_126_G14_carry_18_port);
   U441 : XOR2_X1 port map( A => n33, B => sub_126_G14_carry_17_port, Z => 
                           A_neg_13_17_port);
   U442 : AND2_X1 port map( A1 => sub_126_G14_carry_16_port, A2 => n31, ZN => 
                           sub_126_G14_carry_17_port);
   U443 : XOR2_X1 port map( A => n30, B => sub_126_G14_carry_16_port, Z => 
                           A_neg_13_16_port);
   U444 : AND2_X1 port map( A1 => sub_126_G14_carry_15_port, A2 => n28, ZN => 
                           sub_126_G14_carry_16_port);
   U445 : XOR2_X1 port map( A => n27, B => sub_126_G14_carry_15_port, Z => 
                           A_neg_13_15_port);
   U446 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G14_carry_15_port);
   U447 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_13_14_port);
   U448 : XOR2_X1 port map( A => n66, B => sub_126_G13_carry_27_port, Z => 
                           A_neg_12_27_port);
   U449 : AND2_X1 port map( A1 => sub_126_G13_carry_26_port, A2 => n64, ZN => 
                           sub_126_G13_carry_27_port);
   U450 : XOR2_X1 port map( A => n63, B => sub_126_G13_carry_26_port, Z => 
                           A_neg_12_26_port);
   U451 : AND2_X1 port map( A1 => sub_126_G13_carry_25_port, A2 => n61, ZN => 
                           sub_126_G13_carry_26_port);
   U452 : XOR2_X1 port map( A => n60, B => sub_126_G13_carry_25_port, Z => 
                           A_neg_12_25_port);
   U453 : AND2_X1 port map( A1 => sub_126_G13_carry_24_port, A2 => n58, ZN => 
                           sub_126_G13_carry_25_port);
   U454 : XOR2_X1 port map( A => n57, B => sub_126_G13_carry_24_port, Z => 
                           A_neg_12_24_port);
   U455 : AND2_X1 port map( A1 => sub_126_G13_carry_23_port, A2 => n55, ZN => 
                           sub_126_G13_carry_24_port);
   U456 : XOR2_X1 port map( A => n54, B => sub_126_G13_carry_23_port, Z => 
                           A_neg_12_23_port);
   U457 : AND2_X1 port map( A1 => sub_126_G13_carry_22_port, A2 => n52, ZN => 
                           sub_126_G13_carry_23_port);
   U458 : XOR2_X1 port map( A => n51, B => sub_126_G13_carry_22_port, Z => 
                           A_neg_12_22_port);
   U459 : AND2_X1 port map( A1 => sub_126_G13_carry_21_port, A2 => n49, ZN => 
                           sub_126_G13_carry_22_port);
   U460 : XOR2_X1 port map( A => n48, B => sub_126_G13_carry_21_port, Z => 
                           A_neg_12_21_port);
   U461 : AND2_X1 port map( A1 => sub_126_G13_carry_20_port, A2 => n46, ZN => 
                           sub_126_G13_carry_21_port);
   U462 : XOR2_X1 port map( A => n45, B => sub_126_G13_carry_20_port, Z => 
                           A_neg_12_20_port);
   U463 : AND2_X1 port map( A1 => sub_126_G13_carry_19_port, A2 => n43, ZN => 
                           sub_126_G13_carry_20_port);
   U464 : XOR2_X1 port map( A => n42, B => sub_126_G13_carry_19_port, Z => 
                           A_neg_12_19_port);
   U465 : AND2_X1 port map( A1 => sub_126_G13_carry_18_port, A2 => n40, ZN => 
                           sub_126_G13_carry_19_port);
   U466 : XOR2_X1 port map( A => n39, B => sub_126_G13_carry_18_port, Z => 
                           A_neg_12_18_port);
   U467 : AND2_X1 port map( A1 => sub_126_G13_carry_17_port, A2 => n37, ZN => 
                           sub_126_G13_carry_18_port);
   U468 : XOR2_X1 port map( A => n36, B => sub_126_G13_carry_17_port, Z => 
                           A_neg_12_17_port);
   U469 : AND2_X1 port map( A1 => sub_126_G13_carry_16_port, A2 => n34, ZN => 
                           sub_126_G13_carry_17_port);
   U470 : XOR2_X1 port map( A => n33, B => sub_126_G13_carry_16_port, Z => 
                           A_neg_12_16_port);
   U471 : AND2_X1 port map( A1 => sub_126_G13_carry_15_port, A2 => n31, ZN => 
                           sub_126_G13_carry_16_port);
   U472 : XOR2_X1 port map( A => n30, B => sub_126_G13_carry_15_port, Z => 
                           A_neg_12_15_port);
   U473 : AND2_X1 port map( A1 => sub_126_G13_carry_14_port, A2 => n28, ZN => 
                           sub_126_G13_carry_15_port);
   U474 : XOR2_X1 port map( A => n27, B => sub_126_G13_carry_14_port, Z => 
                           A_neg_12_14_port);
   U475 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G13_carry_14_port);
   U476 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_12_13_port);
   U477 : XOR2_X1 port map( A => n66, B => sub_126_G16_carry_30_port, Z => 
                           A_neg_15_30_port);
   U478 : AND2_X1 port map( A1 => sub_126_G16_carry_29_port, A2 => n64, ZN => 
                           sub_126_G16_carry_30_port);
   U479 : XOR2_X1 port map( A => n63, B => sub_126_G16_carry_29_port, Z => 
                           A_neg_15_29_port);
   U480 : AND2_X1 port map( A1 => sub_126_G16_carry_28_port, A2 => n61, ZN => 
                           sub_126_G16_carry_29_port);
   U481 : XOR2_X1 port map( A => n60, B => sub_126_G16_carry_28_port, Z => 
                           A_neg_15_28_port);
   U482 : AND2_X1 port map( A1 => sub_126_G16_carry_27_port, A2 => n58, ZN => 
                           sub_126_G16_carry_28_port);
   U483 : XOR2_X1 port map( A => n57, B => sub_126_G16_carry_27_port, Z => 
                           A_neg_15_27_port);
   U484 : AND2_X1 port map( A1 => sub_126_G16_carry_26_port, A2 => n55, ZN => 
                           sub_126_G16_carry_27_port);
   U485 : XOR2_X1 port map( A => n54, B => sub_126_G16_carry_26_port, Z => 
                           A_neg_15_26_port);
   U486 : AND2_X1 port map( A1 => sub_126_G16_carry_25_port, A2 => n52, ZN => 
                           sub_126_G16_carry_26_port);
   U487 : XOR2_X1 port map( A => n51, B => sub_126_G16_carry_25_port, Z => 
                           A_neg_15_25_port);
   U488 : AND2_X1 port map( A1 => sub_126_G16_carry_24_port, A2 => n49, ZN => 
                           sub_126_G16_carry_25_port);
   U489 : XOR2_X1 port map( A => n48, B => sub_126_G16_carry_24_port, Z => 
                           A_neg_15_24_port);
   U490 : AND2_X1 port map( A1 => sub_126_G16_carry_23_port, A2 => n46, ZN => 
                           sub_126_G16_carry_24_port);
   U491 : XOR2_X1 port map( A => n45, B => sub_126_G16_carry_23_port, Z => 
                           A_neg_15_23_port);
   U492 : AND2_X1 port map( A1 => sub_126_G16_carry_22_port, A2 => n43, ZN => 
                           sub_126_G16_carry_23_port);
   U493 : XOR2_X1 port map( A => n42, B => sub_126_G16_carry_22_port, Z => 
                           A_neg_15_22_port);
   U494 : AND2_X1 port map( A1 => sub_126_G16_carry_21_port, A2 => n40, ZN => 
                           sub_126_G16_carry_22_port);
   U495 : XOR2_X1 port map( A => n39, B => sub_126_G16_carry_21_port, Z => 
                           A_neg_15_21_port);
   U496 : AND2_X1 port map( A1 => sub_126_G16_carry_20_port, A2 => n37, ZN => 
                           sub_126_G16_carry_21_port);
   U497 : XOR2_X1 port map( A => n36, B => sub_126_G16_carry_20_port, Z => 
                           A_neg_15_20_port);
   U498 : AND2_X1 port map( A1 => sub_126_G16_carry_19_port, A2 => n34, ZN => 
                           sub_126_G16_carry_20_port);
   U499 : XOR2_X1 port map( A => n33, B => sub_126_G16_carry_19_port, Z => 
                           A_neg_15_19_port);
   U500 : AND2_X1 port map( A1 => sub_126_G16_carry_18_port, A2 => n31, ZN => 
                           sub_126_G16_carry_19_port);
   U501 : XOR2_X1 port map( A => n30, B => sub_126_G16_carry_18_port, Z => 
                           A_neg_15_18_port);
   U502 : AND2_X1 port map( A1 => sub_126_G16_carry_17_port, A2 => n28, ZN => 
                           sub_126_G16_carry_18_port);
   U503 : XOR2_X1 port map( A => n27, B => sub_126_G16_carry_17_port, Z => 
                           A_neg_15_17_port);
   U504 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G16_carry_17_port);
   U505 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_15_16_port);
   U506 : XOR2_X1 port map( A => n66, B => sub_126_G15_carry_29_port, Z => 
                           A_neg_14_29_port);
   U507 : AND2_X1 port map( A1 => sub_126_G15_carry_28_port, A2 => n64, ZN => 
                           sub_126_G15_carry_29_port);
   U508 : XOR2_X1 port map( A => n63, B => sub_126_G15_carry_28_port, Z => 
                           A_neg_14_28_port);
   U509 : AND2_X1 port map( A1 => sub_126_G15_carry_27_port, A2 => n61, ZN => 
                           sub_126_G15_carry_28_port);
   U510 : XOR2_X1 port map( A => n60, B => sub_126_G15_carry_27_port, Z => 
                           A_neg_14_27_port);
   U511 : AND2_X1 port map( A1 => sub_126_G15_carry_26_port, A2 => n58, ZN => 
                           sub_126_G15_carry_27_port);
   U512 : XOR2_X1 port map( A => n57, B => sub_126_G15_carry_26_port, Z => 
                           A_neg_14_26_port);
   U513 : AND2_X1 port map( A1 => sub_126_G15_carry_25_port, A2 => n55, ZN => 
                           sub_126_G15_carry_26_port);
   U514 : XOR2_X1 port map( A => n54, B => sub_126_G15_carry_25_port, Z => 
                           A_neg_14_25_port);
   U515 : AND2_X1 port map( A1 => sub_126_G15_carry_24_port, A2 => n52, ZN => 
                           sub_126_G15_carry_25_port);
   U516 : XOR2_X1 port map( A => n51, B => sub_126_G15_carry_24_port, Z => 
                           A_neg_14_24_port);
   U517 : AND2_X1 port map( A1 => sub_126_G15_carry_23_port, A2 => n49, ZN => 
                           sub_126_G15_carry_24_port);
   U518 : XOR2_X1 port map( A => n48, B => sub_126_G15_carry_23_port, Z => 
                           A_neg_14_23_port);
   U519 : AND2_X1 port map( A1 => sub_126_G15_carry_22_port, A2 => n46, ZN => 
                           sub_126_G15_carry_23_port);
   U520 : XOR2_X1 port map( A => n45, B => sub_126_G15_carry_22_port, Z => 
                           A_neg_14_22_port);
   U521 : AND2_X1 port map( A1 => sub_126_G15_carry_21_port, A2 => n43, ZN => 
                           sub_126_G15_carry_22_port);
   U522 : XOR2_X1 port map( A => n42, B => sub_126_G15_carry_21_port, Z => 
                           A_neg_14_21_port);
   U523 : AND2_X1 port map( A1 => sub_126_G15_carry_20_port, A2 => n40, ZN => 
                           sub_126_G15_carry_21_port);
   U524 : XOR2_X1 port map( A => n39, B => sub_126_G15_carry_20_port, Z => 
                           A_neg_14_20_port);
   U525 : AND2_X1 port map( A1 => sub_126_G15_carry_19_port, A2 => n37, ZN => 
                           sub_126_G15_carry_20_port);
   U526 : XOR2_X1 port map( A => n36, B => sub_126_G15_carry_19_port, Z => 
                           A_neg_14_19_port);
   U527 : AND2_X1 port map( A1 => sub_126_G15_carry_18_port, A2 => n34, ZN => 
                           sub_126_G15_carry_19_port);
   U528 : XOR2_X1 port map( A => n33, B => sub_126_G15_carry_18_port, Z => 
                           A_neg_14_18_port);
   U529 : AND2_X1 port map( A1 => sub_126_G15_carry_17_port, A2 => n31, ZN => 
                           sub_126_G15_carry_18_port);
   U530 : XOR2_X1 port map( A => n30, B => sub_126_G15_carry_17_port, Z => 
                           A_neg_14_17_port);
   U531 : AND2_X1 port map( A1 => sub_126_G15_carry_16_port, A2 => n28, ZN => 
                           sub_126_G15_carry_17_port);
   U532 : XOR2_X1 port map( A => n27, B => sub_126_G15_carry_16_port, Z => 
                           A_neg_14_16_port);
   U533 : AND2_X1 port map( A1 => n18, A2 => n25, ZN => 
                           sub_126_G15_carry_16_port);
   U534 : XOR2_X1 port map( A => n24, B => n17, Z => A_neg_14_15_port);
   n69 <= '0';

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CMP_NBIT32 is

   port( SUM : in std_logic_vector (31 downto 0);  Cout : in std_logic;  A_L_B,
         A_LE_B, A_G_B, A_GE_B, A_E_B, A_NE_B : out std_logic);

end CMP_NBIT32;

architecture SYN_structural of CMP_NBIT32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal A_L_B_port, A_LE_B_port, N29, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      A_E_B_port : std_logic;

begin
   A_L_B <= A_L_B_port;
   A_LE_B <= A_LE_B_port;
   A_E_B <= A_E_B_port;
   A_NE_B <= N29;
   
   U1 : NOR4_X1 port map( A1 => SUM(19), A2 => SUM(18), A3 => SUM(17), A4 => 
                           SUM(16), ZN => n4);
   U2 : NOR4_X1 port map( A1 => SUM(22), A2 => SUM(21), A3 => SUM(20), A4 => 
                           SUM(1), ZN => n5);
   U3 : NOR4_X1 port map( A1 => n12, A2 => SUM(0), A3 => SUM(11), A4 => SUM(10)
                           , ZN => n6);
   U4 : NOR4_X1 port map( A1 => SUM(9), A2 => SUM(8), A3 => SUM(7), A4 => 
                           SUM(6), ZN => n11);
   U5 : OR4_X1 port map( A1 => SUM(13), A2 => SUM(12), A3 => SUM(15), A4 => 
                           SUM(14), ZN => n12);
   U6 : INV_X1 port map( A => A_LE_B_port, ZN => A_G_B);
   U7 : NOR4_X1 port map( A1 => SUM(26), A2 => SUM(25), A3 => SUM(24), A4 => 
                           SUM(23), ZN => n8);
   U8 : NOR4_X1 port map( A1 => SUM(2), A2 => SUM(29), A3 => SUM(28), A4 => 
                           SUM(27), ZN => n9);
   U9 : NAND2_X1 port map( A1 => Cout, A2 => N29, ZN => A_LE_B_port);
   U10 : NAND4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => N29);
   U11 : AND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n7);
   U12 : INV_X1 port map( A => A_L_B_port, ZN => A_GE_B);
   U13 : NOR2_X1 port map( A1 => A_E_B_port, A2 => Cout, ZN => A_L_B_port);
   U14 : INV_X1 port map( A => N29, ZN => A_E_B_port);
   U15 : NOR4_X1 port map( A1 => SUM(30), A2 => SUM(4), A3 => SUM(3), A4 => 
                           SUM(5), ZN => n10);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LOGIC_NBIT32_N_SELECTOR4 is

   port( S : in std_logic_vector (3 downto 0);  A, B : in std_logic_vector (31 
         downto 0);  O : out std_logic_vector (31 downto 0));

end LOGIC_NBIT32_N_SELECTOR4;

architecture SYN_structural of LOGIC_NBIT32_N_SELECTOR4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4_1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_2
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_3
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_4
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_2
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_5
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_6
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_7
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_8
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_3
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_9
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_10
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_11
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_12
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_4
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_13
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_14
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_15
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_16
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_5
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_17
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_18
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_19
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_20
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_6
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_21
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_22
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_23
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_24
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_7
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_25
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_26
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_27
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_28
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_8
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_29
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_30
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_31
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_32
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_9
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_33
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_34
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_35
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_36
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_10
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_37
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_38
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_39
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_40
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_11
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_41
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_42
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_43
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_44
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_12
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_45
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_46
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_47
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_48
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_13
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_49
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_50
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_51
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_52
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_14
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_53
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_54
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_55
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_56
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_15
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_57
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_58
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_59
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_60
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_16
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_61
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_62
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_63
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_64
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_17
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_65
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_66
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_67
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_68
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_18
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_69
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_70
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_71
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_72
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_19
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_73
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_74
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_75
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_76
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_20
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_77
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_78
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_79
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_80
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_21
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_81
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_82
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_83
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_84
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_22
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_85
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_86
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_87
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_88
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_23
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_89
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_90
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_91
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_92
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_24
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_93
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_94
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_95
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_96
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_25
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_97
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_98
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_99
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_100
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_26
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_101
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_102
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_103
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_104
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_27
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_105
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_106
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_107
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_108
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_28
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_109
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_110
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_111
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_112
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_29
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_113
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_114
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_115
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_116
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_30
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_117
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_118
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_119
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_120
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_31
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_121
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_122
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_123
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_124
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND4_0
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_125
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_126
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_127
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component ND3_0
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal An_31_port, An_30_port, An_29_port, An_28_port, An_27_port, 
      An_26_port, An_25_port, An_24_port, An_23_port, An_22_port, An_21_port, 
      An_20_port, An_19_port, An_18_port, An_17_port, An_16_port, An_15_port, 
      An_14_port, An_13_port, An_12_port, An_11_port, An_10_port, An_9_port, 
      An_8_port, An_7_port, An_6_port, An_5_port, An_4_port, An_3_port, 
      An_2_port, An_1_port, An_0_port, Bn_31_port, Bn_30_port, Bn_29_port, 
      Bn_28_port, Bn_27_port, Bn_26_port, Bn_25_port, Bn_24_port, Bn_23_port, 
      Bn_22_port, Bn_21_port, Bn_20_port, Bn_19_port, Bn_18_port, Bn_17_port, 
      Bn_16_port, Bn_15_port, Bn_14_port, Bn_13_port, Bn_12_port, Bn_11_port, 
      Bn_10_port, Bn_9_port, Bn_8_port, Bn_7_port, Bn_6_port, Bn_5_port, 
      Bn_4_port, Bn_3_port, Bn_2_port, Bn_1_port, Bn_0_port, l0_31_port, 
      l0_30_port, l0_29_port, l0_28_port, l0_27_port, l0_26_port, l0_25_port, 
      l0_24_port, l0_23_port, l0_22_port, l0_21_port, l0_20_port, l0_19_port, 
      l0_18_port, l0_17_port, l0_16_port, l0_15_port, l0_14_port, l0_13_port, 
      l0_12_port, l0_11_port, l0_10_port, l0_9_port, l0_8_port, l0_7_port, 
      l0_6_port, l0_5_port, l0_4_port, l0_3_port, l0_2_port, l0_1_port, 
      l0_0_port, l1_31_port, l1_30_port, l1_29_port, l1_28_port, l1_27_port, 
      l1_26_port, l1_25_port, l1_24_port, l1_23_port, l1_22_port, l1_21_port, 
      l1_20_port, l1_19_port, l1_18_port, l1_17_port, l1_16_port, l1_15_port, 
      l1_14_port, l1_13_port, l1_12_port, l1_11_port, l1_10_port, l1_9_port, 
      l1_8_port, l1_7_port, l1_6_port, l1_5_port, l1_4_port, l1_3_port, 
      l1_2_port, l1_1_port, l1_0_port, l2_31_port, l2_30_port, l2_29_port, 
      l2_28_port, l2_27_port, l2_26_port, l2_25_port, l2_24_port, l2_23_port, 
      l2_22_port, l2_21_port, l2_20_port, l2_19_port, l2_18_port, l2_17_port, 
      l2_16_port, l2_15_port, l2_14_port, l2_13_port, l2_12_port, l2_11_port, 
      l2_10_port, l2_9_port, l2_8_port, l2_7_port, l2_6_port, l2_5_port, 
      l2_4_port, l2_3_port, l2_2_port, l2_1_port, l2_0_port, l3_31_port, 
      l3_30_port, l3_29_port, l3_28_port, l3_27_port, l3_26_port, l3_25_port, 
      l3_24_port, l3_23_port, l3_22_port, l3_21_port, l3_20_port, l3_19_port, 
      l3_18_port, l3_17_port, l3_16_port, l3_15_port, l3_14_port, l3_13_port, 
      l3_12_port, l3_11_port, l3_10_port, l3_9_port, l3_8_port, l3_7_port, 
      l3_6_port, l3_5_port, l3_4_port, l3_3_port, l3_2_port, l3_1_port, 
      l3_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16 : std_logic;

begin
   
   A_i_0 : IV_0 port map( A => A(0), Y => An_0_port);
   A_i_1 : IV_63 port map( A => A(1), Y => An_1_port);
   A_i_2 : IV_62 port map( A => A(2), Y => An_2_port);
   A_i_3 : IV_61 port map( A => A(3), Y => An_3_port);
   A_i_4 : IV_60 port map( A => A(4), Y => An_4_port);
   A_i_5 : IV_59 port map( A => A(5), Y => An_5_port);
   A_i_6 : IV_58 port map( A => A(6), Y => An_6_port);
   A_i_7 : IV_57 port map( A => A(7), Y => An_7_port);
   A_i_8 : IV_56 port map( A => A(8), Y => An_8_port);
   A_i_9 : IV_55 port map( A => A(9), Y => An_9_port);
   A_i_10 : IV_54 port map( A => A(10), Y => An_10_port);
   A_i_11 : IV_53 port map( A => A(11), Y => An_11_port);
   A_i_12 : IV_52 port map( A => A(12), Y => An_12_port);
   A_i_13 : IV_51 port map( A => A(13), Y => An_13_port);
   A_i_14 : IV_50 port map( A => A(14), Y => An_14_port);
   A_i_15 : IV_49 port map( A => A(15), Y => An_15_port);
   A_i_16 : IV_48 port map( A => A(16), Y => An_16_port);
   A_i_17 : IV_47 port map( A => A(17), Y => An_17_port);
   A_i_18 : IV_46 port map( A => A(18), Y => An_18_port);
   A_i_19 : IV_45 port map( A => A(19), Y => An_19_port);
   A_i_20 : IV_44 port map( A => A(20), Y => An_20_port);
   A_i_21 : IV_43 port map( A => A(21), Y => An_21_port);
   A_i_22 : IV_42 port map( A => A(22), Y => An_22_port);
   A_i_23 : IV_41 port map( A => A(23), Y => An_23_port);
   A_i_24 : IV_40 port map( A => A(24), Y => An_24_port);
   A_i_25 : IV_39 port map( A => A(25), Y => An_25_port);
   A_i_26 : IV_38 port map( A => A(26), Y => An_26_port);
   A_i_27 : IV_37 port map( A => A(27), Y => An_27_port);
   A_i_28 : IV_36 port map( A => A(28), Y => An_28_port);
   A_i_29 : IV_35 port map( A => A(29), Y => An_29_port);
   A_i_30 : IV_34 port map( A => A(30), Y => An_30_port);
   A_i_31 : IV_33 port map( A => A(31), Y => An_31_port);
   B_i_0 : IV_32 port map( A => B(0), Y => Bn_0_port);
   B_i_1 : IV_31 port map( A => B(1), Y => Bn_1_port);
   B_i_2 : IV_30 port map( A => B(2), Y => Bn_2_port);
   B_i_3 : IV_29 port map( A => B(3), Y => Bn_3_port);
   B_i_4 : IV_28 port map( A => B(4), Y => Bn_4_port);
   B_i_5 : IV_27 port map( A => B(5), Y => Bn_5_port);
   B_i_6 : IV_26 port map( A => B(6), Y => Bn_6_port);
   B_i_7 : IV_25 port map( A => B(7), Y => Bn_7_port);
   B_i_8 : IV_24 port map( A => B(8), Y => Bn_8_port);
   B_i_9 : IV_23 port map( A => B(9), Y => Bn_9_port);
   B_i_10 : IV_22 port map( A => B(10), Y => Bn_10_port);
   B_i_11 : IV_21 port map( A => B(11), Y => Bn_11_port);
   B_i_12 : IV_20 port map( A => B(12), Y => Bn_12_port);
   B_i_13 : IV_19 port map( A => B(13), Y => Bn_13_port);
   B_i_14 : IV_18 port map( A => B(14), Y => Bn_14_port);
   B_i_15 : IV_17 port map( A => B(15), Y => Bn_15_port);
   B_i_16 : IV_16 port map( A => B(16), Y => Bn_16_port);
   B_i_17 : IV_15 port map( A => B(17), Y => Bn_17_port);
   B_i_18 : IV_14 port map( A => B(18), Y => Bn_18_port);
   B_i_19 : IV_13 port map( A => B(19), Y => Bn_19_port);
   B_i_20 : IV_12 port map( A => B(20), Y => Bn_20_port);
   B_i_21 : IV_11 port map( A => B(21), Y => Bn_21_port);
   B_i_22 : IV_10 port map( A => B(22), Y => Bn_22_port);
   B_i_23 : IV_9 port map( A => B(23), Y => Bn_23_port);
   B_i_24 : IV_8 port map( A => B(24), Y => Bn_24_port);
   B_i_25 : IV_7 port map( A => B(25), Y => Bn_25_port);
   B_i_26 : IV_6 port map( A => B(26), Y => Bn_26_port);
   B_i_27 : IV_5 port map( A => B(27), Y => Bn_27_port);
   B_i_28 : IV_4 port map( A => B(28), Y => Bn_28_port);
   B_i_29 : IV_3 port map( A => B(29), Y => Bn_29_port);
   B_i_30 : IV_2 port map( A => B(30), Y => Bn_30_port);
   B_i_31 : IV_1 port map( A => B(31), Y => Bn_31_port);
   U0_0 : ND3_0 port map( A => n3, B => An_0_port, C => Bn_0_port, Y => 
                           l0_0_port);
   U1_0 : ND3_127 port map( A => n5, B => An_0_port, C => B(0), Y => l1_0_port)
                           ;
   U2_0 : ND3_126 port map( A => n9, B => A(0), C => Bn_0_port, Y => l2_0_port)
                           ;
   U3_0 : ND3_125 port map( A => n13, B => A(0), C => B(0), Y => l3_0_port);
   U4_0 : ND4_0 port map( A => l0_0_port, B => l1_0_port, C => l2_0_port, D => 
                           l3_0_port, Y => O(0));
   U0_1 : ND3_124 port map( A => n1, B => An_1_port, C => Bn_1_port, Y => 
                           l0_1_port);
   U1_1 : ND3_123 port map( A => n5, B => An_1_port, C => B(1), Y => l1_1_port)
                           ;
   U2_1 : ND3_122 port map( A => n9, B => A(1), C => Bn_1_port, Y => l2_1_port)
                           ;
   U3_1 : ND3_121 port map( A => n13, B => A(1), C => B(1), Y => l3_1_port);
   U4_1 : ND4_31 port map( A => l0_1_port, B => l1_1_port, C => l2_1_port, D =>
                           l3_1_port, Y => O(1));
   U0_2 : ND3_120 port map( A => n1, B => An_2_port, C => Bn_2_port, Y => 
                           l0_2_port);
   U1_2 : ND3_119 port map( A => n5, B => An_2_port, C => B(2), Y => l1_2_port)
                           ;
   U2_2 : ND3_118 port map( A => n9, B => A(2), C => Bn_2_port, Y => l2_2_port)
                           ;
   U3_2 : ND3_117 port map( A => n13, B => A(2), C => B(2), Y => l3_2_port);
   U4_2 : ND4_30 port map( A => l0_2_port, B => l1_2_port, C => l2_2_port, D =>
                           l3_2_port, Y => O(2));
   U0_3 : ND3_116 port map( A => n1, B => An_3_port, C => Bn_3_port, Y => 
                           l0_3_port);
   U1_3 : ND3_115 port map( A => n5, B => An_3_port, C => B(3), Y => l1_3_port)
                           ;
   U2_3 : ND3_114 port map( A => n9, B => A(3), C => Bn_3_port, Y => l2_3_port)
                           ;
   U3_3 : ND3_113 port map( A => n13, B => A(3), C => B(3), Y => l3_3_port);
   U4_3 : ND4_29 port map( A => l0_3_port, B => l1_3_port, C => l2_3_port, D =>
                           l3_3_port, Y => O(3));
   U0_4 : ND3_112 port map( A => n1, B => An_4_port, C => Bn_4_port, Y => 
                           l0_4_port);
   U1_4 : ND3_111 port map( A => n5, B => An_4_port, C => B(4), Y => l1_4_port)
                           ;
   U2_4 : ND3_110 port map( A => n9, B => A(4), C => Bn_4_port, Y => l2_4_port)
                           ;
   U3_4 : ND3_109 port map( A => n13, B => A(4), C => B(4), Y => l3_4_port);
   U4_4 : ND4_28 port map( A => l0_4_port, B => l1_4_port, C => l2_4_port, D =>
                           l3_4_port, Y => O(4));
   U0_5 : ND3_108 port map( A => n1, B => An_5_port, C => Bn_5_port, Y => 
                           l0_5_port);
   U1_5 : ND3_107 port map( A => n5, B => An_5_port, C => B(5), Y => l1_5_port)
                           ;
   U2_5 : ND3_106 port map( A => n9, B => A(5), C => Bn_5_port, Y => l2_5_port)
                           ;
   U3_5 : ND3_105 port map( A => n13, B => A(5), C => B(5), Y => l3_5_port);
   U4_5 : ND4_27 port map( A => l0_5_port, B => l1_5_port, C => l2_5_port, D =>
                           l3_5_port, Y => O(5));
   U0_6 : ND3_104 port map( A => n1, B => An_6_port, C => Bn_6_port, Y => 
                           l0_6_port);
   U1_6 : ND3_103 port map( A => n5, B => An_6_port, C => B(6), Y => l1_6_port)
                           ;
   U2_6 : ND3_102 port map( A => n9, B => A(6), C => Bn_6_port, Y => l2_6_port)
                           ;
   U3_6 : ND3_101 port map( A => n13, B => A(6), C => B(6), Y => l3_6_port);
   U4_6 : ND4_26 port map( A => l0_6_port, B => l1_6_port, C => l2_6_port, D =>
                           l3_6_port, Y => O(6));
   U0_7 : ND3_100 port map( A => n1, B => An_7_port, C => Bn_7_port, Y => 
                           l0_7_port);
   U1_7 : ND3_99 port map( A => n5, B => An_7_port, C => B(7), Y => l1_7_port);
   U2_7 : ND3_98 port map( A => n9, B => A(7), C => Bn_7_port, Y => l2_7_port);
   U3_7 : ND3_97 port map( A => n13, B => A(7), C => B(7), Y => l3_7_port);
   U4_7 : ND4_25 port map( A => l0_7_port, B => l1_7_port, C => l2_7_port, D =>
                           l3_7_port, Y => O(7));
   U0_8 : ND3_96 port map( A => n1, B => An_8_port, C => Bn_8_port, Y => 
                           l0_8_port);
   U1_8 : ND3_95 port map( A => n5, B => An_8_port, C => B(8), Y => l1_8_port);
   U2_8 : ND3_94 port map( A => n9, B => A(8), C => Bn_8_port, Y => l2_8_port);
   U3_8 : ND3_93 port map( A => n13, B => A(8), C => B(8), Y => l3_8_port);
   U4_8 : ND4_24 port map( A => l0_8_port, B => l1_8_port, C => l2_8_port, D =>
                           l3_8_port, Y => O(8));
   U0_9 : ND3_92 port map( A => n1, B => An_9_port, C => Bn_9_port, Y => 
                           l0_9_port);
   U1_9 : ND3_91 port map( A => n5, B => An_9_port, C => B(9), Y => l1_9_port);
   U2_9 : ND3_90 port map( A => n9, B => A(9), C => Bn_9_port, Y => l2_9_port);
   U3_9 : ND3_89 port map( A => n13, B => A(9), C => B(9), Y => l3_9_port);
   U4_9 : ND4_23 port map( A => l0_9_port, B => l1_9_port, C => l2_9_port, D =>
                           l3_9_port, Y => O(9));
   U0_10 : ND3_88 port map( A => n1, B => An_10_port, C => Bn_10_port, Y => 
                           l0_10_port);
   U1_10 : ND3_87 port map( A => n5, B => An_10_port, C => B(10), Y => 
                           l1_10_port);
   U2_10 : ND3_86 port map( A => n9, B => A(10), C => Bn_10_port, Y => 
                           l2_10_port);
   U3_10 : ND3_85 port map( A => n13, B => A(10), C => B(10), Y => l3_10_port);
   U4_10 : ND4_22 port map( A => l0_10_port, B => l1_10_port, C => l2_10_port, 
                           D => l3_10_port, Y => O(10));
   U0_11 : ND3_84 port map( A => n1, B => An_11_port, C => Bn_11_port, Y => 
                           l0_11_port);
   U1_11 : ND3_83 port map( A => n6, B => An_11_port, C => B(11), Y => 
                           l1_11_port);
   U2_11 : ND3_82 port map( A => n10, B => A(11), C => Bn_11_port, Y => 
                           l2_11_port);
   U3_11 : ND3_81 port map( A => n14, B => A(11), C => B(11), Y => l3_11_port);
   U4_11 : ND4_21 port map( A => l0_11_port, B => l1_11_port, C => l2_11_port, 
                           D => l3_11_port, Y => O(11));
   U0_12 : ND3_80 port map( A => n2, B => An_12_port, C => Bn_12_port, Y => 
                           l0_12_port);
   U1_12 : ND3_79 port map( A => n6, B => An_12_port, C => B(12), Y => 
                           l1_12_port);
   U2_12 : ND3_78 port map( A => n10, B => A(12), C => Bn_12_port, Y => 
                           l2_12_port);
   U3_12 : ND3_77 port map( A => n14, B => A(12), C => B(12), Y => l3_12_port);
   U4_12 : ND4_20 port map( A => l0_12_port, B => l1_12_port, C => l2_12_port, 
                           D => l3_12_port, Y => O(12));
   U0_13 : ND3_76 port map( A => n2, B => An_13_port, C => Bn_13_port, Y => 
                           l0_13_port);
   U1_13 : ND3_75 port map( A => n6, B => An_13_port, C => B(13), Y => 
                           l1_13_port);
   U2_13 : ND3_74 port map( A => n10, B => A(13), C => Bn_13_port, Y => 
                           l2_13_port);
   U3_13 : ND3_73 port map( A => n14, B => A(13), C => B(13), Y => l3_13_port);
   U4_13 : ND4_19 port map( A => l0_13_port, B => l1_13_port, C => l2_13_port, 
                           D => l3_13_port, Y => O(13));
   U0_14 : ND3_72 port map( A => n2, B => An_14_port, C => Bn_14_port, Y => 
                           l0_14_port);
   U1_14 : ND3_71 port map( A => n6, B => An_14_port, C => B(14), Y => 
                           l1_14_port);
   U2_14 : ND3_70 port map( A => n10, B => A(14), C => Bn_14_port, Y => 
                           l2_14_port);
   U3_14 : ND3_69 port map( A => n14, B => A(14), C => B(14), Y => l3_14_port);
   U4_14 : ND4_18 port map( A => l0_14_port, B => l1_14_port, C => l2_14_port, 
                           D => l3_14_port, Y => O(14));
   U0_15 : ND3_68 port map( A => n2, B => An_15_port, C => Bn_15_port, Y => 
                           l0_15_port);
   U1_15 : ND3_67 port map( A => n6, B => An_15_port, C => B(15), Y => 
                           l1_15_port);
   U2_15 : ND3_66 port map( A => n10, B => A(15), C => Bn_15_port, Y => 
                           l2_15_port);
   U3_15 : ND3_65 port map( A => n14, B => A(15), C => B(15), Y => l3_15_port);
   U4_15 : ND4_17 port map( A => l0_15_port, B => l1_15_port, C => l2_15_port, 
                           D => l3_15_port, Y => O(15));
   U0_16 : ND3_64 port map( A => n2, B => An_16_port, C => Bn_16_port, Y => 
                           l0_16_port);
   U1_16 : ND3_63 port map( A => n6, B => An_16_port, C => B(16), Y => 
                           l1_16_port);
   U2_16 : ND3_62 port map( A => n10, B => A(16), C => Bn_16_port, Y => 
                           l2_16_port);
   U3_16 : ND3_61 port map( A => n14, B => A(16), C => B(16), Y => l3_16_port);
   U4_16 : ND4_16 port map( A => l0_16_port, B => l1_16_port, C => l2_16_port, 
                           D => l3_16_port, Y => O(16));
   U0_17 : ND3_60 port map( A => n2, B => An_17_port, C => Bn_17_port, Y => 
                           l0_17_port);
   U1_17 : ND3_59 port map( A => n6, B => An_17_port, C => B(17), Y => 
                           l1_17_port);
   U2_17 : ND3_58 port map( A => n10, B => A(17), C => Bn_17_port, Y => 
                           l2_17_port);
   U3_17 : ND3_57 port map( A => n14, B => A(17), C => B(17), Y => l3_17_port);
   U4_17 : ND4_15 port map( A => l0_17_port, B => l1_17_port, C => l2_17_port, 
                           D => l3_17_port, Y => O(17));
   U0_18 : ND3_56 port map( A => n2, B => An_18_port, C => Bn_18_port, Y => 
                           l0_18_port);
   U1_18 : ND3_55 port map( A => n6, B => An_18_port, C => B(18), Y => 
                           l1_18_port);
   U2_18 : ND3_54 port map( A => n10, B => A(18), C => Bn_18_port, Y => 
                           l2_18_port);
   U3_18 : ND3_53 port map( A => n14, B => A(18), C => B(18), Y => l3_18_port);
   U4_18 : ND4_14 port map( A => l0_18_port, B => l1_18_port, C => l2_18_port, 
                           D => l3_18_port, Y => O(18));
   U0_19 : ND3_52 port map( A => n2, B => An_19_port, C => Bn_19_port, Y => 
                           l0_19_port);
   U1_19 : ND3_51 port map( A => n6, B => An_19_port, C => B(19), Y => 
                           l1_19_port);
   U2_19 : ND3_50 port map( A => n10, B => A(19), C => Bn_19_port, Y => 
                           l2_19_port);
   U3_19 : ND3_49 port map( A => n14, B => A(19), C => B(19), Y => l3_19_port);
   U4_19 : ND4_13 port map( A => l0_19_port, B => l1_19_port, C => l2_19_port, 
                           D => l3_19_port, Y => O(19));
   U0_20 : ND3_48 port map( A => n2, B => An_20_port, C => Bn_20_port, Y => 
                           l0_20_port);
   U1_20 : ND3_47 port map( A => n6, B => An_20_port, C => B(20), Y => 
                           l1_20_port);
   U2_20 : ND3_46 port map( A => n10, B => A(20), C => Bn_20_port, Y => 
                           l2_20_port);
   U3_20 : ND3_45 port map( A => n14, B => A(20), C => B(20), Y => l3_20_port);
   U4_20 : ND4_12 port map( A => l0_20_port, B => l1_20_port, C => l2_20_port, 
                           D => l3_20_port, Y => O(20));
   U0_21 : ND3_44 port map( A => n2, B => An_21_port, C => Bn_21_port, Y => 
                           l0_21_port);
   U1_21 : ND3_43 port map( A => n6, B => An_21_port, C => B(21), Y => 
                           l1_21_port);
   U2_21 : ND3_42 port map( A => n10, B => A(21), C => Bn_21_port, Y => 
                           l2_21_port);
   U3_21 : ND3_41 port map( A => n14, B => A(21), C => B(21), Y => l3_21_port);
   U4_21 : ND4_11 port map( A => l0_21_port, B => l1_21_port, C => l2_21_port, 
                           D => l3_21_port, Y => O(21));
   U0_22 : ND3_40 port map( A => n2, B => An_22_port, C => Bn_22_port, Y => 
                           l0_22_port);
   U1_22 : ND3_39 port map( A => n7, B => An_22_port, C => B(22), Y => 
                           l1_22_port);
   U2_22 : ND3_38 port map( A => n11, B => A(22), C => Bn_22_port, Y => 
                           l2_22_port);
   U3_22 : ND3_37 port map( A => n15, B => A(22), C => B(22), Y => l3_22_port);
   U4_22 : ND4_10 port map( A => l0_22_port, B => l1_22_port, C => l2_22_port, 
                           D => l3_22_port, Y => O(22));
   U0_23 : ND3_36 port map( A => n3, B => An_23_port, C => Bn_23_port, Y => 
                           l0_23_port);
   U1_23 : ND3_35 port map( A => n7, B => An_23_port, C => B(23), Y => 
                           l1_23_port);
   U2_23 : ND3_34 port map( A => n11, B => A(23), C => Bn_23_port, Y => 
                           l2_23_port);
   U3_23 : ND3_33 port map( A => n15, B => A(23), C => B(23), Y => l3_23_port);
   U4_23 : ND4_9 port map( A => l0_23_port, B => l1_23_port, C => l2_23_port, D
                           => l3_23_port, Y => O(23));
   U0_24 : ND3_32 port map( A => n3, B => An_24_port, C => Bn_24_port, Y => 
                           l0_24_port);
   U1_24 : ND3_31 port map( A => n7, B => An_24_port, C => B(24), Y => 
                           l1_24_port);
   U2_24 : ND3_30 port map( A => n11, B => A(24), C => Bn_24_port, Y => 
                           l2_24_port);
   U3_24 : ND3_29 port map( A => n15, B => A(24), C => B(24), Y => l3_24_port);
   U4_24 : ND4_8 port map( A => l0_24_port, B => l1_24_port, C => l2_24_port, D
                           => l3_24_port, Y => O(24));
   U0_25 : ND3_28 port map( A => n3, B => An_25_port, C => Bn_25_port, Y => 
                           l0_25_port);
   U1_25 : ND3_27 port map( A => n7, B => An_25_port, C => B(25), Y => 
                           l1_25_port);
   U2_25 : ND3_26 port map( A => n11, B => A(25), C => Bn_25_port, Y => 
                           l2_25_port);
   U3_25 : ND3_25 port map( A => n15, B => A(25), C => B(25), Y => l3_25_port);
   U4_25 : ND4_7 port map( A => l0_25_port, B => l1_25_port, C => l2_25_port, D
                           => l3_25_port, Y => O(25));
   U0_26 : ND3_24 port map( A => n3, B => An_26_port, C => Bn_26_port, Y => 
                           l0_26_port);
   U1_26 : ND3_23 port map( A => n7, B => An_26_port, C => B(26), Y => 
                           l1_26_port);
   U2_26 : ND3_22 port map( A => n11, B => A(26), C => Bn_26_port, Y => 
                           l2_26_port);
   U3_26 : ND3_21 port map( A => n15, B => A(26), C => B(26), Y => l3_26_port);
   U4_26 : ND4_6 port map( A => l0_26_port, B => l1_26_port, C => l2_26_port, D
                           => l3_26_port, Y => O(26));
   U0_27 : ND3_20 port map( A => n3, B => An_27_port, C => Bn_27_port, Y => 
                           l0_27_port);
   U1_27 : ND3_19 port map( A => n7, B => An_27_port, C => B(27), Y => 
                           l1_27_port);
   U2_27 : ND3_18 port map( A => n11, B => A(27), C => Bn_27_port, Y => 
                           l2_27_port);
   U3_27 : ND3_17 port map( A => n15, B => A(27), C => B(27), Y => l3_27_port);
   U4_27 : ND4_5 port map( A => l0_27_port, B => l1_27_port, C => l2_27_port, D
                           => l3_27_port, Y => O(27));
   U0_28 : ND3_16 port map( A => n3, B => An_28_port, C => Bn_28_port, Y => 
                           l0_28_port);
   U1_28 : ND3_15 port map( A => n7, B => An_28_port, C => B(28), Y => 
                           l1_28_port);
   U2_28 : ND3_14 port map( A => n11, B => A(28), C => Bn_28_port, Y => 
                           l2_28_port);
   U3_28 : ND3_13 port map( A => n15, B => A(28), C => B(28), Y => l3_28_port);
   U4_28 : ND4_4 port map( A => l0_28_port, B => l1_28_port, C => l2_28_port, D
                           => l3_28_port, Y => O(28));
   U0_29 : ND3_12 port map( A => n3, B => An_29_port, C => Bn_29_port, Y => 
                           l0_29_port);
   U1_29 : ND3_11 port map( A => n7, B => An_29_port, C => B(29), Y => 
                           l1_29_port);
   U2_29 : ND3_10 port map( A => n11, B => A(29), C => Bn_29_port, Y => 
                           l2_29_port);
   U3_29 : ND3_9 port map( A => n15, B => A(29), C => B(29), Y => l3_29_port);
   U4_29 : ND4_3 port map( A => l0_29_port, B => l1_29_port, C => l2_29_port, D
                           => l3_29_port, Y => O(29));
   U0_30 : ND3_8 port map( A => n3, B => An_30_port, C => Bn_30_port, Y => 
                           l0_30_port);
   U1_30 : ND3_7 port map( A => n7, B => An_30_port, C => B(30), Y => 
                           l1_30_port);
   U2_30 : ND3_6 port map( A => n11, B => A(30), C => Bn_30_port, Y => 
                           l2_30_port);
   U3_30 : ND3_5 port map( A => n15, B => A(30), C => B(30), Y => l3_30_port);
   U4_30 : ND4_2 port map( A => l0_30_port, B => l1_30_port, C => l2_30_port, D
                           => l3_30_port, Y => O(30));
   U0_31 : ND3_4 port map( A => n3, B => An_31_port, C => Bn_31_port, Y => 
                           l0_31_port);
   U1_31 : ND3_3 port map( A => n7, B => An_31_port, C => B(31), Y => 
                           l1_31_port);
   U2_31 : ND3_2 port map( A => n11, B => A(31), C => Bn_31_port, Y => 
                           l2_31_port);
   U3_31 : ND3_1 port map( A => n15, B => A(31), C => B(31), Y => l3_31_port);
   U4_31 : ND4_1 port map( A => l0_31_port, B => l1_31_port, C => l2_31_port, D
                           => l3_31_port, Y => O(31));
   U1 : BUF_X1 port map( A => S(0), Z => n4);
   U2 : BUF_X1 port map( A => S(1), Z => n8);
   U3 : BUF_X1 port map( A => S(2), Z => n12);
   U4 : BUF_X1 port map( A => S(3), Z => n16);
   U5 : BUF_X1 port map( A => n8, Z => n5);
   U6 : BUF_X1 port map( A => n12, Z => n9);
   U7 : BUF_X1 port map( A => n16, Z => n13);
   U8 : BUF_X1 port map( A => n4, Z => n1);
   U9 : BUF_X1 port map( A => n8, Z => n6);
   U10 : BUF_X1 port map( A => n12, Z => n10);
   U11 : BUF_X1 port map( A => n16, Z => n14);
   U12 : BUF_X1 port map( A => n4, Z => n2);
   U13 : BUF_X1 port map( A => n4, Z => n3);
   U14 : BUF_X1 port map( A => n8, Z => n7);
   U15 : BUF_X1 port map( A => n12, Z => n11);
   U16 : BUF_X1 port map( A => n16, Z => n15);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SHIFTER is

   port( data_in : in std_logic_vector (31 downto 0);  R : in std_logic_vector 
         (4 downto 0);  conf : in std_logic_vector (1 downto 0);  data_out : 
         out std_logic_vector (31 downto 0));

end SHIFTER;

architecture SYN_Behavioral of SHIFTER is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal mask_0_39_port, mask_0_38_port, mask_0_37_port, mask_0_36_port, 
      mask_0_35_port, mask_0_34_port, mask_0_33_port, mask_0_32_port, 
      mask_0_31_port, mask_0_30_port, mask_0_29_port, mask_0_28_port, 
      mask_0_27_port, mask_0_26_port, mask_0_25_port, mask_0_24_port, 
      mask_0_23_port, mask_0_22_port, mask_0_21_port, mask_0_20_port, 
      mask_0_19_port, mask_0_18_port, mask_0_17_port, mask_0_16_port, 
      mask_0_15_port, mask_0_14_port, mask_0_13_port, mask_0_12_port, 
      mask_0_11_port, mask_0_10_port, mask_0_9_port, mask_0_8_port, 
      mask_0_7_port, mask_0_6_port, mask_0_5_port, mask_0_4_port, mask_0_3_port
      , mask_0_2_port, mask_0_1_port, mask_0_0_port, mask_1_39_port, 
      mask_1_38_port, mask_1_37_port, mask_1_36_port, mask_1_35_port, 
      mask_1_34_port, mask_1_33_port, mask_1_32_port, mask_1_31_port, 
      mask_1_30_port, mask_1_29_port, mask_1_28_port, mask_1_27_port, 
      mask_1_26_port, mask_1_25_port, mask_1_24_port, mask_1_23_port, 
      mask_1_22_port, mask_1_21_port, mask_1_20_port, mask_1_19_port, 
      mask_1_18_port, mask_1_17_port, mask_1_16_port, mask_1_15_port, 
      mask_1_14_port, mask_1_13_port, mask_1_12_port, mask_1_11_port, 
      mask_1_10_port, mask_1_9_port, mask_1_8_port, mask_1_7_port, 
      mask_1_6_port, mask_1_5_port, mask_1_4_port, mask_1_3_port, mask_1_2_port
      , mask_1_1_port, mask_1_0_port, mask_2_39_port, mask_2_38_port, 
      mask_2_37_port, mask_2_36_port, mask_2_35_port, mask_2_34_port, 
      mask_2_33_port, mask_2_32_port, mask_2_31_port, mask_2_30_port, 
      mask_2_29_port, mask_2_28_port, mask_2_27_port, mask_2_26_port, 
      mask_2_25_port, mask_2_24_port, mask_2_23_port, mask_2_22_port, 
      mask_2_21_port, mask_2_20_port, mask_2_19_port, mask_2_18_port, 
      mask_2_17_port, mask_2_16_port, mask_2_15_port, mask_2_14_port, 
      mask_2_13_port, mask_2_12_port, mask_2_11_port, mask_2_10_port, 
      mask_2_9_port, mask_2_8_port, mask_2_7_port, mask_2_6_port, mask_2_5_port
      , mask_2_4_port, mask_2_3_port, mask_2_2_port, mask_2_1_port, 
      mask_2_0_port, mask_3_39_port, mask_3_38_port, mask_3_37_port, 
      mask_3_36_port, mask_3_35_port, mask_3_34_port, mask_3_33_port, 
      mask_3_32_port, mask_3_31_port, mask_3_30_port, mask_3_29_port, 
      mask_3_28_port, mask_3_27_port, mask_3_26_port, mask_3_25_port, 
      mask_3_24_port, mask_3_23_port, mask_3_22_port, mask_3_21_port, 
      mask_3_20_port, mask_3_19_port, mask_3_18_port, mask_3_17_port, 
      mask_3_16_port, mask_3_15_port, mask_3_14_port, mask_3_13_port, 
      mask_3_12_port, mask_3_11_port, mask_3_10_port, mask_3_9_port, 
      mask_3_8_port, mask_3_7_port, mask_3_6_port, mask_3_5_port, mask_3_4_port
      , mask_3_3_port, mask_3_2_port, mask_3_1_port, mask_3_0_port, N28, N35, 
      N37, N38, N39, N40, N41, N42, N43, N45, N46, N47, N48, N49, N50, N51, N53
      , N54, N55, N56, N57, N58, N59, N60, N68, N69, N70, N71, N72, N73, N74, 
      N75, N76, N77, N78, N79, N80, N81, N82, N83, N85, N86, N87, N88, N89, N90
      , N91, N92, N93, N94, N95, N96, N97, N98, N99, N108, N109, N110, N111, 
      N112, N113, N114, N115, N116, out_mask_39_port, out_mask_37_port, 
      out_mask_36_port, out_mask_35_port, out_mask_34_port, out_mask_33_port, 
      out_mask_32_port, out_mask_31_port, out_mask_30_port, out_mask_29_port, 
      out_mask_28_port, out_mask_27_port, out_mask_26_port, out_mask_25_port, 
      out_mask_24_port, out_mask_23_port, out_mask_22_port, out_mask_21_port, 
      out_mask_20_port, out_mask_19_port, out_mask_18_port, out_mask_17_port, 
      out_mask_16_port, out_mask_15_port, out_mask_14_port, out_mask_13_port, 
      out_mask_12_port, out_mask_11_port, out_mask_10_port, out_mask_9_port, 
      out_mask_8_port, out_mask_7_port, out_mask_6_port, out_mask_5_port, 
      out_mask_4_port, out_mask_3_port, out_mask_2_port, out_mask_0_port, N158,
      N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
      N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, 
      N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, 
      N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, 
      N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, 
      N219, N220, N221, n86_port, n87_port, n90_port, n91_port, n92_port, 
      n93_port, n94_port, n95_port, n96_port, n97_port, n98_port, n99_port, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108_port, n109_port, 
      n110_port, n111_port, n112_port, n113_port, n114_port, n115_port, 
      n116_port, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158_port, n159_port, n160_port
      , n161_port, n162_port, n163_port, n164_port, n165_port, n166_port, 
      n167_port, n168_port, n169_port, n170_port, n172_port, n173_port, 
      n174_port, n175_port, n176_port, n177_port, n178_port, n179_port, 
      n180_port, n181_port, n182_port, n183_port, n184_port, n185_port, 
      n186_port, n187_port, n188_port, n189_port, n190_port, n191_port, 
      n192_port, n193_port, n194_port, n195_port, n196_port, n197_port, 
      n198_port, n199_port, n200_port, n201_port, n202_port, n203_port, 
      n204_port, n205_port, n206_port, n207_port, n208_port, n209_port, 
      n210_port, n211_port, n212_port, n213_port, n214_port, n215_port, 
      n216_port, n217_port, n219_port, n220_port, n221_port, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n1, n2,
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28_port, n29, n30, n31, n32
      , n33, n34, n35_port, n36, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44, n45_port, n46_port, n47_port, n48_port
      , n49_port, n50_port, n51_port, n52, n53_port, n54_port, n55_port, 
      n56_port, n57_port, n58_port, n59_port, n60_port, n61, n62, n63, n64, n65
      , n66, n67, n68_port, n69_port, n70_port, n71_port, n72_port, n73_port, 
      n74_port, n75_port, n76_port, n77_port, n78_port, n79_port, n80_port, 
      n81_port, n82_port, n83_port, n84, n85_port, n88_port, n89_port, 
      n171_port, n218_port, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n532, n533, n534 : std_logic;

begin
   
   mask_reg_0_39_inst : DLH_X1 port map( G => n443, D => n453, Q => 
                           mask_0_39_port);
   mask_reg_0_38_inst : DLH_X1 port map( G => n443, D => n454, Q => 
                           mask_0_38_port);
   mask_reg_0_37_inst : DLH_X1 port map( G => n443, D => n455, Q => 
                           mask_0_37_port);
   mask_reg_0_36_inst : DLH_X1 port map( G => n443, D => n456, Q => 
                           mask_0_36_port);
   mask_reg_0_35_inst : DLH_X1 port map( G => n443, D => n457, Q => 
                           mask_0_35_port);
   mask_reg_0_34_inst : DLH_X1 port map( G => n443, D => n458, Q => 
                           mask_0_34_port);
   mask_reg_0_33_inst : DLH_X1 port map( G => n443, D => n459, Q => 
                           mask_0_33_port);
   mask_reg_0_32_inst : DLH_X1 port map( G => n443, D => n460, Q => 
                           mask_0_32_port);
   mask_reg_0_31_inst : DLH_X1 port map( G => n443, D => N116, Q => 
                           mask_0_31_port);
   mask_reg_0_30_inst : DLH_X1 port map( G => n443, D => N115, Q => 
                           mask_0_30_port);
   mask_reg_0_29_inst : DLH_X1 port map( G => n442, D => N114, Q => 
                           mask_0_29_port);
   mask_reg_0_28_inst : DLH_X1 port map( G => n442, D => N113, Q => 
                           mask_0_28_port);
   mask_reg_0_27_inst : DLH_X1 port map( G => n442, D => N112, Q => 
                           mask_0_27_port);
   mask_reg_0_26_inst : DLH_X1 port map( G => n442, D => N111, Q => 
                           mask_0_26_port);
   mask_reg_0_25_inst : DLH_X1 port map( G => n442, D => N110, Q => 
                           mask_0_25_port);
   mask_reg_0_24_inst : DLH_X1 port map( G => n442, D => N109, Q => 
                           mask_0_24_port);
   mask_reg_0_23_inst : DLH_X1 port map( G => n442, D => N108, Q => 
                           mask_0_23_port);
   mask_reg_0_22_inst : DLH_X1 port map( G => n442, D => n470, Q => 
                           mask_0_22_port);
   mask_reg_0_21_inst : DLH_X1 port map( G => n442, D => n472, Q => 
                           mask_0_21_port);
   mask_reg_0_20_inst : DLH_X1 port map( G => n442, D => n474, Q => 
                           mask_0_20_port);
   mask_reg_0_19_inst : DLH_X1 port map( G => n441, D => n476, Q => 
                           mask_0_19_port);
   mask_reg_0_18_inst : DLH_X1 port map( G => n441, D => n478, Q => 
                           mask_0_18_port);
   mask_reg_0_17_inst : DLH_X1 port map( G => n441, D => n480, Q => 
                           mask_0_17_port);
   mask_reg_0_16_inst : DLH_X1 port map( G => n441, D => n482, Q => 
                           mask_0_16_port);
   mask_reg_0_15_inst : DLH_X1 port map( G => n441, D => n484, Q => 
                           mask_0_15_port);
   mask_reg_0_14_inst : DLH_X1 port map( G => n441, D => N99, Q => 
                           mask_0_14_port);
   mask_reg_0_13_inst : DLH_X1 port map( G => n441, D => N98, Q => 
                           mask_0_13_port);
   mask_reg_0_12_inst : DLH_X1 port map( G => n441, D => N97, Q => 
                           mask_0_12_port);
   mask_reg_0_11_inst : DLH_X1 port map( G => n441, D => N96, Q => 
                           mask_0_11_port);
   mask_reg_0_10_inst : DLH_X1 port map( G => n441, D => N95, Q => 
                           mask_0_10_port);
   mask_reg_0_9_inst : DLH_X1 port map( G => n440, D => N94, Q => mask_0_9_port
                           );
   mask_reg_0_8_inst : DLH_X1 port map( G => n440, D => N93, Q => mask_0_8_port
                           );
   mask_reg_0_7_inst : DLH_X1 port map( G => n440, D => N92, Q => mask_0_7_port
                           );
   mask_reg_0_6_inst : DLH_X1 port map( G => n440, D => N91, Q => mask_0_6_port
                           );
   mask_reg_0_5_inst : DLH_X1 port map( G => n440, D => N90, Q => mask_0_5_port
                           );
   mask_reg_0_4_inst : DLH_X1 port map( G => n440, D => N89, Q => mask_0_4_port
                           );
   mask_reg_0_3_inst : DLH_X1 port map( G => n440, D => N88, Q => mask_0_3_port
                           );
   mask_reg_0_2_inst : DLH_X1 port map( G => n440, D => N87, Q => mask_0_2_port
                           );
   mask_reg_0_1_inst : DLH_X1 port map( G => n440, D => N86, Q => mask_0_1_port
                           );
   mask_reg_0_0_inst : DLH_X1 port map( G => n440, D => N85, Q => mask_0_0_port
                           );
   mask_reg_1_39_inst : DLH_X1 port map( G => n439, D => n461, Q => 
                           mask_1_39_port);
   mask_reg_1_38_inst : DLH_X1 port map( G => n439, D => N83, Q => 
                           mask_1_38_port);
   mask_reg_1_37_inst : DLH_X1 port map( G => n439, D => N82, Q => 
                           mask_1_37_port);
   mask_reg_1_36_inst : DLH_X1 port map( G => n439, D => N81, Q => 
                           mask_1_36_port);
   mask_reg_1_35_inst : DLH_X1 port map( G => n439, D => N80, Q => 
                           mask_1_35_port);
   mask_reg_1_34_inst : DLH_X1 port map( G => n439, D => N79, Q => 
                           mask_1_34_port);
   mask_reg_1_33_inst : DLH_X1 port map( G => n439, D => N78, Q => 
                           mask_1_33_port);
   mask_reg_1_32_inst : DLH_X1 port map( G => n439, D => N77, Q => 
                           mask_1_32_port);
   mask_reg_1_31_inst : DLH_X1 port map( G => n439, D => N60, Q => 
                           mask_1_31_port);
   mask_reg_1_30_inst : DLH_X1 port map( G => n439, D => N59, Q => 
                           mask_1_30_port);
   mask_reg_1_29_inst : DLH_X1 port map( G => n438, D => N58, Q => 
                           mask_1_29_port);
   mask_reg_1_28_inst : DLH_X1 port map( G => n438, D => N57, Q => 
                           mask_1_28_port);
   mask_reg_1_27_inst : DLH_X1 port map( G => n438, D => N56, Q => 
                           mask_1_27_port);
   mask_reg_1_26_inst : DLH_X1 port map( G => n438, D => N55, Q => 
                           mask_1_26_port);
   mask_reg_1_25_inst : DLH_X1 port map( G => n438, D => N54, Q => 
                           mask_1_25_port);
   mask_reg_1_24_inst : DLH_X1 port map( G => n438, D => N53, Q => 
                           mask_1_24_port);
   mask_reg_1_23_inst : DLH_X1 port map( G => n438, D => N76, Q => 
                           mask_1_23_port);
   mask_reg_1_22_inst : DLH_X1 port map( G => n438, D => N75, Q => 
                           mask_1_22_port);
   mask_reg_1_21_inst : DLH_X1 port map( G => n438, D => N74, Q => 
                           mask_1_21_port);
   mask_reg_1_20_inst : DLH_X1 port map( G => n438, D => N73, Q => 
                           mask_1_20_port);
   mask_reg_1_19_inst : DLH_X1 port map( G => n437, D => N72, Q => 
                           mask_1_19_port);
   mask_reg_1_18_inst : DLH_X1 port map( G => n437, D => N71, Q => 
                           mask_1_18_port);
   mask_reg_1_17_inst : DLH_X1 port map( G => n437, D => N70, Q => 
                           mask_1_17_port);
   mask_reg_1_16_inst : DLH_X1 port map( G => n437, D => N69, Q => 
                           mask_1_16_port);
   mask_reg_1_15_inst : DLH_X1 port map( G => n437, D => n469, Q => 
                           mask_1_15_port);
   mask_reg_1_14_inst : DLH_X1 port map( G => n437, D => N51, Q => 
                           mask_1_14_port);
   mask_reg_1_13_inst : DLH_X1 port map( G => n437, D => N50, Q => 
                           mask_1_13_port);
   mask_reg_1_12_inst : DLH_X1 port map( G => n437, D => N49, Q => 
                           mask_1_12_port);
   mask_reg_1_11_inst : DLH_X1 port map( G => n437, D => N48, Q => 
                           mask_1_11_port);
   mask_reg_1_10_inst : DLH_X1 port map( G => n437, D => N47, Q => 
                           mask_1_10_port);
   mask_reg_1_9_inst : DLH_X1 port map( G => n436, D => N46, Q => mask_1_9_port
                           );
   mask_reg_1_8_inst : DLH_X1 port map( G => n436, D => N45, Q => mask_1_8_port
                           );
   mask_reg_1_7_inst : DLH_X1 port map( G => n436, D => N68, Q => mask_1_7_port
                           );
   mask_reg_1_6_inst : DLH_X1 port map( G => n436, D => n487, Q => 
                           mask_1_6_port);
   mask_reg_1_5_inst : DLH_X1 port map( G => n436, D => n489, Q => 
                           mask_1_5_port);
   mask_reg_1_4_inst : DLH_X1 port map( G => n436, D => n491, Q => 
                           mask_1_4_port);
   mask_reg_1_3_inst : DLH_X1 port map( G => n436, D => n493, Q => 
                           mask_1_3_port);
   mask_reg_1_2_inst : DLH_X1 port map( G => n436, D => n495, Q => 
                           mask_1_2_port);
   mask_reg_1_1_inst : DLH_X1 port map( G => n436, D => n497, Q => 
                           mask_1_1_port);
   mask_reg_1_0_inst : DLH_X1 port map( G => n436, D => n499, Q => 
                           mask_1_0_port);
   mask_reg_2_39_inst : DLH_X1 port map( G => n435, D => N60, Q => 
                           mask_2_39_port);
   mask_reg_2_38_inst : DLH_X1 port map( G => n435, D => N59, Q => 
                           mask_2_38_port);
   mask_reg_2_37_inst : DLH_X1 port map( G => n435, D => N58, Q => 
                           mask_2_37_port);
   mask_reg_2_36_inst : DLH_X1 port map( G => n435, D => N57, Q => 
                           mask_2_36_port);
   mask_reg_2_35_inst : DLH_X1 port map( G => n435, D => N56, Q => 
                           mask_2_35_port);
   mask_reg_2_34_inst : DLH_X1 port map( G => n435, D => N55, Q => 
                           mask_2_34_port);
   mask_reg_2_33_inst : DLH_X1 port map( G => n435, D => N54, Q => 
                           mask_2_33_port);
   mask_reg_2_32_inst : DLH_X1 port map( G => n435, D => N53, Q => 
                           mask_2_32_port);
   mask_reg_2_31_inst : DLH_X1 port map( G => n435, D => n452, Q => 
                           mask_2_31_port);
   mask_reg_2_30_inst : DLH_X1 port map( G => n435, D => N43, Q => 
                           mask_2_30_port);
   mask_reg_2_29_inst : DLH_X1 port map( G => n434, D => N42, Q => 
                           mask_2_29_port);
   mask_reg_2_28_inst : DLH_X1 port map( G => n434, D => N41, Q => 
                           mask_2_28_port);
   mask_reg_2_27_inst : DLH_X1 port map( G => n434, D => N40, Q => 
                           mask_2_27_port);
   mask_reg_2_26_inst : DLH_X1 port map( G => n434, D => N39, Q => 
                           mask_2_26_port);
   mask_reg_2_25_inst : DLH_X1 port map( G => n434, D => N38, Q => 
                           mask_2_25_port);
   mask_reg_2_24_inst : DLH_X1 port map( G => n434, D => N37, Q => 
                           mask_2_24_port);
   mask_reg_2_23_inst : DLH_X1 port map( G => n434, D => n397, Q => 
                           mask_2_23_port);
   mask_reg_2_22_inst : DLH_X1 port map( G => n434, D => n397, Q => 
                           mask_2_22_port);
   mask_reg_2_21_inst : DLH_X1 port map( G => n434, D => n397, Q => 
                           mask_2_21_port);
   mask_reg_2_20_inst : DLH_X1 port map( G => n434, D => n397, Q => 
                           mask_2_20_port);
   mask_reg_2_19_inst : DLH_X1 port map( G => n433, D => n397, Q => 
                           mask_2_19_port);
   mask_reg_2_18_inst : DLH_X1 port map( G => n433, D => n390, Q => 
                           mask_2_18_port);
   mask_reg_2_17_inst : DLH_X1 port map( G => n433, D => n390, Q => 
                           mask_2_17_port);
   mask_reg_2_16_inst : DLH_X1 port map( G => n433, D => n390, Q => 
                           mask_2_16_port);
   mask_reg_2_15_inst : DLH_X1 port map( G => n433, D => N35, Q => 
                           mask_2_15_port);
   mask_reg_2_14_inst : DLH_X1 port map( G => n433, D => n462, Q => 
                           mask_2_14_port);
   mask_reg_2_13_inst : DLH_X1 port map( G => n433, D => n463, Q => 
                           mask_2_13_port);
   mask_reg_2_12_inst : DLH_X1 port map( G => n433, D => n464, Q => 
                           mask_2_12_port);
   mask_reg_2_11_inst : DLH_X1 port map( G => n433, D => n465, Q => 
                           mask_2_11_port);
   mask_reg_2_10_inst : DLH_X1 port map( G => n433, D => n466, Q => 
                           mask_2_10_port);
   mask_reg_2_9_inst : DLH_X1 port map( G => n432, D => n467, Q => 
                           mask_2_9_port);
   mask_reg_2_8_inst : DLH_X1 port map( G => n432, D => n468, Q => 
                           mask_2_8_port);
   mask_reg_2_7_inst : DLH_X1 port map( G => n432, D => n469, Q => 
                           mask_2_7_port);
   mask_reg_2_6_inst : DLH_X1 port map( G => n432, D => N51, Q => mask_2_6_port
                           );
   mask_reg_2_5_inst : DLH_X1 port map( G => n432, D => N50, Q => mask_2_5_port
                           );
   mask_reg_2_4_inst : DLH_X1 port map( G => n432, D => N49, Q => mask_2_4_port
                           );
   mask_reg_2_3_inst : DLH_X1 port map( G => n432, D => N48, Q => mask_2_3_port
                           );
   mask_reg_2_2_inst : DLH_X1 port map( G => n432, D => N47, Q => mask_2_2_port
                           );
   mask_reg_2_1_inst : DLH_X1 port map( G => n432, D => N46, Q => mask_2_1_port
                           );
   mask_reg_2_0_inst : DLH_X1 port map( G => n432, D => N45, Q => mask_2_0_port
                           );
   mask_reg_3_39_inst : DLH_X1 port map( G => n431, D => n452, Q => 
                           mask_3_39_port);
   mask_reg_3_38_inst : DLH_X1 port map( G => n431, D => N43, Q => 
                           mask_3_38_port);
   mask_reg_3_37_inst : DLH_X1 port map( G => n431, D => N42, Q => 
                           mask_3_37_port);
   mask_reg_3_36_inst : DLH_X1 port map( G => n431, D => N41, Q => 
                           mask_3_36_port);
   mask_reg_3_35_inst : DLH_X1 port map( G => n431, D => N40, Q => 
                           mask_3_35_port);
   mask_reg_3_34_inst : DLH_X1 port map( G => n431, D => N39, Q => 
                           mask_3_34_port);
   mask_reg_3_33_inst : DLH_X1 port map( G => n431, D => N38, Q => 
                           mask_3_33_port);
   mask_reg_3_32_inst : DLH_X1 port map( G => n431, D => N37, Q => 
                           mask_3_32_port);
   mask_reg_3_31_inst : DLH_X1 port map( G => n431, D => n390, Q => 
                           mask_3_31_port);
   mask_reg_3_30_inst : DLH_X1 port map( G => n431, D => n390, Q => 
                           mask_3_30_port);
   mask_reg_3_29_inst : DLH_X1 port map( G => n430, D => n390, Q => 
                           mask_3_29_port);
   mask_reg_3_28_inst : DLH_X1 port map( G => n430, D => n390, Q => 
                           mask_3_28_port);
   mask_reg_3_27_inst : DLH_X1 port map( G => n430, D => n390, Q => 
                           mask_3_27_port);
   mask_reg_3_26_inst : DLH_X1 port map( G => n430, D => n390, Q => 
                           mask_3_26_port);
   mask_reg_3_25_inst : DLH_X1 port map( G => n430, D => n391, Q => 
                           mask_3_25_port);
   mask_reg_3_24_inst : DLH_X1 port map( G => n430, D => n391, Q => 
                           mask_3_24_port);
   mask_reg_3_23_inst : DLH_X1 port map( G => n430, D => n391, Q => 
                           mask_3_23_port);
   mask_reg_3_22_inst : DLH_X1 port map( G => n430, D => n391, Q => 
                           mask_3_22_port);
   mask_reg_3_21_inst : DLH_X1 port map( G => n430, D => n391, Q => 
                           mask_3_21_port);
   mask_reg_3_20_inst : DLH_X1 port map( G => n430, D => n391, Q => 
                           mask_3_20_port);
   mask_reg_3_19_inst : DLH_X1 port map( G => n429, D => n391, Q => 
                           mask_3_19_port);
   mask_reg_3_18_inst : DLH_X1 port map( G => n429, D => n391, Q => 
                           mask_3_18_port);
   mask_reg_3_17_inst : DLH_X1 port map( G => n429, D => n391, Q => 
                           mask_3_17_port);
   mask_reg_3_16_inst : DLH_X1 port map( G => n429, D => n390, Q => 
                           mask_3_16_port);
   mask_reg_3_15_inst : DLH_X1 port map( G => n429, D => n391, Q => 
                           mask_3_15_port);
   mask_reg_3_14_inst : DLH_X1 port map( G => n429, D => n392, Q => 
                           mask_3_14_port);
   mask_reg_3_13_inst : DLH_X1 port map( G => n429, D => n392, Q => 
                           mask_3_13_port);
   mask_reg_3_12_inst : DLH_X1 port map( G => n429, D => n392, Q => 
                           mask_3_12_port);
   mask_reg_3_11_inst : DLH_X1 port map( G => n429, D => n392, Q => 
                           mask_3_11_port);
   mask_reg_3_10_inst : DLH_X1 port map( G => n429, D => n392, Q => 
                           mask_3_10_port);
   mask_reg_3_9_inst : DLH_X1 port map( G => n428, D => n392, Q => 
                           mask_3_9_port);
   mask_reg_3_8_inst : DLH_X1 port map( G => n428, D => n397, Q => 
                           mask_3_8_port);
   mask_reg_3_7_inst : DLH_X1 port map( G => n428, D => N35, Q => mask_3_7_port
                           );
   mask_reg_3_6_inst : DLH_X1 port map( G => n428, D => n462, Q => 
                           mask_3_6_port);
   mask_reg_3_5_inst : DLH_X1 port map( G => n428, D => n463, Q => 
                           mask_3_5_port);
   mask_reg_3_4_inst : DLH_X1 port map( G => n428, D => n464, Q => 
                           mask_3_4_port);
   mask_reg_3_3_inst : DLH_X1 port map( G => n428, D => n465, Q => 
                           mask_3_3_port);
   mask_reg_3_2_inst : DLH_X1 port map( G => n428, D => n466, Q => 
                           mask_3_2_port);
   mask_reg_3_1_inst : DLH_X1 port map( G => n428, D => n467, Q => 
                           mask_3_1_port);
   mask_reg_3_0_inst : DLH_X1 port map( G => n428, D => n468, Q => 
                           mask_3_0_port);
   U3 : BUF_X1 port map( A => n91_port, Z => n414);
   U4 : INV_X1 port map( A => R(0), ZN => n338);
   U5 : OR2_X1 port map( A1 => conf(1), A2 => conf(0), ZN => n1);
   U6 : BUF_X1 port map( A => n451, Z => n446);
   U7 : BUF_X1 port map( A => n451, Z => n445);
   U8 : BUF_X1 port map( A => n451, Z => n444);
   U9 : BUF_X1 port map( A => n450, Z => n448);
   U10 : BUF_X1 port map( A => n450, Z => n447);
   U11 : BUF_X1 port map( A => n427, Z => n451);
   U12 : BUF_X1 port map( A => n427, Z => n450);
   U13 : BUF_X1 port map( A => n345, Z => n347);
   U14 : BUF_X1 port map( A => n345, Z => n346);
   U15 : BUF_X1 port map( A => n354, Z => n356);
   U16 : BUF_X1 port map( A => n354, Z => n355);
   U17 : BUF_X1 port map( A => n2, Z => n421);
   U18 : BUF_X1 port map( A => n3, Z => n415);
   U19 : BUF_X1 port map( A => n414, Z => n412);
   U20 : BUF_X1 port map( A => n8, Z => n397);
   U21 : BUF_X1 port map( A => n406, Z => n403);
   U22 : AND2_X1 port map( A1 => R(4), A2 => R(3), ZN => n2);
   U23 : AND2_X1 port map( A1 => R(4), A2 => n532, ZN => n3);
   U24 : BUF_X1 port map( A => n8, Z => n398);
   U25 : BUF_X1 port map( A => n406, Z => n404);
   U26 : BUF_X1 port map( A => n338, Z => n363);
   U27 : BUF_X1 port map( A => n338, Z => n364);
   U28 : NOR2_X1 port map( A1 => n239, A2 => n238, ZN => n229);
   U29 : BUF_X1 port map( A => n1, Z => n406);
   U30 : BUF_X1 port map( A => n407, Z => n402);
   U31 : AND2_X1 port map( A1 => n106, A2 => n107, ZN => n4);
   U32 : AND2_X1 port map( A1 => n146, A2 => n147, ZN => n5);
   U33 : BUF_X1 port map( A => n448, Z => n429);
   U34 : BUF_X1 port map( A => n448, Z => n430);
   U35 : BUF_X1 port map( A => n448, Z => n431);
   U36 : BUF_X1 port map( A => n447, Z => n432);
   U37 : BUF_X1 port map( A => n447, Z => n433);
   U38 : BUF_X1 port map( A => n447, Z => n434);
   U39 : BUF_X1 port map( A => n446, Z => n435);
   U40 : BUF_X1 port map( A => n446, Z => n436);
   U41 : BUF_X1 port map( A => n446, Z => n437);
   U42 : BUF_X1 port map( A => n445, Z => n438);
   U43 : BUF_X1 port map( A => n445, Z => n439);
   U44 : BUF_X1 port map( A => n445, Z => n440);
   U45 : BUF_X1 port map( A => n444, Z => n441);
   U46 : BUF_X1 port map( A => n444, Z => n442);
   U47 : BUF_X1 port map( A => n444, Z => n443);
   U48 : BUF_X1 port map( A => n412, Z => n409);
   U49 : BUF_X1 port map( A => n412, Z => n410);
   U50 : BUF_X1 port map( A => n412, Z => n411);
   U51 : BUF_X1 port map( A => n421, Z => n423);
   U52 : BUF_X1 port map( A => n415, Z => n417);
   U53 : BUF_X1 port map( A => n347, Z => n348);
   U54 : BUF_X1 port map( A => n347, Z => n349);
   U55 : BUF_X1 port map( A => n421, Z => n424);
   U56 : BUF_X1 port map( A => n415, Z => n419);
   U57 : BUF_X1 port map( A => n415, Z => n418);
   U58 : BUF_X1 port map( A => n421, Z => n425);
   U59 : BUF_X1 port map( A => n346, Z => n351);
   U60 : BUF_X1 port map( A => n346, Z => n352);
   U61 : BUF_X1 port map( A => n347, Z => n350);
   U62 : BUF_X1 port map( A => n346, Z => n353);
   U63 : BUF_X1 port map( A => n356, Z => n358);
   U64 : BUF_X1 port map( A => n356, Z => n359);
   U65 : BUF_X1 port map( A => n356, Z => n357);
   U66 : BUF_X1 port map( A => n355, Z => n360);
   U67 : BUF_X1 port map( A => n355, Z => n361);
   U68 : BUF_X1 port map( A => n355, Z => n362);
   U69 : BUF_X1 port map( A => n449, Z => n428);
   U70 : BUF_X1 port map( A => n450, Z => n449);
   U71 : INV_X1 port map( A => n189_port, ZN => data_out(21));
   U72 : INV_X1 port map( A => n188_port, ZN => data_out(22));
   U73 : INV_X1 port map( A => n185_port, ZN => data_out(25));
   U74 : AOI22_X1 port map( A1 => N184, A2 => n400, B1 => N216, B2 => n393, ZN 
                           => n184_port);
   U75 : INV_X1 port map( A => n179_port, ZN => data_out(30));
   U76 : AOI22_X1 port map( A1 => N188, A2 => n399, B1 => N220, B2 => n403, ZN 
                           => n179_port);
   U77 : INV_X1 port map( A => n181_port, ZN => data_out(29));
   U78 : AOI22_X1 port map( A1 => N187, A2 => n399, B1 => N219, B2 => n403, ZN 
                           => n181_port);
   U79 : BUF_X1 port map( A => n416, Z => n420);
   U80 : BUF_X1 port map( A => n3, Z => n416);
   U81 : BUF_X1 port map( A => n413, Z => n408);
   U82 : CLKBUF_X1 port map( A => n414, Z => n413);
   U83 : BUF_X1 port map( A => n422, Z => n426);
   U84 : BUF_X1 port map( A => n2, Z => n422);
   U85 : INV_X1 port map( A => n342, ZN => n344);
   U86 : INV_X1 port map( A => n342, ZN => n343);
   U87 : BUF_X1 port map( A => n363, Z => n370);
   U88 : BUF_X1 port map( A => n363, Z => n369);
   U89 : BUF_X1 port map( A => n363, Z => n368);
   U90 : BUF_X1 port map( A => n364, Z => n367);
   U91 : BUF_X1 port map( A => n364, Z => n366);
   U92 : BUF_X1 port map( A => n364, Z => n365);
   U93 : BUF_X1 port map( A => n340, Z => n341);
   U94 : INV_X1 port map( A => n6, ZN => n373);
   U95 : INV_X1 port map( A => n6, ZN => n372);
   U96 : INV_X1 port map( A => n6, ZN => n371);
   U97 : INV_X1 port map( A => n7, ZN => n376);
   U98 : INV_X1 port map( A => n7, ZN => n375);
   U99 : INV_X1 port map( A => n7, ZN => n374);
   U100 : NAND2_X1 port map( A1 => n227, A2 => n216_port, ZN => N69);
   U101 : NAND2_X1 port map( A1 => n226, A2 => n214_port, ZN => N70);
   U102 : NAND2_X1 port map( A1 => n225, A2 => n212_port, ZN => N71);
   U103 : NAND2_X1 port map( A1 => n224, A2 => n210_port, ZN => N72);
   U104 : NAND2_X1 port map( A1 => n223, A2 => n208_port, ZN => N73);
   U105 : NAND2_X1 port map( A1 => n222, A2 => n206_port, ZN => N74);
   U106 : NAND2_X1 port map( A1 => n221_port, A2 => n204_port, ZN => N75);
   U107 : NAND2_X1 port map( A1 => n396, A2 => n216_port, ZN => N37);
   U108 : NAND2_X1 port map( A1 => n396, A2 => n214_port, ZN => N38);
   U109 : NAND2_X1 port map( A1 => n396, A2 => n212_port, ZN => N39);
   U110 : NAND2_X1 port map( A1 => n396, A2 => n210_port, ZN => N40);
   U111 : NAND2_X1 port map( A1 => n396, A2 => n208_port, ZN => N41);
   U112 : NAND2_X1 port map( A1 => n396, A2 => n206_port, ZN => N42);
   U113 : NAND2_X1 port map( A1 => n396, A2 => n204_port, ZN => N43);
   U114 : INV_X1 port map( A => n227, ZN => n468);
   U115 : INV_X1 port map( A => n226, ZN => n467);
   U116 : INV_X1 port map( A => n225, ZN => n466);
   U117 : INV_X1 port map( A => n224, ZN => n465);
   U118 : INV_X1 port map( A => n223, ZN => n464);
   U119 : INV_X1 port map( A => n222, ZN => n463);
   U120 : INV_X1 port map( A => n221_port, ZN => n462);
   U121 : NAND2_X1 port map( A1 => n215_port, A2 => n216_port, ZN => N93);
   U122 : NAND2_X1 port map( A1 => n213_port, A2 => n214_port, ZN => N94);
   U123 : NAND2_X1 port map( A1 => n211_port, A2 => n212_port, ZN => N95);
   U124 : NAND2_X1 port map( A1 => n209_port, A2 => n210_port, ZN => N96);
   U125 : NAND2_X1 port map( A1 => n207_port, A2 => n208_port, ZN => N97);
   U126 : NAND2_X1 port map( A1 => n205_port, A2 => n206_port, ZN => N98);
   U127 : NAND2_X1 port map( A1 => n203_port, A2 => n204_port, ZN => N99);
   U128 : INV_X1 port map( A => n228, ZN => n469);
   U129 : INV_X1 port map( A => n220_port, ZN => n452);
   U130 : INV_X1 port map( A => n215_port, ZN => n499);
   U131 : INV_X1 port map( A => n213_port, ZN => n497);
   U132 : INV_X1 port map( A => n211_port, ZN => n495);
   U133 : INV_X1 port map( A => n209_port, ZN => n493);
   U134 : INV_X1 port map( A => n207_port, ZN => n491);
   U135 : INV_X1 port map( A => n205_port, ZN => n489);
   U136 : INV_X1 port map( A => n203_port, ZN => n487);
   U137 : BUF_X1 port map( A => n404, Z => n394);
   U138 : INV_X1 port map( A => n217_port, ZN => n461);
   U139 : BUF_X1 port map( A => n404, Z => n395);
   U140 : INV_X1 port map( A => n397, ZN => n396);
   U141 : BUF_X1 port map( A => n404, Z => n393);
   U142 : INV_X1 port map( A => n403, ZN => n400);
   U143 : INV_X1 port map( A => n403, ZN => n399);
   U144 : BUF_X1 port map( A => n398, Z => n391);
   U145 : BUF_X1 port map( A => n398, Z => n390);
   U146 : BUF_X1 port map( A => n398, Z => n392);
   U147 : INV_X1 port map( A => n190_port, ZN => data_out(20));
   U148 : INV_X1 port map( A => n183_port, ZN => data_out(27));
   U149 : AOI22_X1 port map( A1 => N186, A2 => n399, B1 => N218, B2 => n403, ZN
                           => n182_port);
   U150 : AOI22_X1 port map( A1 => N182, A2 => n400, B1 => N214, B2 => n393, ZN
                           => n186_port);
   U151 : AOI22_X1 port map( A1 => N189, A2 => n399, B1 => N221, B2 => n403, ZN
                           => n178_port);
   U152 : NOR2_X1 port map( A1 => R(3), A2 => R(4), ZN => n91_port);
   U153 : INV_X1 port map( A => n193_port, ZN => data_out(18));
   U154 : INV_X1 port map( A => n197_port, ZN => data_out(14));
   U155 : AOI22_X1 port map( A1 => N172, A2 => n400, B1 => N204, B2 => n393, ZN
                           => n197_port);
   U156 : INV_X1 port map( A => n196_port, ZN => data_out(15));
   U157 : INV_X1 port map( A => n194_port, ZN => data_out(17));
   U158 : INV_X1 port map( A => n195_port, ZN => data_out(16));
   U159 : AOI22_X1 port map( A1 => N174, A2 => n400, B1 => N206, B2 => n393, ZN
                           => n195_port);
   U160 : AOI22_X1 port map( A1 => N159, A2 => n400, B1 => N191, B2 => n393, ZN
                           => n191_port);
   U161 : INV_X1 port map( A => n199_port, ZN => data_out(12));
   U162 : AOI22_X1 port map( A1 => N170, A2 => n399, B1 => N202, B2 => n394, ZN
                           => n199_port);
   U163 : AOI22_X1 port map( A1 => N177, A2 => n400, B1 => N209, B2 => n393, ZN
                           => n192_port);
   U164 : INV_X1 port map( A => n200_port, ZN => data_out(11));
   U165 : INV_X1 port map( A => n176_port, ZN => data_out(4));
   U166 : INV_X1 port map( A => n177_port, ZN => data_out(3));
   U167 : AOI22_X1 port map( A1 => N171, A2 => n401, B1 => N203, B2 => n394, ZN
                           => n198_port);
   U168 : INV_X1 port map( A => n174_port, ZN => data_out(6));
   U169 : AOI22_X1 port map( A1 => N169, A2 => n400, B1 => N201, B2 => n394, ZN
                           => n200_port);
   U170 : INV_X1 port map( A => n175_port, ZN => data_out(5));
   U171 : AOI22_X1 port map( A1 => N165, A2 => n399, B1 => N197, B2 => n403, ZN
                           => n173_port);
   U172 : AOI22_X1 port map( A1 => N167, A2 => n399, B1 => N199, B2 => n394, ZN
                           => n170_port);
   U173 : AOI22_X1 port map( A1 => N168, A2 => n401, B1 => N200, B2 => n394, ZN
                           => n201_port);
   U174 : BUF_X1 port map( A => n297, Z => n345);
   U175 : INV_X1 port map( A => R(2), ZN => n301);
   U176 : BUF_X1 port map( A => n298, Z => n354);
   U177 : BUF_X1 port map( A => n339, Z => n342);
   U178 : BUF_X1 port map( A => n338, Z => n339);
   U179 : AND2_X1 port map( A1 => R(1), A2 => n301, ZN => n6);
   U180 : AND2_X1 port map( A1 => R(1), A2 => R(2), ZN => n7);
   U181 : INV_X1 port map( A => n229, ZN => n533);
   U182 : AOI21_X1 port map( B1 => n401, B2 => data_in(7), A => n397, ZN => 
                           n220_port);
   U183 : AOI21_X1 port map( B1 => n401, B2 => data_in(23), A => n397, ZN => 
                           n217_port);
   U184 : NAND2_X1 port map( A1 => data_in(24), A2 => n533, ZN => n227);
   U185 : NAND2_X1 port map( A1 => data_in(25), A2 => n533, ZN => n226);
   U186 : NAND2_X1 port map( A1 => data_in(26), A2 => n533, ZN => n225);
   U187 : NAND2_X1 port map( A1 => data_in(27), A2 => n533, ZN => n224);
   U188 : NAND2_X1 port map( A1 => data_in(28), A2 => n533, ZN => n223);
   U189 : NAND2_X1 port map( A1 => data_in(29), A2 => n533, ZN => n222);
   U190 : NAND2_X1 port map( A1 => data_in(30), A2 => n533, ZN => n221_port);
   U191 : NOR2_X1 port map( A1 => n483, A2 => n229, ZN => N45);
   U192 : NOR2_X1 port map( A1 => n481, A2 => n229, ZN => N46);
   U193 : NOR2_X1 port map( A1 => n479, A2 => n229, ZN => N47);
   U194 : NOR2_X1 port map( A1 => n477, A2 => n229, ZN => N48);
   U195 : NOR2_X1 port map( A1 => n475, A2 => n229, ZN => N49);
   U196 : NOR2_X1 port map( A1 => n473, A2 => n229, ZN => N50);
   U197 : NOR2_X1 port map( A1 => n471, A2 => n229, ZN => N51);
   U198 : NAND2_X1 port map( A1 => data_in(8), A2 => n533, ZN => n215_port);
   U199 : NAND2_X1 port map( A1 => data_in(9), A2 => n533, ZN => n213_port);
   U200 : NAND2_X1 port map( A1 => data_in(10), A2 => n533, ZN => n211_port);
   U201 : NAND2_X1 port map( A1 => data_in(11), A2 => n533, ZN => n209_port);
   U202 : NAND2_X1 port map( A1 => data_in(12), A2 => n533, ZN => n207_port);
   U203 : NAND2_X1 port map( A1 => data_in(13), A2 => n533, ZN => n205_port);
   U204 : NAND2_X1 port map( A1 => data_in(14), A2 => n533, ZN => n203_port);
   U205 : NAND2_X1 port map( A1 => data_in(23), A2 => n533, ZN => n228);
   U206 : NOR2_X1 port map( A1 => n485, A2 => n229, ZN => N68);
   U207 : NAND2_X1 port map( A1 => data_in(0), A2 => n401, ZN => n216_port);
   U208 : NAND2_X1 port map( A1 => data_in(1), A2 => n401, ZN => n214_port);
   U209 : NAND2_X1 port map( A1 => data_in(2), A2 => n401, ZN => n212_port);
   U210 : NAND2_X1 port map( A1 => data_in(3), A2 => n401, ZN => n210_port);
   U211 : NAND2_X1 port map( A1 => data_in(4), A2 => n400, ZN => n208_port);
   U212 : NAND2_X1 port map( A1 => data_in(5), A2 => n399, ZN => n206_port);
   U213 : NAND2_X1 port map( A1 => data_in(6), A2 => n401, ZN => n204_port);
   U214 : OAI21_X1 port map( B1 => n395, B2 => n498, A => n396, ZN => N53);
   U215 : INV_X1 port map( A => data_in(8), ZN => n498);
   U216 : OAI21_X1 port map( B1 => n395, B2 => n496, A => n396, ZN => N54);
   U217 : INV_X1 port map( A => data_in(9), ZN => n496);
   U218 : OAI21_X1 port map( B1 => n395, B2 => n494, A => n396, ZN => N55);
   U219 : INV_X1 port map( A => data_in(10), ZN => n494);
   U220 : OAI21_X1 port map( B1 => n395, B2 => n492, A => n396, ZN => N56);
   U221 : INV_X1 port map( A => data_in(11), ZN => n492);
   U222 : OAI21_X1 port map( B1 => n395, B2 => n490, A => n396, ZN => N57);
   U223 : INV_X1 port map( A => data_in(12), ZN => n490);
   U224 : OAI21_X1 port map( B1 => n395, B2 => n488, A => n396, ZN => N58);
   U225 : INV_X1 port map( A => data_in(13), ZN => n488);
   U226 : OAI21_X1 port map( B1 => n395, B2 => n486, A => n396, ZN => N59);
   U227 : INV_X1 port map( A => data_in(14), ZN => n486);
   U228 : OAI21_X1 port map( B1 => n395, B2 => n485, A => n396, ZN => N60);
   U229 : OAI21_X1 port map( B1 => n395, B2 => n483, A => n396, ZN => N77);
   U230 : OAI21_X1 port map( B1 => n394, B2 => n481, A => n396, ZN => N78);
   U231 : OAI21_X1 port map( B1 => n394, B2 => n479, A => n396, ZN => N79);
   U232 : OAI21_X1 port map( B1 => n394, B2 => n477, A => n396, ZN => N80);
   U233 : OAI21_X1 port map( B1 => n394, B2 => n475, A => n396, ZN => N81);
   U234 : OAI21_X1 port map( B1 => n394, B2 => n473, A => n396, ZN => N82);
   U235 : OAI21_X1 port map( B1 => n394, B2 => n471, A => n396, ZN => N83);
   U236 : OAI21_X1 port map( B1 => n405, B2 => n485, A => n228, ZN => N108);
   U237 : OAI21_X1 port map( B1 => n405, B2 => n483, A => n227, ZN => N109);
   U238 : OAI21_X1 port map( B1 => n405, B2 => n481, A => n226, ZN => N110);
   U239 : OAI21_X1 port map( B1 => n405, B2 => n479, A => n225, ZN => N111);
   U240 : OAI21_X1 port map( B1 => n405, B2 => n477, A => n224, ZN => N112);
   U241 : OAI21_X1 port map( B1 => n405, B2 => n475, A => n223, ZN => N113);
   U242 : OAI21_X1 port map( B1 => n405, B2 => n473, A => n222, ZN => N114);
   U243 : OAI21_X1 port map( B1 => n395, B2 => n471, A => n221_port, ZN => N115
                           );
   U244 : NAND2_X1 port map( A1 => n396, A2 => n219_port, ZN => N35);
   U245 : AND2_X1 port map( A1 => n533, A2 => data_in(0), ZN => N85);
   U246 : AND2_X1 port map( A1 => n533, A2 => data_in(1), ZN => N86);
   U247 : AND2_X1 port map( A1 => n533, A2 => data_in(2), ZN => N87);
   U248 : AND2_X1 port map( A1 => n533, A2 => data_in(3), ZN => N88);
   U249 : AND2_X1 port map( A1 => n533, A2 => data_in(4), ZN => N89);
   U250 : AND2_X1 port map( A1 => n533, A2 => data_in(5), ZN => N90);
   U251 : AND2_X1 port map( A1 => n533, A2 => data_in(6), ZN => N91);
   U252 : AND2_X1 port map( A1 => n533, A2 => data_in(7), ZN => N92);
   U253 : BUF_X1 port map( A => N28, Z => n427);
   U254 : NAND2_X1 port map( A1 => n229, A2 => n403, ZN => N28);
   U255 : NAND2_X1 port map( A1 => n219_port, A2 => n220_port, ZN => N76);
   U256 : NAND2_X1 port map( A1 => n219_port, A2 => n217_port, ZN => N116);
   U257 : INV_X1 port map( A => n402, ZN => n401);
   U258 : BUF_X1 port map( A => n406, Z => n405);
   U259 : INV_X1 port map( A => n247, ZN => n484);
   U260 : AOI21_X1 port map( B1 => n400, B2 => data_in(7), A => N68, ZN => n247
                           );
   U261 : INV_X1 port map( A => n246, ZN => n482);
   U262 : AOI21_X1 port map( B1 => n400, B2 => data_in(8), A => N45, ZN => n246
                           );
   U263 : INV_X1 port map( A => n245, ZN => n480);
   U264 : AOI21_X1 port map( B1 => n399, B2 => data_in(9), A => N46, ZN => n245
                           );
   U265 : INV_X1 port map( A => n244, ZN => n478);
   U266 : AOI21_X1 port map( B1 => n401, B2 => data_in(10), A => N47, ZN => 
                           n244);
   U267 : INV_X1 port map( A => n243, ZN => n476);
   U268 : AOI21_X1 port map( B1 => n399, B2 => data_in(11), A => N48, ZN => 
                           n243);
   U269 : INV_X1 port map( A => n242, ZN => n474);
   U270 : AOI21_X1 port map( B1 => n400, B2 => data_in(12), A => N49, ZN => 
                           n242);
   U271 : INV_X1 port map( A => n241, ZN => n472);
   U272 : AOI21_X1 port map( B1 => n399, B2 => data_in(13), A => N50, ZN => 
                           n241);
   U273 : INV_X1 port map( A => n240, ZN => n470);
   U274 : AOI21_X1 port map( B1 => n401, B2 => data_in(14), A => N51, ZN => 
                           n240);
   U275 : INV_X1 port map( A => n237, ZN => n460);
   U276 : AOI21_X1 port map( B1 => n401, B2 => data_in(24), A => n397, ZN => 
                           n237);
   U277 : INV_X1 port map( A => n236, ZN => n459);
   U278 : AOI21_X1 port map( B1 => n401, B2 => data_in(25), A => n397, ZN => 
                           n236);
   U279 : INV_X1 port map( A => n235, ZN => n458);
   U280 : AOI21_X1 port map( B1 => n401, B2 => data_in(26), A => n397, ZN => 
                           n235);
   U281 : INV_X1 port map( A => n234, ZN => n457);
   U282 : AOI21_X1 port map( B1 => n401, B2 => data_in(27), A => n397, ZN => 
                           n234);
   U283 : INV_X1 port map( A => n233, ZN => n456);
   U284 : AOI21_X1 port map( B1 => n401, B2 => data_in(28), A => n397, ZN => 
                           n233);
   U285 : INV_X1 port map( A => n232, ZN => n455);
   U286 : AOI21_X1 port map( B1 => n401, B2 => data_in(29), A => n397, ZN => 
                           n232);
   U287 : INV_X1 port map( A => n231, ZN => n454);
   U288 : AOI21_X1 port map( B1 => n401, B2 => data_in(30), A => n397, ZN => 
                           n231);
   U289 : INV_X1 port map( A => n230, ZN => n453);
   U290 : AOI21_X1 port map( B1 => n401, B2 => data_in(31), A => n397, ZN => 
                           n230);
   U291 : INV_X1 port map( A => out_mask_23_port, ZN => n324);
   U292 : INV_X1 port map( A => out_mask_25_port, ZN => n322);
   U293 : INV_X1 port map( A => out_mask_26_port, ZN => n321);
   U294 : INV_X1 port map( A => out_mask_27_port, ZN => n320);
   U295 : INV_X1 port map( A => out_mask_22_port, ZN => n325);
   U296 : INV_X1 port map( A => out_mask_24_port, ZN => n323);
   U297 : INV_X1 port map( A => out_mask_34_port, ZN => n312);
   U298 : INV_X1 port map( A => out_mask_32_port, ZN => n314);
   U299 : INV_X1 port map( A => out_mask_20_port, ZN => n327);
   U300 : INV_X1 port map( A => out_mask_30_port, ZN => n316);
   U301 : INV_X1 port map( A => out_mask_21_port, ZN => n326);
   U302 : INV_X1 port map( A => out_mask_29_port, ZN => n318);
   U303 : INV_X1 port map( A => out_mask_31_port, ZN => n315);
   U304 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => out_mask_39_port);
   U305 : INV_X1 port map( A => out_mask_33_port, ZN => n313);
   U306 : INV_X1 port map( A => out_mask_28_port, ZN => n319);
   U307 : AOI22_X1 port map( A1 => N158, A2 => n400, B1 => N190, B2 => n394, ZN
                           => n202_port);
   U308 : INV_X1 port map( A => out_mask_5_port, ZN => n306);
   U309 : INV_X1 port map( A => out_mask_2_port, ZN => n317);
   U310 : INV_X1 port map( A => out_mask_6_port, ZN => n305);
   U311 : INV_X1 port map( A => out_mask_36_port, ZN => n310);
   U312 : INV_X1 port map( A => out_mask_4_port, ZN => n307);
   U313 : INV_X1 port map( A => out_mask_7_port, ZN => n304);
   U314 : INV_X1 port map( A => out_mask_8_port, ZN => n303);
   U315 : INV_X1 port map( A => out_mask_9_port, ZN => n302);
   U316 : INV_X1 port map( A => out_mask_35_port, ZN => n311);
   U317 : INV_X1 port map( A => out_mask_3_port, ZN => n308);
   U318 : INV_X1 port map( A => out_mask_37_port, ZN => n309);
   U319 : INV_X1 port map( A => out_mask_19_port, ZN => n328);
   U320 : INV_X1 port map( A => out_mask_16_port, ZN => n331);
   U321 : INV_X1 port map( A => out_mask_15_port, ZN => n332);
   U322 : INV_X1 port map( A => out_mask_18_port, ZN => n329);
   U323 : INV_X1 port map( A => out_mask_10_port, ZN => n337);
   U324 : INV_X1 port map( A => out_mask_11_port, ZN => n336);
   U325 : INV_X1 port map( A => out_mask_12_port, ZN => n335);
   U326 : INV_X1 port map( A => out_mask_17_port, ZN => n330);
   U327 : INV_X1 port map( A => out_mask_14_port, ZN => n333);
   U328 : INV_X1 port map( A => out_mask_13_port, ZN => n334);
   U329 : NAND2_X1 port map( A1 => n239, A2 => data_in(31), ZN => n219_port);
   U330 : INV_X1 port map( A => data_in(15), ZN => n485);
   U331 : INV_X1 port map( A => data_in(16), ZN => n483);
   U332 : INV_X1 port map( A => data_in(17), ZN => n481);
   U333 : INV_X1 port map( A => data_in(18), ZN => n479);
   U334 : INV_X1 port map( A => data_in(19), ZN => n477);
   U335 : INV_X1 port map( A => data_in(20), ZN => n475);
   U336 : INV_X1 port map( A => data_in(21), ZN => n473);
   U337 : INV_X1 port map( A => data_in(22), ZN => n471);
   U338 : BUF_X1 port map( A => n1, Z => n407);
   U339 : AND2_X1 port map( A1 => data_in(31), A2 => n238, ZN => n8);
   U340 : NAND2_X1 port map( A1 => n138, A2 => n139, ZN => out_mask_23_port);
   U341 : AOI22_X1 port map( A1 => mask_3_23_port, A2 => n424, B1 => 
                           mask_2_23_port, B2 => n418, ZN => n139);
   U342 : AOI22_X1 port map( A1 => mask_1_23_port, A2 => n382, B1 => 
                           mask_0_23_port, B2 => n409, ZN => n138);
   U343 : NAND2_X1 port map( A1 => n134, A2 => n135, ZN => out_mask_25_port);
   U344 : AOI22_X1 port map( A1 => mask_3_25_port, A2 => n424, B1 => 
                           mask_2_25_port, B2 => n418, ZN => n135);
   U345 : AOI22_X1 port map( A1 => mask_1_25_port, A2 => n384, B1 => 
                           mask_0_25_port, B2 => n409, ZN => n134);
   U346 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => out_mask_26_port);
   U347 : AOI22_X1 port map( A1 => mask_3_26_port, A2 => n424, B1 => 
                           mask_2_26_port, B2 => n418, ZN => n133);
   U348 : AOI22_X1 port map( A1 => mask_1_26_port, A2 => n382, B1 => 
                           mask_0_26_port, B2 => n409, ZN => n132);
   U349 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => out_mask_27_port);
   U350 : AOI22_X1 port map( A1 => mask_3_27_port, A2 => n424, B1 => 
                           mask_2_27_port, B2 => n418, ZN => n131);
   U351 : AOI22_X1 port map( A1 => mask_1_27_port, A2 => n383, B1 => 
                           mask_0_27_port, B2 => n409, ZN => n130);
   U352 : NAND2_X1 port map( A1 => n140, A2 => n141, ZN => out_mask_22_port);
   U353 : AOI22_X1 port map( A1 => mask_3_22_port, A2 => n424, B1 => 
                           mask_2_22_port, B2 => n418, ZN => n141);
   U354 : AOI22_X1 port map( A1 => mask_1_22_port, A2 => n90_port, B1 => 
                           mask_0_22_port, B2 => n409, ZN => n140);
   U355 : NAND2_X1 port map( A1 => n136, A2 => n137, ZN => out_mask_24_port);
   U356 : AOI22_X1 port map( A1 => mask_3_24_port, A2 => n424, B1 => 
                           mask_2_24_port, B2 => n418, ZN => n137);
   U357 : AOI22_X1 port map( A1 => mask_1_24_port, A2 => n383, B1 => 
                           mask_0_24_port, B2 => n409, ZN => n136);
   U358 : NAND2_X1 port map( A1 => n114_port, A2 => n115_port, ZN => 
                           out_mask_34_port);
   U359 : AOI22_X1 port map( A1 => mask_3_34_port, A2 => n425, B1 => 
                           mask_2_34_port, B2 => n419, ZN => n115_port);
   U360 : AOI22_X1 port map( A1 => mask_1_34_port, A2 => n380, B1 => 
                           mask_0_34_port, B2 => n410, ZN => n114_port);
   U361 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => out_mask_32_port);
   U362 : AOI22_X1 port map( A1 => mask_3_32_port, A2 => n425, B1 => 
                           mask_2_32_port, B2 => n419, ZN => n119);
   U363 : AOI22_X1 port map( A1 => mask_1_32_port, A2 => n385, B1 => 
                           mask_0_32_port, B2 => n410, ZN => n118);
   U364 : NAND2_X1 port map( A1 => n144, A2 => n145, ZN => out_mask_20_port);
   U365 : AOI22_X1 port map( A1 => mask_3_20_port, A2 => n424, B1 => 
                           mask_2_20_port, B2 => n418, ZN => n145);
   U366 : AOI22_X1 port map( A1 => mask_1_20_port, A2 => n386, B1 => 
                           mask_0_20_port, B2 => n409, ZN => n144);
   U367 : NAND2_X1 port map( A1 => n122, A2 => n123, ZN => out_mask_30_port);
   U368 : AOI22_X1 port map( A1 => mask_3_30_port, A2 => n424, B1 => 
                           mask_2_30_port, B2 => n418, ZN => n123);
   U369 : AOI22_X1 port map( A1 => mask_1_30_port, A2 => n381, B1 => 
                           mask_0_30_port, B2 => n409, ZN => n122);
   U370 : NAND2_X1 port map( A1 => n142, A2 => n143, ZN => out_mask_21_port);
   U371 : AOI22_X1 port map( A1 => mask_3_21_port, A2 => n424, B1 => 
                           mask_2_21_port, B2 => n418, ZN => n143);
   U372 : AOI22_X1 port map( A1 => mask_1_21_port, A2 => n389, B1 => 
                           mask_0_21_port, B2 => n409, ZN => n142);
   U373 : NAND2_X1 port map( A1 => n126, A2 => n127, ZN => out_mask_29_port);
   U374 : AOI22_X1 port map( A1 => mask_3_29_port, A2 => n424, B1 => 
                           mask_2_29_port, B2 => n418, ZN => n127);
   U375 : AOI22_X1 port map( A1 => mask_1_29_port, A2 => n379, B1 => 
                           mask_0_29_port, B2 => n409, ZN => n126);
   U376 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => out_mask_31_port);
   U377 : AOI22_X1 port map( A1 => mask_3_31_port, A2 => n425, B1 => 
                           mask_2_31_port, B2 => n419, ZN => n121);
   U378 : AOI22_X1 port map( A1 => mask_1_31_port, A2 => n381, B1 => 
                           mask_0_31_port, B2 => n410, ZN => n120);
   U379 : NAND2_X1 port map( A1 => n116_port, A2 => n117, ZN => 
                           out_mask_33_port);
   U380 : AOI22_X1 port map( A1 => mask_3_33_port, A2 => n425, B1 => 
                           mask_2_33_port, B2 => n419, ZN => n117);
   U381 : AOI22_X1 port map( A1 => mask_1_33_port, A2 => n387, B1 => 
                           mask_0_33_port, B2 => n410, ZN => n116_port);
   U382 : NAND2_X1 port map( A1 => n128, A2 => n129, ZN => out_mask_28_port);
   U383 : AOI22_X1 port map( A1 => mask_3_28_port, A2 => n424, B1 => 
                           mask_2_28_port, B2 => n418, ZN => n129);
   U384 : AOI22_X1 port map( A1 => mask_1_28_port, A2 => n389, B1 => 
                           mask_0_28_port, B2 => n409, ZN => n128);
   U385 : NAND2_X1 port map( A1 => n98_port, A2 => n99_port, ZN => 
                           out_mask_5_port);
   U386 : AOI22_X1 port map( A1 => mask_3_5_port, A2 => n425, B1 => 
                           mask_2_5_port, B2 => n419, ZN => n99_port);
   U387 : AOI22_X1 port map( A1 => mask_1_5_port, A2 => n388, B1 => 
                           mask_0_5_port, B2 => n410, ZN => n98_port);
   U388 : NAND2_X1 port map( A1 => n168_port, A2 => n169_port, ZN => 
                           out_mask_0_port);
   U389 : AOI22_X1 port map( A1 => mask_3_0_port, A2 => n423, B1 => 
                           mask_2_0_port, B2 => n417, ZN => n169_port);
   U390 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => out_mask_2_port);
   U391 : AOI22_X1 port map( A1 => mask_3_2_port, A2 => n424, B1 => 
                           mask_2_2_port, B2 => n418, ZN => n125);
   U392 : AOI22_X1 port map( A1 => mask_1_2_port, A2 => n380, B1 => 
                           mask_0_2_port, B2 => n409, ZN => n124);
   U393 : NAND2_X1 port map( A1 => n96_port, A2 => n97_port, ZN => 
                           out_mask_6_port);
   U394 : AOI22_X1 port map( A1 => mask_3_6_port, A2 => n426, B1 => 
                           mask_2_6_port, B2 => n420, ZN => n97_port);
   U395 : AOI22_X1 port map( A1 => mask_1_6_port, A2 => n379, B1 => 
                           mask_0_6_port, B2 => n411, ZN => n96_port);
   U396 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => out_mask_4_port);
   U397 : AOI22_X1 port map( A1 => mask_3_4_port, A2 => n425, B1 => 
                           mask_2_4_port, B2 => n419, ZN => n101);
   U398 : AOI22_X1 port map( A1 => mask_1_4_port, A2 => n387, B1 => 
                           mask_0_4_port, B2 => n410, ZN => n100);
   U399 : NAND2_X1 port map( A1 => n94_port, A2 => n95_port, ZN => 
                           out_mask_7_port);
   U400 : AOI22_X1 port map( A1 => mask_3_7_port, A2 => n426, B1 => 
                           mask_2_7_port, B2 => n420, ZN => n95_port);
   U401 : AOI22_X1 port map( A1 => mask_1_7_port, A2 => n381, B1 => 
                           mask_0_7_port, B2 => n411, ZN => n94_port);
   U402 : AOI22_X1 port map( A1 => mask_3_38_port, A2 => n425, B1 => 
                           mask_2_38_port, B2 => n419, ZN => n107);
   U403 : AOI22_X1 port map( A1 => mask_1_38_port, A2 => n387, B1 => 
                           mask_0_38_port, B2 => n410, ZN => n106);
   U404 : NAND2_X1 port map( A1 => n92_port, A2 => n93_port, ZN => 
                           out_mask_8_port);
   U405 : AOI22_X1 port map( A1 => mask_3_8_port, A2 => n426, B1 => 
                           mask_2_8_port, B2 => n420, ZN => n93_port);
   U406 : AOI22_X1 port map( A1 => mask_1_8_port, A2 => n385, B1 => 
                           mask_0_8_port, B2 => n411, ZN => n92_port);
   U407 : NAND2_X1 port map( A1 => n86_port, A2 => n87_port, ZN => 
                           out_mask_9_port);
   U408 : AOI22_X1 port map( A1 => mask_3_9_port, A2 => n426, B1 => 
                           mask_2_9_port, B2 => n420, ZN => n87_port);
   U409 : AOI22_X1 port map( A1 => mask_1_9_port, A2 => n384, B1 => 
                           mask_0_9_port, B2 => n411, ZN => n86_port);
   U410 : NAND2_X1 port map( A1 => n112_port, A2 => n113_port, ZN => 
                           out_mask_35_port);
   U411 : AOI22_X1 port map( A1 => mask_3_35_port, A2 => n425, B1 => 
                           mask_2_35_port, B2 => n419, ZN => n113_port);
   U412 : AOI22_X1 port map( A1 => mask_1_35_port, A2 => n383, B1 => 
                           mask_0_35_port, B2 => n410, ZN => n112_port);
   U413 : NAND2_X1 port map( A1 => n108_port, A2 => n109_port, ZN => 
                           out_mask_37_port);
   U414 : AOI22_X1 port map( A1 => mask_3_37_port, A2 => n425, B1 => 
                           mask_2_37_port, B2 => n419, ZN => n109_port);
   U415 : AOI22_X1 port map( A1 => mask_1_37_port, A2 => n389, B1 => 
                           mask_0_37_port, B2 => n410, ZN => n108_port);
   U416 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => out_mask_3_port);
   U417 : AOI22_X1 port map( A1 => mask_3_3_port, A2 => n425, B1 => 
                           mask_2_3_port, B2 => n419, ZN => n103);
   U418 : AOI22_X1 port map( A1 => mask_1_3_port, A2 => n388, B1 => 
                           mask_0_3_port, B2 => n410, ZN => n102);
   U419 : NAND2_X1 port map( A1 => n148, A2 => n149, ZN => out_mask_19_port);
   U420 : AOI22_X1 port map( A1 => mask_3_19_port, A2 => n423, B1 => 
                           mask_2_19_port, B2 => n417, ZN => n149);
   U421 : AOI22_X1 port map( A1 => mask_1_19_port, A2 => n386, B1 => 
                           mask_0_19_port, B2 => n408, ZN => n148);
   U422 : NAND2_X1 port map( A1 => n154, A2 => n155, ZN => out_mask_16_port);
   U423 : AOI22_X1 port map( A1 => mask_3_16_port, A2 => n423, B1 => 
                           mask_2_16_port, B2 => n417, ZN => n155);
   U424 : AOI22_X1 port map( A1 => mask_1_16_port, A2 => n379, B1 => 
                           mask_0_16_port, B2 => n408, ZN => n154);
   U425 : NAND2_X1 port map( A1 => n156, A2 => n157, ZN => out_mask_15_port);
   U426 : AOI22_X1 port map( A1 => mask_3_15_port, A2 => n423, B1 => 
                           mask_2_15_port, B2 => n417, ZN => n157);
   U427 : AOI22_X1 port map( A1 => mask_1_15_port, A2 => n389, B1 => 
                           mask_0_15_port, B2 => n408, ZN => n156);
   U428 : NAND2_X1 port map( A1 => n150, A2 => n151, ZN => out_mask_18_port);
   U429 : AOI22_X1 port map( A1 => mask_3_18_port, A2 => n423, B1 => 
                           mask_2_18_port, B2 => n417, ZN => n151);
   U430 : AOI22_X1 port map( A1 => mask_1_18_port, A2 => n385, B1 => 
                           mask_0_18_port, B2 => n408, ZN => n150);
   U431 : NAND2_X1 port map( A1 => n166_port, A2 => n167_port, ZN => 
                           out_mask_10_port);
   U432 : AOI22_X1 port map( A1 => mask_3_10_port, A2 => n423, B1 => 
                           mask_2_10_port, B2 => n417, ZN => n167_port);
   U433 : AOI22_X1 port map( A1 => mask_1_10_port, A2 => n384, B1 => 
                           mask_0_10_port, B2 => n408, ZN => n166_port);
   U434 : NAND2_X1 port map( A1 => n164_port, A2 => n165_port, ZN => 
                           out_mask_11_port);
   U435 : AOI22_X1 port map( A1 => mask_3_11_port, A2 => n423, B1 => 
                           mask_2_11_port, B2 => n417, ZN => n165_port);
   U436 : AOI22_X1 port map( A1 => mask_1_11_port, A2 => n386, B1 => 
                           mask_0_11_port, B2 => n408, ZN => n164_port);
   U437 : NAND2_X1 port map( A1 => n162_port, A2 => n163_port, ZN => 
                           out_mask_12_port);
   U438 : AOI22_X1 port map( A1 => mask_3_12_port, A2 => n423, B1 => 
                           mask_2_12_port, B2 => n417, ZN => n163_port);
   U439 : AOI22_X1 port map( A1 => mask_1_12_port, A2 => n380, B1 => 
                           mask_0_12_port, B2 => n408, ZN => n162_port);
   U440 : NAND2_X1 port map( A1 => n152, A2 => n153, ZN => out_mask_17_port);
   U441 : AOI22_X1 port map( A1 => mask_3_17_port, A2 => n423, B1 => 
                           mask_2_17_port, B2 => n417, ZN => n153);
   U442 : AOI22_X1 port map( A1 => mask_1_17_port, A2 => n383, B1 => 
                           mask_0_17_port, B2 => n408, ZN => n152);
   U443 : NAND2_X1 port map( A1 => n110_port, A2 => n111_port, ZN => 
                           out_mask_36_port);
   U444 : AOI22_X1 port map( A1 => mask_3_36_port, A2 => n425, B1 => 
                           mask_2_36_port, B2 => n419, ZN => n111_port);
   U445 : AOI22_X1 port map( A1 => mask_1_36_port, A2 => n384, B1 => 
                           mask_0_36_port, B2 => n410, ZN => n110_port);
   U446 : NAND2_X1 port map( A1 => n158_port, A2 => n159_port, ZN => 
                           out_mask_14_port);
   U447 : AOI22_X1 port map( A1 => mask_3_14_port, A2 => n423, B1 => 
                           mask_2_14_port, B2 => n417, ZN => n159_port);
   U448 : AOI22_X1 port map( A1 => mask_1_14_port, A2 => n387, B1 => 
                           mask_0_14_port, B2 => n408, ZN => n158_port);
   U449 : NAND2_X1 port map( A1 => n160_port, A2 => n161_port, ZN => 
                           out_mask_13_port);
   U450 : AOI22_X1 port map( A1 => mask_3_13_port, A2 => n423, B1 => 
                           mask_2_13_port, B2 => n417, ZN => n161_port);
   U451 : AOI22_X1 port map( A1 => mask_1_13_port, A2 => n388, B1 => 
                           mask_0_13_port, B2 => n408, ZN => n160_port);
   U452 : AOI22_X1 port map( A1 => mask_3_1_port, A2 => n423, B1 => 
                           mask_2_1_port, B2 => n417, ZN => n147);
   U453 : AOI22_X1 port map( A1 => mask_1_1_port, A2 => n382, B1 => 
                           mask_0_1_port, B2 => n408, ZN => n146);
   U454 : AOI22_X1 port map( A1 => mask_1_39_port, A2 => n386, B1 => 
                           mask_0_39_port, B2 => n410, ZN => n104);
   U455 : AOI22_X1 port map( A1 => mask_1_0_port, A2 => n385, B1 => 
                           mask_0_0_port, B2 => n408, ZN => n168_port);
   U456 : AOI22_X1 port map( A1 => mask_3_39_port, A2 => n425, B1 => 
                           mask_2_39_port, B2 => n419, ZN => n105);
   U457 : NOR2_X1 port map( A1 => n534, A2 => conf(1), ZN => n239);
   U458 : AND2_X1 port map( A1 => conf(1), A2 => n534, ZN => n238);
   U459 : INV_X1 port map( A => conf(0), ZN => n534);
   U460 : NOR2_X1 port map( A1 => R(2), A2 => R(1), ZN => n298);
   U461 : NOR2_X1 port map( A1 => n301, A2 => R(1), ZN => n297);
   U462 : AOI22_X1 port map( A1 => n362, A2 => n5, B1 => n353, B2 => n306, ZN 
                           => n9);
   U463 : OAI221_X1 port map( B1 => out_mask_3_port, B2 => n372, C1 => 
                           out_mask_7_port, C2 => n375, A => n9, ZN => n13);
   U464 : OAI22_X1 port map( A1 => n376, A2 => n305, B1 => n373, B2 => n317, ZN
                           => n10);
   U465 : AOI221_X1 port map( B1 => out_mask_0_port, B2 => n357, C1 => 
                           out_mask_4_port, C2 => n353, A => n10, ZN => n11);
   U466 : OAI22_X1 port map( A1 => n13, A2 => n366, B1 => R(0), B2 => n11, ZN 
                           => N190);
   U467 : AOI22_X1 port map( A1 => n357, A2 => n317, B1 => n348, B2 => n305, ZN
                           => n12);
   U468 : OAI221_X1 port map( B1 => out_mask_4_port, B2 => n371, C1 => 
                           out_mask_8_port, C2 => n375, A => n12, ZN => n15);
   U469 : OAI22_X1 port map( A1 => n343, A2 => n13, B1 => n15, B2 => n370, ZN 
                           => N191);
   U470 : AOI22_X1 port map( A1 => n357, A2 => n308, B1 => n348, B2 => n304, ZN
                           => n14);
   U471 : OAI221_X1 port map( B1 => out_mask_5_port, B2 => n373, C1 => 
                           out_mask_9_port, C2 => n376, A => n14, ZN => n17);
   U472 : OAI22_X1 port map( A1 => n344, A2 => n15, B1 => n17, B2 => n370, ZN 
                           => N192);
   U473 : AOI22_X1 port map( A1 => n357, A2 => n307, B1 => n348, B2 => n303, ZN
                           => n16);
   U474 : OAI221_X1 port map( B1 => out_mask_6_port, B2 => n371, C1 => 
                           out_mask_10_port, C2 => n374, A => n16, ZN => n19);
   U475 : OAI22_X1 port map( A1 => R(0), A2 => n17, B1 => n19, B2 => n370, ZN 
                           => N193);
   U476 : AOI22_X1 port map( A1 => n357, A2 => n306, B1 => n348, B2 => n302, ZN
                           => n18);
   U477 : OAI221_X1 port map( B1 => out_mask_7_port, B2 => n371, C1 => 
                           out_mask_11_port, C2 => n374, A => n18, ZN => n21);
   U478 : OAI22_X1 port map( A1 => n343, A2 => n19, B1 => n21, B2 => n370, ZN 
                           => N194);
   U479 : AOI22_X1 port map( A1 => n357, A2 => n305, B1 => n348, B2 => n337, ZN
                           => n20);
   U480 : OAI221_X1 port map( B1 => out_mask_8_port, B2 => n373, C1 => 
                           out_mask_12_port, C2 => n376, A => n20, ZN => n23);
   U481 : OAI22_X1 port map( A1 => n343, A2 => n21, B1 => n23, B2 => n370, ZN 
                           => N195);
   U482 : AOI22_X1 port map( A1 => n357, A2 => n304, B1 => n348, B2 => n336, ZN
                           => n22);
   U483 : OAI221_X1 port map( B1 => out_mask_9_port, B2 => n373, C1 => 
                           out_mask_13_port, C2 => n376, A => n22, ZN => n25);
   U484 : OAI22_X1 port map( A1 => n344, A2 => n23, B1 => n25, B2 => n370, ZN 
                           => N196);
   U485 : AOI22_X1 port map( A1 => n357, A2 => n303, B1 => n348, B2 => n335, ZN
                           => n24);
   U486 : OAI221_X1 port map( B1 => out_mask_10_port, B2 => n372, C1 => 
                           out_mask_14_port, C2 => n376, A => n24, ZN => n27);
   U487 : OAI22_X1 port map( A1 => R(0), A2 => n25, B1 => n27, B2 => n370, ZN 
                           => N197);
   U488 : AOI22_X1 port map( A1 => n358, A2 => n302, B1 => n348, B2 => n334, ZN
                           => n26);
   U489 : OAI221_X1 port map( B1 => out_mask_11_port, B2 => n371, C1 => 
                           out_mask_15_port, C2 => n374, A => n26, ZN => n29);
   U490 : OAI22_X1 port map( A1 => n344, A2 => n27, B1 => n29, B2 => n370, ZN 
                           => N198);
   U491 : AOI22_X1 port map( A1 => n358, A2 => n337, B1 => n348, B2 => n333, ZN
                           => n28_port);
   U492 : OAI221_X1 port map( B1 => out_mask_12_port, B2 => n373, C1 => 
                           out_mask_16_port, C2 => n376, A => n28_port, ZN => 
                           n31);
   U493 : OAI22_X1 port map( A1 => n343, A2 => n29, B1 => n31, B2 => n370, ZN 
                           => N199);
   U494 : AOI22_X1 port map( A1 => n358, A2 => n336, B1 => n348, B2 => n332, ZN
                           => n30);
   U495 : OAI221_X1 port map( B1 => out_mask_13_port, B2 => n373, C1 => 
                           out_mask_17_port, C2 => n376, A => n30, ZN => n33);
   U496 : OAI22_X1 port map( A1 => n344, A2 => n31, B1 => n33, B2 => n369, ZN 
                           => N200);
   U497 : AOI22_X1 port map( A1 => n358, A2 => n335, B1 => n348, B2 => n331, ZN
                           => n32);
   U498 : OAI221_X1 port map( B1 => out_mask_14_port, B2 => n372, C1 => 
                           out_mask_18_port, C2 => n374, A => n32, ZN => 
                           n35_port);
   U499 : OAI22_X1 port map( A1 => R(0), A2 => n33, B1 => n35_port, B2 => n369,
                           ZN => N201);
   U500 : AOI22_X1 port map( A1 => n358, A2 => n334, B1 => n349, B2 => n330, ZN
                           => n34);
   U501 : OAI221_X1 port map( B1 => out_mask_15_port, B2 => n373, C1 => 
                           out_mask_19_port, C2 => n376, A => n34, ZN => 
                           n37_port);
   U502 : OAI22_X1 port map( A1 => n344, A2 => n35_port, B1 => n37_port, B2 => 
                           n369, ZN => N202);
   U503 : AOI22_X1 port map( A1 => n358, A2 => n333, B1 => n349, B2 => n329, ZN
                           => n36);
   U504 : OAI221_X1 port map( B1 => out_mask_16_port, B2 => n371, C1 => 
                           out_mask_20_port, C2 => n375, A => n36, ZN => 
                           n39_port);
   U505 : OAI22_X1 port map( A1 => R(0), A2 => n37_port, B1 => n39_port, B2 => 
                           n369, ZN => N203);
   U506 : AOI22_X1 port map( A1 => n358, A2 => n332, B1 => n349, B2 => n328, ZN
                           => n38_port);
   U507 : OAI221_X1 port map( B1 => out_mask_17_port, B2 => n373, C1 => 
                           out_mask_21_port, C2 => n375, A => n38_port, ZN => 
                           n41_port);
   U508 : OAI22_X1 port map( A1 => R(0), A2 => n39_port, B1 => n41_port, B2 => 
                           n369, ZN => N204);
   U509 : AOI22_X1 port map( A1 => n358, A2 => n331, B1 => n349, B2 => n327, ZN
                           => n40_port);
   U510 : OAI221_X1 port map( B1 => out_mask_18_port, B2 => n371, C1 => 
                           out_mask_22_port, C2 => n375, A => n40_port, ZN => 
                           n43_port);
   U511 : OAI22_X1 port map( A1 => n344, A2 => n41_port, B1 => n43_port, B2 => 
                           n368, ZN => N205);
   U512 : AOI22_X1 port map( A1 => n358, A2 => n330, B1 => n349, B2 => n326, ZN
                           => n42_port);
   U513 : OAI221_X1 port map( B1 => out_mask_19_port, B2 => n373, C1 => 
                           out_mask_23_port, C2 => n376, A => n42_port, ZN => 
                           n45_port);
   U514 : OAI22_X1 port map( A1 => n343, A2 => n43_port, B1 => n45_port, B2 => 
                           n369, ZN => N206);
   U515 : AOI22_X1 port map( A1 => n358, A2 => n329, B1 => n349, B2 => n325, ZN
                           => n44);
   U516 : OAI221_X1 port map( B1 => out_mask_20_port, B2 => n372, C1 => 
                           out_mask_24_port, C2 => n375, A => n44, ZN => 
                           n47_port);
   U517 : OAI22_X1 port map( A1 => n344, A2 => n45_port, B1 => n47_port, B2 => 
                           n369, ZN => N207);
   U518 : AOI22_X1 port map( A1 => n358, A2 => n328, B1 => n349, B2 => n324, ZN
                           => n46_port);
   U519 : OAI221_X1 port map( B1 => out_mask_21_port, B2 => n371, C1 => 
                           out_mask_25_port, C2 => n374, A => n46_port, ZN => 
                           n49_port);
   U520 : OAI22_X1 port map( A1 => R(0), A2 => n47_port, B1 => n49_port, B2 => 
                           n369, ZN => N208);
   U521 : AOI22_X1 port map( A1 => n359, A2 => n327, B1 => n349, B2 => n323, ZN
                           => n48_port);
   U522 : OAI221_X1 port map( B1 => out_mask_22_port, B2 => n372, C1 => 
                           out_mask_26_port, C2 => n375, A => n48_port, ZN => 
                           n51_port);
   U523 : OAI22_X1 port map( A1 => n343, A2 => n49_port, B1 => n51_port, B2 => 
                           n369, ZN => N209);
   U524 : AOI22_X1 port map( A1 => n359, A2 => n326, B1 => n349, B2 => n322, ZN
                           => n50_port);
   U525 : OAI221_X1 port map( B1 => out_mask_23_port, B2 => n372, C1 => 
                           out_mask_27_port, C2 => n375, A => n50_port, ZN => 
                           n53_port);
   U526 : OAI22_X1 port map( A1 => R(0), A2 => n51_port, B1 => n53_port, B2 => 
                           n369, ZN => N210);
   U527 : AOI22_X1 port map( A1 => n359, A2 => n325, B1 => n349, B2 => n321, ZN
                           => n52);
   U528 : OAI221_X1 port map( B1 => out_mask_24_port, B2 => n371, C1 => 
                           out_mask_28_port, C2 => n374, A => n52, ZN => 
                           n55_port);
   U529 : OAI22_X1 port map( A1 => n343, A2 => n53_port, B1 => n55_port, B2 => 
                           n369, ZN => N211);
   U530 : AOI22_X1 port map( A1 => n359, A2 => n324, B1 => n349, B2 => n320, ZN
                           => n54_port);
   U531 : OAI221_X1 port map( B1 => out_mask_25_port, B2 => n372, C1 => 
                           out_mask_29_port, C2 => n375, A => n54_port, ZN => 
                           n57_port);
   U532 : OAI22_X1 port map( A1 => n344, A2 => n55_port, B1 => n57_port, B2 => 
                           n368, ZN => N212);
   U533 : AOI22_X1 port map( A1 => n359, A2 => n323, B1 => n350, B2 => n319, ZN
                           => n56_port);
   U534 : OAI221_X1 port map( B1 => out_mask_26_port, B2 => n372, C1 => 
                           out_mask_30_port, C2 => n375, A => n56_port, ZN => 
                           n59_port);
   U535 : OAI22_X1 port map( A1 => R(0), A2 => n57_port, B1 => n59_port, B2 => 
                           n368, ZN => N213);
   U536 : AOI22_X1 port map( A1 => n359, A2 => n322, B1 => n350, B2 => n318, ZN
                           => n58_port);
   U537 : OAI221_X1 port map( B1 => out_mask_27_port, B2 => n372, C1 => 
                           out_mask_31_port, C2 => n375, A => n58_port, ZN => 
                           n61);
   U538 : OAI22_X1 port map( A1 => R(0), A2 => n59_port, B1 => n61, B2 => n368,
                           ZN => N214);
   U539 : AOI22_X1 port map( A1 => n359, A2 => n321, B1 => n350, B2 => n316, ZN
                           => n60_port);
   U540 : OAI221_X1 port map( B1 => out_mask_28_port, B2 => n372, C1 => 
                           out_mask_32_port, C2 => n374, A => n60_port, ZN => 
                           n63);
   U541 : OAI22_X1 port map( A1 => n343, A2 => n61, B1 => n63, B2 => n368, ZN 
                           => N215);
   U542 : AOI22_X1 port map( A1 => n359, A2 => n320, B1 => n350, B2 => n315, ZN
                           => n62);
   U543 : OAI221_X1 port map( B1 => out_mask_29_port, B2 => n371, C1 => 
                           out_mask_33_port, C2 => n374, A => n62, ZN => n65);
   U544 : OAI22_X1 port map( A1 => R(0), A2 => n63, B1 => n65, B2 => n368, ZN 
                           => N216);
   U545 : AOI22_X1 port map( A1 => n359, A2 => n319, B1 => n350, B2 => n314, ZN
                           => n64);
   U546 : OAI221_X1 port map( B1 => out_mask_30_port, B2 => n373, C1 => 
                           out_mask_34_port, C2 => n374, A => n64, ZN => n67);
   U547 : OAI22_X1 port map( A1 => R(0), A2 => n65, B1 => n67, B2 => n368, ZN 
                           => N217);
   U548 : AOI22_X1 port map( A1 => n359, A2 => n318, B1 => n350, B2 => n313, ZN
                           => n66);
   U549 : OAI221_X1 port map( B1 => out_mask_31_port, B2 => n372, C1 => 
                           out_mask_35_port, C2 => n375, A => n66, ZN => 
                           n69_port);
   U550 : OAI22_X1 port map( A1 => R(0), A2 => n67, B1 => n69_port, B2 => n368,
                           ZN => N218);
   U551 : AOI22_X1 port map( A1 => n359, A2 => n316, B1 => n350, B2 => n312, ZN
                           => n68_port);
   U552 : OAI221_X1 port map( B1 => out_mask_32_port, B2 => n371, C1 => 
                           out_mask_36_port, C2 => n374, A => n68_port, ZN => 
                           n71_port);
   U553 : OAI22_X1 port map( A1 => R(0), A2 => n69_port, B1 => n71_port, B2 => 
                           n368, ZN => N219);
   U554 : AOI22_X1 port map( A1 => n360, A2 => n315, B1 => n350, B2 => n311, ZN
                           => n70_port);
   U555 : OAI221_X1 port map( B1 => out_mask_33_port, B2 => n373, C1 => 
                           out_mask_37_port, C2 => n375, A => n70_port, ZN => 
                           n74_port);
   U556 : OAI22_X1 port map( A1 => R(0), A2 => n71_port, B1 => n74_port, B2 => 
                           n368, ZN => N220);
   U557 : OAI22_X1 port map( A1 => n375, A2 => n4, B1 => n372, B2 => n312, ZN 
                           => n72_port);
   U558 : AOI221_X1 port map( B1 => out_mask_32_port, B2 => n357, C1 => 
                           out_mask_36_port, C2 => n353, A => n72_port, ZN => 
                           n73_port);
   U559 : OAI22_X1 port map( A1 => R(0), A2 => n74_port, B1 => n370, B2 => 
                           n73_port, ZN => N221);
   U560 : AOI22_X1 port map( A1 => n360, A2 => n303, B1 => n350, B2 => n307, ZN
                           => n75_port);
   U561 : OAI221_X1 port map( B1 => out_mask_6_port, B2 => n372, C1 => 
                           out_mask_2_port, C2 => n375, A => n75_port, ZN => 
                           n79_port);
   U562 : OAI22_X1 port map( A1 => n374, A2 => n5, B1 => n371, B2 => n306, ZN 
                           => n76_port);
   U563 : AOI221_X1 port map( B1 => out_mask_7_port, B2 => n357, C1 => 
                           out_mask_3_port, C2 => n353, A => n76_port, ZN => 
                           n77_port);
   U564 : OAI22_X1 port map( A1 => R(0), A2 => n79_port, B1 => n370, B2 => 
                           n77_port, ZN => N158);
   U565 : AOI22_X1 port map( A1 => n360, A2 => n302, B1 => n351, B2 => n306, ZN
                           => n78_port);
   U566 : OAI221_X1 port map( B1 => out_mask_7_port, B2 => n371, C1 => 
                           out_mask_3_port, C2 => n374, A => n78_port, ZN => 
                           n81_port);
   U567 : OAI22_X1 port map( A1 => n79_port, A2 => n367, B1 => n344, B2 => 
                           n81_port, ZN => N159);
   U568 : AOI22_X1 port map( A1 => n360, A2 => n337, B1 => n351, B2 => n305, ZN
                           => n80_port);
   U569 : OAI221_X1 port map( B1 => out_mask_8_port, B2 => n372, C1 => 
                           out_mask_4_port, C2 => n375, A => n80_port, ZN => 
                           n83_port);
   U570 : OAI22_X1 port map( A1 => n81_port, A2 => n367, B1 => n344, B2 => 
                           n83_port, ZN => N160);
   U571 : AOI22_X1 port map( A1 => n360, A2 => n336, B1 => n351, B2 => n304, ZN
                           => n82_port);
   U572 : OAI221_X1 port map( B1 => out_mask_9_port, B2 => n373, C1 => 
                           out_mask_5_port, C2 => n374, A => n82_port, ZN => 
                           n85_port);
   U573 : OAI22_X1 port map( A1 => n83_port, A2 => n367, B1 => n344, B2 => 
                           n85_port, ZN => N161);
   U574 : AOI22_X1 port map( A1 => n360, A2 => n335, B1 => n351, B2 => n303, ZN
                           => n84);
   U575 : OAI221_X1 port map( B1 => out_mask_10_port, B2 => n372, C1 => 
                           out_mask_6_port, C2 => n376, A => n84, ZN => 
                           n89_port);
   U576 : OAI22_X1 port map( A1 => n85_port, A2 => n367, B1 => n344, B2 => 
                           n89_port, ZN => N162);
   U577 : AOI22_X1 port map( A1 => n360, A2 => n334, B1 => n351, B2 => n302, ZN
                           => n88_port);
   U578 : OAI221_X1 port map( B1 => out_mask_11_port, B2 => n371, C1 => 
                           out_mask_7_port, C2 => n376, A => n88_port, ZN => 
                           n218_port);
   U579 : OAI22_X1 port map( A1 => n89_port, A2 => n367, B1 => n344, B2 => 
                           n218_port, ZN => N163);
   U580 : AOI22_X1 port map( A1 => n360, A2 => n333, B1 => n351, B2 => n337, ZN
                           => n171_port);
   U581 : OAI221_X1 port map( B1 => out_mask_12_port, B2 => n372, C1 => 
                           out_mask_8_port, C2 => n376, A => n171_port, ZN => 
                           n249);
   U582 : OAI22_X1 port map( A1 => n218_port, A2 => n367, B1 => n344, B2 => 
                           n249, ZN => N164);
   U583 : AOI22_X1 port map( A1 => n360, A2 => n332, B1 => n351, B2 => n336, ZN
                           => n248);
   U584 : OAI221_X1 port map( B1 => out_mask_13_port, B2 => n372, C1 => 
                           out_mask_9_port, C2 => n375, A => n248, ZN => n251);
   U585 : OAI22_X1 port map( A1 => n249, A2 => n367, B1 => n344, B2 => n251, ZN
                           => N165);
   U586 : AOI22_X1 port map( A1 => n360, A2 => n331, B1 => n351, B2 => n335, ZN
                           => n250);
   U587 : OAI221_X1 port map( B1 => out_mask_14_port, B2 => n372, C1 => 
                           out_mask_10_port, C2 => n375, A => n250, ZN => n253)
                           ;
   U588 : OAI22_X1 port map( A1 => n251, A2 => n367, B1 => n344, B2 => n253, ZN
                           => N166);
   U589 : AOI22_X1 port map( A1 => n361, A2 => n330, B1 => n351, B2 => n334, ZN
                           => n252);
   U590 : OAI221_X1 port map( B1 => out_mask_15_port, B2 => n373, C1 => 
                           out_mask_11_port, C2 => n376, A => n252, ZN => n255)
                           ;
   U591 : OAI22_X1 port map( A1 => n253, A2 => n367, B1 => n344, B2 => n255, ZN
                           => N167);
   U592 : AOI22_X1 port map( A1 => n361, A2 => n329, B1 => n351, B2 => n333, ZN
                           => n254);
   U593 : OAI221_X1 port map( B1 => out_mask_16_port, B2 => n372, C1 => 
                           out_mask_12_port, C2 => n376, A => n254, ZN => n257)
                           ;
   U594 : OAI22_X1 port map( A1 => n255, A2 => n367, B1 => n344, B2 => n257, ZN
                           => N168);
   U595 : AOI22_X1 port map( A1 => n361, A2 => n328, B1 => n351, B2 => n332, ZN
                           => n256);
   U596 : OAI221_X1 port map( B1 => out_mask_17_port, B2 => n373, C1 => 
                           out_mask_13_port, C2 => n376, A => n256, ZN => n259)
                           ;
   U597 : OAI22_X1 port map( A1 => n257, A2 => n366, B1 => n344, B2 => n259, ZN
                           => N169);
   U598 : AOI22_X1 port map( A1 => n361, A2 => n327, B1 => n352, B2 => n331, ZN
                           => n258);
   U599 : OAI221_X1 port map( B1 => out_mask_18_port, B2 => n371, C1 => 
                           out_mask_14_port, C2 => n376, A => n258, ZN => n261)
                           ;
   U600 : OAI22_X1 port map( A1 => n259, A2 => n366, B1 => n343, B2 => n261, ZN
                           => N170);
   U601 : AOI22_X1 port map( A1 => n361, A2 => n326, B1 => n352, B2 => n330, ZN
                           => n260);
   U602 : OAI221_X1 port map( B1 => out_mask_19_port, B2 => n373, C1 => 
                           out_mask_15_port, C2 => n376, A => n260, ZN => n263)
                           ;
   U603 : OAI22_X1 port map( A1 => n261, A2 => n366, B1 => n343, B2 => n263, ZN
                           => N171);
   U604 : AOI22_X1 port map( A1 => n361, A2 => n325, B1 => n350, B2 => n329, ZN
                           => n262);
   U605 : OAI221_X1 port map( B1 => out_mask_20_port, B2 => n373, C1 => 
                           out_mask_16_port, C2 => n374, A => n262, ZN => n265)
                           ;
   U606 : OAI22_X1 port map( A1 => n263, A2 => n366, B1 => n343, B2 => n265, ZN
                           => N172);
   U607 : AOI22_X1 port map( A1 => n360, A2 => n324, B1 => n350, B2 => n328, ZN
                           => n264);
   U608 : OAI221_X1 port map( B1 => out_mask_21_port, B2 => n371, C1 => 
                           out_mask_17_port, C2 => n375, A => n264, ZN => n267)
                           ;
   U609 : OAI22_X1 port map( A1 => n265, A2 => n366, B1 => n343, B2 => n267, ZN
                           => N173);
   U610 : AOI22_X1 port map( A1 => n361, A2 => n323, B1 => n352, B2 => n327, ZN
                           => n266);
   U611 : OAI221_X1 port map( B1 => out_mask_22_port, B2 => n372, C1 => 
                           out_mask_18_port, C2 => n375, A => n266, ZN => n269)
                           ;
   U612 : OAI22_X1 port map( A1 => n267, A2 => n366, B1 => n343, B2 => n269, ZN
                           => N174);
   U613 : AOI22_X1 port map( A1 => n361, A2 => n322, B1 => n352, B2 => n326, ZN
                           => n268);
   U614 : OAI221_X1 port map( B1 => out_mask_23_port, B2 => n373, C1 => 
                           out_mask_19_port, C2 => n374, A => n268, ZN => n271)
                           ;
   U615 : OAI22_X1 port map( A1 => n269, A2 => n366, B1 => n343, B2 => n271, ZN
                           => N175);
   U616 : AOI22_X1 port map( A1 => n361, A2 => n321, B1 => n352, B2 => n325, ZN
                           => n270);
   U617 : OAI221_X1 port map( B1 => out_mask_24_port, B2 => n371, C1 => 
                           out_mask_20_port, C2 => n376, A => n270, ZN => n273)
                           ;
   U618 : OAI22_X1 port map( A1 => n271, A2 => n366, B1 => n343, B2 => n273, ZN
                           => N176);
   U619 : AOI22_X1 port map( A1 => n361, A2 => n320, B1 => n352, B2 => n324, ZN
                           => n272);
   U620 : OAI221_X1 port map( B1 => out_mask_25_port, B2 => n372, C1 => 
                           out_mask_21_port, C2 => n376, A => n272, ZN => n275)
                           ;
   U621 : OAI22_X1 port map( A1 => n273, A2 => n366, B1 => n343, B2 => n275, ZN
                           => N177);
   U622 : AOI22_X1 port map( A1 => n361, A2 => n319, B1 => n352, B2 => n323, ZN
                           => n274);
   U623 : OAI221_X1 port map( B1 => out_mask_26_port, B2 => n371, C1 => 
                           out_mask_22_port, C2 => n375, A => n274, ZN => n277)
                           ;
   U624 : OAI22_X1 port map( A1 => n275, A2 => n366, B1 => n343, B2 => n277, ZN
                           => N178);
   U625 : AOI22_X1 port map( A1 => n362, A2 => n318, B1 => n352, B2 => n322, ZN
                           => n276);
   U626 : OAI221_X1 port map( B1 => out_mask_27_port, B2 => n371, C1 => 
                           out_mask_23_port, C2 => n374, A => n276, ZN => n279)
                           ;
   U627 : OAI22_X1 port map( A1 => n277, A2 => n367, B1 => n343, B2 => n279, ZN
                           => N179);
   U628 : AOI22_X1 port map( A1 => n362, A2 => n316, B1 => n352, B2 => n321, ZN
                           => n278);
   U629 : OAI221_X1 port map( B1 => out_mask_28_port, B2 => n373, C1 => 
                           out_mask_24_port, C2 => n375, A => n278, ZN => n281)
                           ;
   U630 : OAI22_X1 port map( A1 => n279, A2 => n365, B1 => n343, B2 => n281, ZN
                           => N180);
   U631 : AOI22_X1 port map( A1 => n362, A2 => n315, B1 => n352, B2 => n320, ZN
                           => n280);
   U632 : OAI221_X1 port map( B1 => out_mask_29_port, B2 => n371, C1 => 
                           out_mask_25_port, C2 => n374, A => n280, ZN => n283)
                           ;
   U633 : OAI22_X1 port map( A1 => n281, A2 => n365, B1 => R(0), B2 => n283, ZN
                           => N181);
   U634 : AOI22_X1 port map( A1 => n362, A2 => n314, B1 => n353, B2 => n319, ZN
                           => n282);
   U635 : OAI221_X1 port map( B1 => out_mask_30_port, B2 => n371, C1 => 
                           out_mask_26_port, C2 => n374, A => n282, ZN => n285)
                           ;
   U636 : OAI22_X1 port map( A1 => n283, A2 => n365, B1 => n343, B2 => n285, ZN
                           => N182);
   U637 : AOI22_X1 port map( A1 => n362, A2 => n313, B1 => n353, B2 => n318, ZN
                           => n284);
   U638 : OAI221_X1 port map( B1 => out_mask_31_port, B2 => n371, C1 => 
                           out_mask_27_port, C2 => n374, A => n284, ZN => n287)
                           ;
   U639 : OAI22_X1 port map( A1 => n285, A2 => n365, B1 => n344, B2 => n287, ZN
                           => N183);
   U640 : AOI22_X1 port map( A1 => n362, A2 => n312, B1 => n353, B2 => n316, ZN
                           => n286);
   U641 : OAI221_X1 port map( B1 => out_mask_32_port, B2 => n372, C1 => 
                           out_mask_28_port, C2 => n374, A => n286, ZN => n289)
                           ;
   U642 : OAI22_X1 port map( A1 => n287, A2 => n365, B1 => R(0), B2 => n289, ZN
                           => N184);
   U643 : AOI22_X1 port map( A1 => n362, A2 => n311, B1 => n353, B2 => n315, ZN
                           => n288);
   U644 : OAI221_X1 port map( B1 => out_mask_33_port, B2 => n373, C1 => 
                           out_mask_29_port, C2 => n374, A => n288, ZN => n291)
                           ;
   U645 : OAI22_X1 port map( A1 => n289, A2 => n365, B1 => n343, B2 => n291, ZN
                           => N185);
   U646 : AOI22_X1 port map( A1 => n362, A2 => n310, B1 => n353, B2 => n314, ZN
                           => n290);
   U647 : OAI221_X1 port map( B1 => out_mask_34_port, B2 => n373, C1 => 
                           out_mask_30_port, C2 => n376, A => n290, ZN => n293)
                           ;
   U648 : OAI22_X1 port map( A1 => n291, A2 => n341, B1 => n344, B2 => n293, ZN
                           => N186);
   U649 : AOI22_X1 port map( A1 => n362, A2 => n309, B1 => n352, B2 => n313, ZN
                           => n292);
   U650 : OAI221_X1 port map( B1 => out_mask_35_port, B2 => n373, C1 => 
                           out_mask_31_port, C2 => n376, A => n292, ZN => n295)
                           ;
   U651 : OAI22_X1 port map( A1 => n293, A2 => n341, B1 => R(0), B2 => n295, ZN
                           => N187);
   U652 : AOI22_X1 port map( A1 => n362, A2 => n4, B1 => n353, B2 => n312, ZN 
                           => n294);
   U653 : OAI221_X1 port map( B1 => out_mask_36_port, B2 => n371, C1 => 
                           out_mask_32_port, C2 => n374, A => n294, ZN => n300)
                           ;
   U654 : OAI22_X1 port map( A1 => n295, A2 => n341, B1 => n343, B2 => n300, ZN
                           => N188);
   U655 : OAI22_X1 port map( A1 => n376, A2 => n313, B1 => n373, B2 => n309, ZN
                           => n296);
   U656 : AOI221_X1 port map( B1 => out_mask_39_port, B2 => n357, C1 => 
                           out_mask_35_port, C2 => n353, A => n296, ZN => n299)
                           ;
   U657 : OAI22_X1 port map( A1 => n300, A2 => n368, B1 => n344, B2 => n299, ZN
                           => N189);
   U658 : CLKBUF_X1 port map( A => n338, Z => n340);
   U659 : INV_X1 port map( A => n90_port, ZN => n377);
   U660 : INV_X1 port map( A => n90_port, ZN => n378);
   U661 : INV_X1 port map( A => n377, ZN => n379);
   U662 : INV_X1 port map( A => n377, ZN => n380);
   U663 : INV_X1 port map( A => n377, ZN => n381);
   U664 : INV_X1 port map( A => n378, ZN => n382);
   U665 : INV_X1 port map( A => n378, ZN => n383);
   U666 : INV_X1 port map( A => n378, ZN => n384);
   U667 : INV_X1 port map( A => n378, ZN => n385);
   U668 : INV_X1 port map( A => n378, ZN => n386);
   U669 : INV_X1 port map( A => n378, ZN => n387);
   U670 : INV_X1 port map( A => n377, ZN => n388);
   U671 : INV_X1 port map( A => n378, ZN => n389);
   U672 : NOR2_X1 port map( A1 => n532, A2 => R(4), ZN => n90_port);
   U673 : AOI22_X1 port map( A1 => N183, A2 => n400, B1 => N215, B2 => n393, ZN
                           => n185_port);
   U674 : AOI22_X1 port map( A1 => N175, A2 => n400, B1 => N207, B2 => n393, ZN
                           => n194_port);
   U675 : AOI22_X1 port map( A1 => N179, A2 => n400, B1 => N211, B2 => n393, ZN
                           => n189_port);
   U676 : AOI22_X1 port map( A1 => N180, A2 => n400, B1 => N212, B2 => n393, ZN
                           => n188_port);
   U677 : AOI22_X1 port map( A1 => N162, A2 => n399, B1 => N194, B2 => n403, ZN
                           => n176_port);
   U678 : AOI22_X1 port map( A1 => N161, A2 => n399, B1 => N193, B2 => n403, ZN
                           => n177_port);
   U679 : AOI22_X1 port map( A1 => N178, A2 => n400, B1 => N210, B2 => n393, ZN
                           => n190_port);
   U680 : AOI22_X1 port map( A1 => N176, A2 => n400, B1 => N208, B2 => n393, ZN
                           => n193_port);
   U681 : AOI22_X1 port map( A1 => N164, A2 => n399, B1 => N196, B2 => n403, ZN
                           => n174_port);
   U682 : AOI22_X1 port map( A1 => N163, A2 => n399, B1 => N195, B2 => n403, ZN
                           => n175_port);
   U683 : INV_X1 port map( A => n184_port, ZN => data_out(26));
   U684 : INV_X1 port map( A => n178_port, ZN => data_out(31));
   U685 : INV_X1 port map( A => n186_port, ZN => data_out(24));
   U686 : INV_X1 port map( A => n187_port, ZN => data_out(23));
   U687 : AOI22_X1 port map( A1 => N181, A2 => n400, B1 => N213, B2 => n395, ZN
                           => n187_port);
   U688 : INV_X1 port map( A => n201_port, ZN => data_out(10));
   U689 : INV_X1 port map( A => n180_port, ZN => data_out(2));
   U690 : AOI22_X1 port map( A1 => N160, A2 => n399, B1 => N192, B2 => n403, ZN
                           => n180_port);
   U691 : INV_X1 port map( A => n192_port, ZN => data_out(19));
   U692 : INV_X1 port map( A => n198_port, ZN => data_out(13));
   U693 : INV_X1 port map( A => n170_port, ZN => data_out(9));
   U694 : AOI22_X1 port map( A1 => N173, A2 => n399, B1 => N205, B2 => n395, ZN
                           => n196_port);
   U695 : INV_X1 port map( A => n182_port, ZN => data_out(28));
   U696 : INV_X1 port map( A => R(3), ZN => n532);
   U697 : INV_X1 port map( A => n173_port, ZN => data_out(7));
   U698 : AOI22_X1 port map( A1 => N185, A2 => n399, B1 => N217, B2 => n395, ZN
                           => n183_port);
   U699 : INV_X1 port map( A => n191_port, ZN => data_out(1));
   U700 : INV_X1 port map( A => n172_port, ZN => data_out(8));
   U701 : AOI22_X1 port map( A1 => N166, A2 => n399, B1 => N198, B2 => n403, ZN
                           => n172_port);
   U702 : INV_X1 port map( A => n202_port, ZN => data_out(0));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in std_logic
         ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end ADDER_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal C_internal, B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, 
      B_in_27_port, B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, 
      B_in_22_port, B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, 
      B_in_17_port, B_in_16_port, B_in_14_port, B_in_12_port, B_in_11_port, 
      B_in_10_port, B_in_9_port, B_in_8_port, B_in_7_port, B_in_6_port, 
      B_in_5_port, B_in_4_port, B_in_3_port, B_in_2_port, B_in_1_port, 
      B_in_0_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, carry_1_port, carry_0_port, n1, n2, n3, n4, 
      n5, n6, n7, n8 : std_logic;

begin
   
   U5 : XOR2_X1 port map( A => B(9), B => n8, Z => B_in_9_port);
   U6 : XOR2_X1 port map( A => B(8), B => n8, Z => B_in_8_port);
   U7 : XOR2_X1 port map( A => B(7), B => n5, Z => B_in_7_port);
   U8 : XOR2_X1 port map( A => B(6), B => n7, Z => B_in_6_port);
   U9 : XOR2_X1 port map( A => B(5), B => n8, Z => B_in_5_port);
   U10 : XOR2_X1 port map( A => B(4), B => n8, Z => B_in_4_port);
   U11 : XOR2_X1 port map( A => B(3), B => n5, Z => B_in_3_port);
   U12 : XOR2_X1 port map( A => B(31), B => n7, Z => B_in_31_port);
   U13 : XOR2_X1 port map( A => B(30), B => n8, Z => B_in_30_port);
   U14 : XOR2_X1 port map( A => B(2), B => n4, Z => B_in_2_port);
   U15 : XOR2_X1 port map( A => B(29), B => n4, Z => B_in_29_port);
   U16 : XOR2_X1 port map( A => B(28), B => n5, Z => B_in_28_port);
   U17 : XOR2_X1 port map( A => B(27), B => n5, Z => B_in_27_port);
   U18 : XOR2_X1 port map( A => B(26), B => n8, Z => B_in_26_port);
   U19 : XOR2_X1 port map( A => B(25), B => n4, Z => B_in_25_port);
   U20 : XOR2_X1 port map( A => B(24), B => n7, Z => B_in_24_port);
   U21 : XOR2_X1 port map( A => B(23), B => n4, Z => B_in_23_port);
   U22 : XOR2_X1 port map( A => B(22), B => n5, Z => B_in_22_port);
   U23 : XOR2_X1 port map( A => B(21), B => n7, Z => B_in_21_port);
   U24 : XOR2_X1 port map( A => B(20), B => n8, Z => B_in_20_port);
   U25 : XOR2_X1 port map( A => B(1), B => n5, Z => B_in_1_port);
   U26 : XOR2_X1 port map( A => B(19), B => n8, Z => B_in_19_port);
   U27 : XOR2_X1 port map( A => B(18), B => n7, Z => B_in_18_port);
   U28 : XOR2_X1 port map( A => B(17), B => n7, Z => B_in_17_port);
   U29 : XOR2_X1 port map( A => B(16), B => n4, Z => B_in_16_port);
   U31 : XOR2_X1 port map( A => B(14), B => n5, Z => B_in_14_port);
   U33 : XOR2_X1 port map( A => B(12), B => n4, Z => B_in_12_port);
   U34 : XOR2_X1 port map( A => B(11), B => n7, Z => B_in_11_port);
   U35 : XOR2_X1 port map( A => B(10), B => n5, Z => B_in_10_port);
   U1 : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           B_in_31_port, B(30) => B_in_30_port, B(29) => 
                           B_in_29_port, B(28) => B_in_28_port, B(27) => 
                           B_in_27_port, B(26) => B_in_26_port, B(25) => 
                           B_in_25_port, B(24) => B_in_24_port, B(23) => 
                           B_in_23_port, B(22) => B_in_22_port, B(21) => 
                           B_in_21_port, B(20) => B_in_20_port, B(19) => 
                           B_in_19_port, B(18) => B_in_18_port, B(17) => 
                           B_in_17_port, B(16) => B_in_16_port, B(15) => n2, 
                           B(14) => B_in_14_port, B(13) => n1, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Cin => C_internal, Co(8) => Cout, Co(7)
                           => carry_7_port, Co(6) => carry_6_port, Co(5) => 
                           carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   U2 : SUM_GEN_N_NBIT_PER_BLOCK4_NBLOCKS8_0 port map( A(31) => A(31), A(30) =>
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B_in_31_port, B(30) 
                           => B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => n2, B(14) => B_in_14_port, 
                           B(13) => n1, B(12) => B_in_12_port, B(11) => 
                           B_in_11_port, B(10) => B_in_10_port, B(9) => 
                           B_in_9_port, B(8) => B_in_8_port, B(7) => 
                           B_in_7_port, B(6) => B_in_6_port, B(5) => 
                           B_in_5_port, B(4) => B_in_4_port, B(3) => 
                           B_in_3_port, B(2) => B_in_2_port, B(1) => 
                           B_in_1_port, B(0) => n3, Ci(7) => carry_7_port, 
                           Ci(6) => carry_6_port, Ci(5) => carry_5_port, Ci(4) 
                           => carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           carry_0_port, S(31) => S(31), S(30) => S(30), S(29) 
                           => S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U4 : BUF_X1 port map( A => ADD_SUB, Z => n5);
   U30 : BUF_X1 port map( A => ADD_SUB, Z => n4);
   U32 : OR2_X1 port map( A1 => n7, A2 => Cin, ZN => C_internal);
   U36 : BUF_X1 port map( A => ADD_SUB, Z => n8);
   U37 : BUF_X1 port map( A => ADD_SUB, Z => n7);
   U38 : XOR2_X1 port map( A => B(13), B => n4, Z => n1);
   U39 : XOR2_X1 port map( A => B(15), B => n4, Z => n2);
   U40 : XOR2_X1 port map( A => B(0), B => n6, Z => n3);
   U41 : XOR2_X1 port map( A => B(0), B => n6, Z => B_in_0_port);
   U42 : CLKBUF_X1 port map( A => ADD_SUB, Z => n6);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_0;

architecture SYN_Behavioral of AND2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_NBIT32_NREG32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_NBIT32_NREG32;

architecture SYN_BEHAVIORAL of RF_NBIT32_NREG32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N193, N194, N195, N196, N197, 
      N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, 
      N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, 
      N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
      N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, 
      N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N259, 
      N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, 
      N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, 
      N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, 
      N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, 
      N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n1, n2, n3, n4, n5, n6, n7, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193_port, n194_port, n195_port, n196_port, n197_port, 
      n198_port, n199_port, n200_port, n201_port, n202_port, n203_port, 
      n204_port, n205_port, n206_port, n207_port, n208_port, n209_port, 
      n210_port, n211_port, n212_port, n213_port, n214_port, n215_port, 
      n216_port, n217_port, n218_port, n219_port, n220_port, n221_port, 
      n222_port, n223_port, n224_port, n225_port, n226_port, n227_port, 
      n228_port, n229_port, n230_port, n231_port, n232_port, n233_port, 
      n234_port, n235_port, n236_port, n237_port, n238_port, n239_port, 
      n240_port, n241_port, n242_port, n243_port, n244_port, n245_port, 
      n246_port, n247_port, n248_port, n249_port, n250_port, n251_port, 
      n252_port, n253_port, n254_port, n255_port, n256_port, n257, n258, 
      n259_port, n260_port, n261_port, n262_port, n263_port, n264_port, 
      n265_port, n266_port, n267_port, n268_port, n269_port, n270_port, 
      n271_port, n272_port, n273_port, n274_port, n275_port, n276_port, 
      n277_port, n278_port, n279_port, n280_port, n281_port, n282_port, 
      n283_port, n284_port, n285_port, n286_port, n287_port, n288_port, 
      n289_port, n290_port, n291_port, n292_port, n293_port, n294_port, 
      n295_port, n296_port, n297_port, n298_port, n299_port, n300_port, 
      n301_port, n302_port, n303_port, n304_port, n305_port, n306_port, 
      n307_port, n308_port, n309_port, n310_port, n311_port, n312_port, 
      n313_port, n314_port, n315_port, n316_port, n317_port, n318_port, 
      n319_port, n320_port, n321_port, n322_port, n323_port, n324_port, 
      n325_port, n326_port, n327_port, n328_port, n329_port, n330_port, 
      n331_port, n332_port, n333_port, n334_port, n335_port, n336_port, 
      n337_port, n338_port, n339_port, n340_port, n341_port, n342_port, 
      n343_port, n344_port, n345_port, n346_port, n347_port, n348_port, 
      n349_port, n350_port, n351_port, n352_port, n353_port, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, 
      n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, 
      n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, 
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, 
      n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, 
      n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
      n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, 
      n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
      n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
      n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
      n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
      n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
      n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
      n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
      n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, 
      n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, 
      n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, 
      n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
      n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, 
      n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
      n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, 
      n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, 
      n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, 
      n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, 
      n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, 
      n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
      n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, 
      n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, 
      n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, 
      n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, 
      n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, 
      n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, 
      n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, 
      n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
      n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, 
      n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, 
      n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, 
      n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
      n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
      n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, 
      n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, 
      n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, 
      n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
      n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, 
      n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, 
      n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, 
      n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, 
      n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
      n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
      n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, 
      n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
      n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, 
      n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, 
      n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, 
      n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
      n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
      n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, 
      n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, 
      n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
      n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, 
      n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
      n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859 : std_logic;

begin
   
   OUT1_reg_31_inst : DLH_X1 port map( G => CLK, D => N256, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => CLK, D => N255, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => CLK, D => N254, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => CLK, D => N253, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => CLK, D => N252, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => CLK, D => N251, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => CLK, D => N250, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => CLK, D => N249, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => CLK, D => N248, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => CLK, D => N247, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => CLK, D => N246, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => CLK, D => N245, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => CLK, D => N244, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => CLK, D => N243, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => CLK, D => N242, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => CLK, D => N241, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => CLK, D => N240, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => CLK, D => N239, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => CLK, D => N238, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => CLK, D => N237, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => CLK, D => N236, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => CLK, D => N235, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => CLK, D => N234, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => CLK, D => N233, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => CLK, D => N232, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => CLK, D => N231, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => CLK, D => N230, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => CLK, D => N229, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => CLK, D => N228, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => CLK, D => N227, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => CLK, D => N226, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => CLK, D => N225, Q => OUT1(0));
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => N353, D => n1774, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => N353, D => n1779, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => N353, D => n1784, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => N353, D => n1789, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => N353, D => n1794, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => N353, D => n1799, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N353, D => n1804, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => N353, D => n1809, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N353, D => n1814, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N353, D => n1819, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => N353, D => n1824, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => N353, D => n1829, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => N353, D => n1834, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => N353, D => n1839, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => N353, D => n1844, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => N352, D => n1774, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => N352, D => n1779, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => N352, D => n1784, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => N352, D => n1789, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => N352, D => n1794, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N352, D => n1799, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => N352, D => n1804, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N352, D => n1809, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N352, D => n1814, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N352, D => n1819, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => N352, D => n1824, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => N352, D => n1829, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => N352, D => n1834, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => N352, D => n1839, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => N352, D => n1844, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => N351, D => n1774, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => N351, D => n1779, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => N351, D => n1784, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => N351, D => n1789, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => N351, D => n1794, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N351, D => n1799, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => N351, D => n1804, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N351, D => n1809, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N351, D => n1814, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N351, D => n1819, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => N351, D => n1824, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => N351, D => n1829, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => N351, D => n1834, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => N351, D => n1839, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => N351, D => n1844, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => N350, D => n1774, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => N350, D => n1779, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => N350, D => n1784, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => N350, D => n1789, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => N350, D => n1794, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N350, D => n1799, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => N350, D => n1804, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N350, D => n1809, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N350, D => n1814, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N350, D => n1819, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => N350, D => n1824, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => N350, D => n1829, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => N350, D => n1834, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => N350, D => n1839, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => N350, D => n1844, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => N349, D => n1774, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => N349, D => n1779, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => N349, D => n1784, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => N349, D => n1789, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => N349, D => n1794, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N349, D => n1799, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => N349, D => n1804, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N349, D => n1809, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N349, D => n1814, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N349, D => n1819, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => N349, D => n1824, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => N349, D => n1829, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => N349, D => n1834, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => N349, D => n1839, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => N349, D => n1844, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => N348, D => n1774, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => N348, D => n1779, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => N348, D => n1784, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => N348, D => n1789, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => N348, D => n1794, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N348, D => n1799, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => N348, D => n1804, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N348, D => n1809, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N348, D => n1814, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N348, D => n1819, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => N348, D => n1824, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => N348, D => n1829, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => N348, D => n1834, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => N348, D => n1839, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => N348, D => n1844, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => N347, D => n1774, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => N347, D => n1779, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => N347, D => n1784, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => N347, D => n1789, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => N347, D => n1794, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N347, D => n1799, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => N347, D => n1804, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N347, D => n1809, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N347, D => n1814, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N347, D => n1819, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => N347, D => n1824, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => N347, D => n1829, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => N347, D => n1834, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => N347, D => n1839, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => N347, D => n1844, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => N346, D => n1779, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => N346, D => n1784, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => N346, D => n1789, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => N346, D => n1794, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => N346, D => n1799, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => N346, D => n1804, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N346, D => n1809, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N346, D => n1814, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N346, D => n1819, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => N346, D => n1824, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => N346, D => n1829, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => N346, D => n1834, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => N346, D => n1839, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N346, D => n1844, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => N345, D => n1829, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => N345, D => n1834, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => N345, D => n1839, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => N345, D => n1844, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => N344, D => n1829, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => N344, D => n1834, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => N344, D => n1839, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N344, D => n1844, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => N343, D => n1747, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => N343, D => n1750, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => N343, D => n1753, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => N343, D => n1756, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => N343, D => n1759, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => N343, D => n1762, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => N343, D => n1765, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => N343, D => n1768, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => N343, D => n1771, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => N343, D => n1775, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => N343, D => n1780, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => N343, D => n1785, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => N343, D => n1790, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => N343, D => n1795, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N343, D => n1800, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => N343, D => n1805, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N343, D => n1810, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N343, D => n1815, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N343, D => n1820, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => N343, D => n1825, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => N343, D => n1830, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => N343, D => n1835, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => N343, D => n1840, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => N343, D => n1845, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => N342, D => n1747, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => N342, D => n1750, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => N342, D => n1753, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => N342, D => n1756, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => N342, D => n1759, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => N342, D => n1762, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => N342, D => n1765, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => N342, D => n1768, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => N342, D => n1771, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => N342, D => n1775, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => N342, D => n1780, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => N342, D => n1785, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => N342, D => n1790, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => N342, D => n1795, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N342, D => n1800, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => N342, D => n1805, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N342, D => n1810, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N342, D => n1815, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N342, D => n1820, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => N342, D => n1825, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => N342, D => n1830, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => N342, D => n1835, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => N342, D => n1840, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => N342, D => n1845, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => N341, D => n1747, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => N341, D => n1750, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => N341, D => n1753, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => N341, D => n1756, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => N341, D => n1759, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => N341, D => n1762, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => N341, D => n1765, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => N341, D => n1768, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => N341, D => n1771, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => N341, D => n1775, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => N341, D => n1780, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => N341, D => n1785, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => N341, D => n1790, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => N341, D => n1795, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N341, D => n1800, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => N341, D => n1805, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N341, D => n1810, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N341, D => n1815, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N341, D => n1820, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => N341, D => n1825, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => N341, D => n1830, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => N341, D => n1835, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => N341, D => n1840, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => N341, D => n1845, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => N340, D => n1747, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => N340, D => n1750, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => N340, D => n1753, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => N340, D => n1756, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => N340, D => n1759, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => N340, D => n1762, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => N340, D => n1765, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => N340, D => n1768, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => N340, D => n1771, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => N340, D => n1775, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => N340, D => n1780, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => N340, D => n1785, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => N340, D => n1790, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => N340, D => n1795, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N340, D => n1800, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => N340, D => n1805, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N340, D => n1810, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N340, D => n1815, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N340, D => n1820, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => N340, D => n1825, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => N340, D => n1830, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => N340, D => n1835, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => N340, D => n1840, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => N340, D => n1845, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => N339, D => n1747, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => N339, D => n1750, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => N339, D => n1753, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => N339, D => n1756, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => N339, D => n1759, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => N339, D => n1762, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => N339, D => n1765, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => N339, D => n1768, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => N339, D => n1771, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => N339, D => n1775, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => N339, D => n1780, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => N339, D => n1785, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => N339, D => n1790, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => N339, D => n1795, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N339, D => n1800, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => N339, D => n1805, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N339, D => n1810, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N339, D => n1815, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N339, D => n1820, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => N339, D => n1825, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => N339, D => n1830, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => N339, D => n1835, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => N339, D => n1840, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => N339, D => n1845, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => N338, D => n1747, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => N338, D => n1750, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => N338, D => n1753, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => N338, D => n1756, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => N338, D => n1759, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => N338, D => n1762, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => N338, D => n1765, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => N338, D => n1768, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => N338, D => n1771, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => N338, D => n1775, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => N338, D => n1780, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => N338, D => n1785, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => N338, D => n1790, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => N338, D => n1795, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N338, D => n1800, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => N338, D => n1805, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N338, D => n1810, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N338, D => n1815, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N338, D => n1820, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => N338, D => n1825, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => N338, D => n1830, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => N338, D => n1835, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => N338, D => n1840, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => N338, D => n1845, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => N337, D => n1747, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => N337, D => n1750, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => N337, D => n1753, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => N337, D => n1756, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => N337, D => n1759, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => N337, D => n1762, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => N337, D => n1765, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => N337, D => n1768, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => N337, D => n1771, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => N337, D => n1775, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => N337, D => n1780, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => N337, D => n1785, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => N337, D => n1790, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => N337, D => n1795, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N337, D => n1800, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => N337, D => n1805, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N337, D => n1810, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N337, D => n1815, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N337, D => n1820, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => N337, D => n1825, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => N337, D => n1830, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => N337, D => n1835, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => N337, D => n1840, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => N337, D => n1845, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => N336, D => n1747, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => N336, D => n1750, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => N336, D => n1753, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => N336, D => n1756, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => N336, D => n1759, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => N336, D => n1762, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => N336, D => n1765, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => N336, D => n1768, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => N336, D => n1771, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => N336, D => n1775, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => N336, D => n1780, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => N336, D => n1785, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => N336, D => n1790, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => N336, D => n1795, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N336, D => n1800, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => N336, D => n1805, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N336, D => n1810, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N336, D => n1815, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N336, D => n1820, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => N336, D => n1825, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => N336, D => n1830, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => N336, D => n1835, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => N336, D => n1840, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => N336, D => n1845, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => N335, D => n1747, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => N335, D => n1750, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => N335, D => n1753, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => N335, D => n1756, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => N335, D => n1759, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => N335, D => n1762, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => N335, D => n1765, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => N335, D => n1768, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => N335, D => n1771, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => N335, D => n1775, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => N335, D => n1780, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => N335, D => n1785, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => N335, D => n1790, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => N335, D => n1795, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N335, D => n1800, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => N335, D => n1805, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N335, D => n1810, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N335, D => n1815, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N335, D => n1820, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => N335, D => n1825, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => N335, D => n1830, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => N335, D => n1835, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => N335, D => n1840, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => N335, D => n1845, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => N334, D => n1747, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => N334, D => n1750, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => N334, D => n1753, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => N334, D => n1756, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => N334, D => n1759, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => N334, D => n1762, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => N334, D => n1765, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => N334, D => n1768, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => N334, D => n1771, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => N334, D => n1775, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => N334, D => n1780, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => N334, D => n1785, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => N334, D => n1790, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => N334, D => n1795, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N334, D => n1800, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => N334, D => n1805, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N334, D => n1810, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N334, D => n1815, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N334, D => n1820, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => N334, D => n1825, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => N334, D => n1830, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => N334, D => n1835, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => N334, D => n1840, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => N334, D => n1845, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => N333, D => n1748, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => N333, D => n1751, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => N333, D => n1754, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => N333, D => n1757, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => N333, D => n1760, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => N333, D => n1763, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => N333, D => n1766, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => N333, D => n1769, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => N333, D => n1772, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => N333, D => n1776, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => N333, D => n1781, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => N333, D => n1786, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => N333, D => n1791, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => N333, D => n1796, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N333, D => n1801, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => N333, D => n1806, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N333, D => n1811, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N333, D => n1816, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N333, D => n1821, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => N333, D => n1826, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => N333, D => n1831, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => N333, D => n1836, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => N333, D => n1841, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => N333, D => n1846, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => N332, D => n1748, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => N332, D => n1751, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => N332, D => n1754, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => N332, D => n1757, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => N332, D => n1760, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => N332, D => n1763, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => N332, D => n1766, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => N332, D => n1769, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => N332, D => n1772, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => N332, D => n1776, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => N332, D => n1781, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => N332, D => n1786, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => N332, D => n1791, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => N332, D => n1796, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N332, D => n1801, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => N332, D => n1806, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N332, D => n1811, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N332, D => n1816, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N332, D => n1821, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => N332, D => n1826, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => N332, D => n1831, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => N332, D => n1836, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => N332, D => n1841, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => N332, D => n1846, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => N331, D => n1748, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => N331, D => n1751, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => N331, D => n1754, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => N331, D => n1757, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => N331, D => n1760, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => N331, D => n1763, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => N331, D => n1766, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => N331, D => n1769, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => N331, D => n1772, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => N331, D => n1776, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => N331, D => n1781, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => N331, D => n1786, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => N331, D => n1791, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => N331, D => n1796, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N331, D => n1801, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => N331, D => n1806, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N331, D => n1811, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N331, D => n1816, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N331, D => n1821, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => N331, D => n1826, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => N331, D => n1831, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => N331, D => n1836, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => N331, D => n1841, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => N331, D => n1846, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => N330, D => n1748, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => N330, D => n1751, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => N330, D => n1754, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => N330, D => n1757, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => N330, D => n1760, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => N330, D => n1763, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => N330, D => n1766, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => N330, D => n1769, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => N330, D => n1772, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => N330, D => n1776, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => N330, D => n1781, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => N330, D => n1786, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => N330, D => n1791, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N330, D => n1796, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N330, D => n1801, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => N330, D => n1806, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N330, D => n1811, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N330, D => n1816, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => N330, D => n1821, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => N330, D => n1826, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => N330, D => n1831, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => N330, D => n1836, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => N330, D => n1841, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => N330, D => n1846, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => N329, D => n1748, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => N329, D => n1751, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => N329, D => n1754, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => N329, D => n1757, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => N329, D => n1760, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => N329, D => n1763, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => N329, D => n1766, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => N329, D => n1769, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => N329, D => n1772, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => N329, D => n1776, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => N329, D => n1781, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => N329, D => n1786, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => N329, D => n1791, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => N329, D => n1796, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N329, D => n1801, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => N329, D => n1806, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N329, D => n1811, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N329, D => n1816, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N329, D => n1821, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => N329, D => n1826, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => N329, D => n1831, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => N329, D => n1836, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => N329, D => n1841, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => N329, D => n1846, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => N328, D => n1748, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => N328, D => n1751, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => N328, D => n1754, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => N328, D => n1757, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => N328, D => n1760, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => N328, D => n1763, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => N328, D => n1766, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => N328, D => n1769, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => N328, D => n1772, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => N328, D => n1776, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => N328, D => n1781, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => N328, D => n1786, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => N328, D => n1791, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => N328, D => n1796, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N328, D => n1801, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => N328, D => n1806, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N328, D => n1811, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N328, D => n1816, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N328, D => n1821, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => N328, D => n1826, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => N328, D => n1831, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => N328, D => n1836, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => N328, D => n1841, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => N328, D => n1846, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => N327, D => n1748, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => N327, D => n1751, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => N327, D => n1754, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => N327, D => n1757, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => N327, D => n1760, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => N327, D => n1763, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => N327, D => n1766, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => N327, D => n1769, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => N327, D => n1772, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => N327, D => n1776, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => N327, D => n1781, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => N327, D => n1786, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => N327, D => n1791, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => N327, D => n1796, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N327, D => n1801, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => N327, D => n1806, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N327, D => n1811, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N327, D => n1816, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N327, D => n1821, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => N327, D => n1826, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => N327, D => n1831, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => N327, D => n1836, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => N327, D => n1841, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => N327, D => n1846, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => N326, D => n1748, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => N326, D => n1751, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => N326, D => n1754, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => N326, D => n1757, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => N326, D => n1760, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => N326, D => n1763, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => N326, D => n1766, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => N326, D => n1769, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => N326, D => n1772, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => N326, D => n1776, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => N326, D => n1781, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => N326, D => n1786, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => N326, D => n1791, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => N326, D => n1796, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N326, D => n1801, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => N326, D => n1806, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N326, D => n1811, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N326, D => n1816, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N326, D => n1821, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => N326, D => n1826, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => N326, D => n1831, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => N326, D => n1836, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => N326, D => n1841, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => N326, D => n1846, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => N325, D => n1748, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => N325, D => n1751, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => N325, D => n1754, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => N325, D => n1757, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => N325, D => n1760, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => N325, D => n1763, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => N325, D => n1766, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => N325, D => n1769, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => N325, D => n1772, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => N325, D => n1776, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => N325, D => n1781, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => N325, D => n1786, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => N325, D => n1791, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => N325, D => n1796, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N325, D => n1801, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => N325, D => n1806, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N325, D => n1811, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N325, D => n1816, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N325, D => n1821, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => N325, D => n1826, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => N325, D => n1831, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => N325, D => n1836, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => N325, D => n1841, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => N325, D => n1846, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => N324, D => n1748, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => N324, D => n1751, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => N324, D => n1754, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => N324, D => n1757, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => N324, D => n1760, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => N324, D => n1763, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => N324, D => n1766, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => N324, D => n1769, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => N324, D => n1772, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => N324, D => n1776, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => N324, D => n1781, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => N324, D => n1786, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => N324, D => n1791, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => N324, D => n1796, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N324, D => n1801, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => N324, D => n1806, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N324, D => n1811, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N324, D => n1816, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N324, D => n1821, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => N324, D => n1826, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => N324, D => n1831, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => N324, D => n1836, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => N324, D => n1841, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => N324, D => n1846, Q => 
                           REGISTERS_30_0_port);
   OUT2_reg_31_inst : DLH_X1 port map( G => CLK, D => N322, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => CLK, D => N321, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => CLK, D => N320, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => CLK, D => N319, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => CLK, D => N318, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => CLK, D => N317, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => CLK, D => N316, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => CLK, D => N315, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => CLK, D => N314, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => CLK, D => N313, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => CLK, D => N312, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => CLK, D => N311, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => CLK, D => N310, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => CLK, D => N309, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => CLK, D => N308, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => CLK, D => N307, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => CLK, D => N306, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => CLK, D => N305, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => CLK, D => N304, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => CLK, D => N303, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => CLK, D => N302, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => CLK, D => N301, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => CLK, D => N300, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => CLK, D => N299, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => CLK, D => N298, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => CLK, D => N297, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => CLK, D => N296, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => CLK, D => N295, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => CLK, D => N294, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => CLK, D => N293, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => CLK, D => N292, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => CLK, D => N291, Q => OUT2(0));
   U35 : OAI21_X2 port map( B1 => n9, B2 => n10, A => n1746, ZN => N353);
   U36 : OAI21_X2 port map( B1 => n9, B2 => n11, A => n1746, ZN => N352);
   U37 : OAI21_X2 port map( B1 => n9, B2 => n12, A => n1746, ZN => N351);
   U38 : OAI21_X2 port map( B1 => n9, B2 => n13, A => n1746, ZN => N350);
   U39 : OAI21_X2 port map( B1 => n9, B2 => n14, A => n1746, ZN => N349);
   U40 : OAI21_X2 port map( B1 => n9, B2 => n15, A => n1746, ZN => N348);
   U41 : OAI21_X2 port map( B1 => n9, B2 => n16, A => n1746, ZN => N347);
   U42 : OAI21_X2 port map( B1 => n18, B2 => n19, A => n1746, ZN => N346);
   U43 : OAI21_X2 port map( B1 => n10, B2 => n18, A => n1746, ZN => N345);
   U44 : OAI21_X2 port map( B1 => n11, B2 => n18, A => n1745, ZN => N344);
   U45 : OAI21_X2 port map( B1 => n12, B2 => n18, A => n1745, ZN => N343);
   U46 : OAI21_X2 port map( B1 => n13, B2 => n18, A => n1745, ZN => N342);
   U47 : OAI21_X2 port map( B1 => n14, B2 => n18, A => n1745, ZN => N341);
   U48 : OAI21_X2 port map( B1 => n15, B2 => n18, A => n1745, ZN => N340);
   U49 : OAI21_X2 port map( B1 => n16, B2 => n18, A => n1745, ZN => N339);
   U50 : OAI21_X2 port map( B1 => n19, B2 => n20, A => n1745, ZN => N338);
   U51 : OAI21_X2 port map( B1 => n10, B2 => n20, A => n1745, ZN => N337);
   U52 : OAI21_X2 port map( B1 => n11, B2 => n20, A => n1745, ZN => N336);
   U53 : OAI21_X2 port map( B1 => n12, B2 => n20, A => n1745, ZN => N335);
   U54 : OAI21_X2 port map( B1 => n13, B2 => n20, A => n1745, ZN => N334);
   U55 : OAI21_X2 port map( B1 => n14, B2 => n20, A => n1744, ZN => N333);
   U56 : OAI21_X2 port map( B1 => n15, B2 => n20, A => n1744, ZN => N332);
   U57 : OAI21_X2 port map( B1 => n16, B2 => n20, A => n1744, ZN => N331);
   U58 : OAI21_X2 port map( B1 => n19, B2 => n21, A => n1744, ZN => N330);
   U59 : OAI21_X2 port map( B1 => n10, B2 => n21, A => n1744, ZN => N329);
   U60 : OAI21_X2 port map( B1 => n11, B2 => n21, A => n1744, ZN => N328);
   U61 : OAI21_X2 port map( B1 => n12, B2 => n21, A => n1744, ZN => N327);
   U62 : OAI21_X2 port map( B1 => n13, B2 => n21, A => n1744, ZN => N326);
   U63 : OAI21_X2 port map( B1 => n14, B2 => n21, A => n1744, ZN => N325);
   U64 : OAI21_X2 port map( B1 => n15, B2 => n21, A => n1744, ZN => N324);
   U65 : OAI21_X2 port map( B1 => n16, B2 => n21, A => n1744, ZN => N323);
   U177 : NAND3_X1 port map( A1 => n1855, A2 => n1854, A3 => n17, ZN => n9);
   U178 : NAND3_X1 port map( A1 => n17, A2 => n1854, A3 => ADD_WR(3), ZN => n18
                           );
   U179 : NAND3_X1 port map( A1 => n17, A2 => n1855, A3 => ADD_WR(4), ZN => n20
                           );
   U180 : NAND3_X1 port map( A1 => n1857, A2 => n1856, A3 => n1858, ZN => n19);
   U181 : NAND3_X1 port map( A1 => n1857, A2 => n1856, A3 => ADD_WR(0), ZN => 
                           n10);
   U182 : NAND3_X1 port map( A1 => n1858, A2 => n1856, A3 => ADD_WR(1), ZN => 
                           n11);
   U183 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1856, A3 => ADD_WR(1), ZN 
                           => n12);
   U184 : NAND3_X1 port map( A1 => n1858, A2 => n1857, A3 => ADD_WR(2), ZN => 
                           n13);
   U185 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1857, A3 => ADD_WR(2), ZN 
                           => n14);
   U186 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n1858, A3 => ADD_WR(2), ZN 
                           => n15);
   U187 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n17, A3 => ADD_WR(4), ZN =>
                           n21);
   U188 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n16);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => N323, D => n56, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => N323, D => n55, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => N323, D => n54, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => N323, D => n53, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => N323, D => n52, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => N323, D => n51, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => N323, D => n50, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => N323, D => n49, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => N323, D => n48, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => N323, D => n47, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => N323, D => n46, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => N323, D => n45, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => N323, D => n44, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => N323, D => n43, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => N323, D => n42, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => N323, D => n41, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => N323, D => n40, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => N323, D => n38, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => N323, D => n37, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => N323, D => n36, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => N323, D => n35, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => N323, D => n34, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N323, D => n33, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => N323, D => n32, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N323, D => n31, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N323, D => n30, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N323, D => n29, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => N323, D => n28, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => N323, D => n7, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => N323, D => n6, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => N323, D => n39, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => N344, D => n56, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => N345, D => n56, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => N346, D => n56, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => N347, D => n56, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => N348, D => n56, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => N349, D => n56, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => N350, D => n56, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => N351, D => n56, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => N352, D => n56, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => N353, D => n56, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => N344, D => n55, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => N344, D => n54, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => N344, D => n53, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => N344, D => n52, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => N344, D => n51, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => N344, D => n50, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => N345, D => n55, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => N345, D => n54, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => N345, D => n53, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => N345, D => n52, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => N345, D => n51, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => N345, D => n50, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => N346, D => n55, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => N346, D => n54, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => N346, D => n53, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => N346, D => n52, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => N346, D => n51, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => N346, D => n50, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => N347, D => n55, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => N347, D => n54, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => N347, D => n53, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => N347, D => n52, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => N347, D => n51, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => N347, D => n50, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => N348, D => n55, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => N348, D => n54, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => N348, D => n53, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => N348, D => n52, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => N348, D => n51, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => N348, D => n50, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => N349, D => n55, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => N349, D => n54, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => N349, D => n53, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => N349, D => n52, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => N349, D => n51, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => N349, D => n50, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => N350, D => n55, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => N350, D => n54, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => N350, D => n53, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => N350, D => n52, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => N350, D => n51, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => N350, D => n50, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => N351, D => n55, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => N351, D => n54, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => N351, D => n53, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => N351, D => n52, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => N351, D => n51, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => N351, D => n50, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => N352, D => n55, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => N352, D => n54, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => N352, D => n53, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => N352, D => n52, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => N352, D => n51, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => N352, D => n50, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => N353, D => n55, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => N353, D => n54, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => N353, D => n53, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => N353, D => n52, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => N353, D => n51, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => N353, D => n50, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => N344, D => n49, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => N345, D => n49, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => N346, D => n49, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => N347, D => n49, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => N348, D => n49, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => N349, D => n49, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => N350, D => n49, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => N351, D => n49, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => N352, D => n49, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => N353, D => n49, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => N323, D => n1, Q => 
                           REGISTERS_31_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => N324, D => n56, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => N325, D => n56, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => N326, D => n56, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => N327, D => n56, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => N328, D => n56, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => N329, D => n56, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => N330, D => n56, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => N331, D => n56, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => N332, D => n56, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => N333, D => n56, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => N334, D => n56, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => N335, D => n56, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => N336, D => n56, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => N337, D => n56, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => N338, D => n56, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => N339, D => n56, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => N340, D => n56, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => N341, D => n56, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => N342, D => n56, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => N343, D => n56, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => N324, D => n55, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => N324, D => n54, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => N324, D => n53, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => N324, D => n52, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => N324, D => n51, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => N324, D => n50, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => N325, D => n55, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => N325, D => n54, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => N325, D => n53, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => N325, D => n52, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => N325, D => n51, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => N325, D => n50, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => N326, D => n55, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => N326, D => n54, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => N326, D => n53, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => N326, D => n52, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => N326, D => n51, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => N326, D => n50, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => N327, D => n55, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => N327, D => n54, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => N327, D => n53, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => N327, D => n52, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => N327, D => n51, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => N327, D => n50, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => N328, D => n55, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => N328, D => n54, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => N328, D => n53, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => N328, D => n52, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => N328, D => n51, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => N328, D => n50, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => N329, D => n55, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => N329, D => n54, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => N329, D => n53, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => N329, D => n52, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => N329, D => n51, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => N329, D => n50, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => N330, D => n55, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => N330, D => n54, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => N330, D => n53, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => N330, D => n52, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => N330, D => n51, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => N330, D => n50, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => N331, D => n55, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => N331, D => n54, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => N331, D => n53, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => N331, D => n52, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => N331, D => n51, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => N331, D => n50, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => N332, D => n55, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => N332, D => n54, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => N332, D => n53, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => N332, D => n52, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => N332, D => n51, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => N332, D => n50, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => N333, D => n55, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => N333, D => n54, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => N333, D => n53, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => N333, D => n52, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => N333, D => n51, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => N333, D => n50, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => N334, D => n55, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => N334, D => n54, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => N334, D => n53, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => N334, D => n52, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => N334, D => n51, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => N334, D => n50, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => N335, D => n55, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => N335, D => n54, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => N335, D => n53, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => N335, D => n52, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => N335, D => n51, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => N335, D => n50, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => N336, D => n55, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => N336, D => n54, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => N336, D => n53, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => N336, D => n52, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => N336, D => n51, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => N336, D => n50, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => N337, D => n55, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => N337, D => n54, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => N337, D => n53, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => N337, D => n52, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => N337, D => n51, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => N337, D => n50, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => N338, D => n55, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => N338, D => n54, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => N338, D => n53, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => N338, D => n52, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => N338, D => n51, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => N338, D => n50, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => N339, D => n55, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => N339, D => n54, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => N339, D => n53, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => N339, D => n52, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => N339, D => n51, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => N339, D => n50, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => N340, D => n55, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => N340, D => n54, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => N340, D => n53, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => N340, D => n52, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => N340, D => n51, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => N340, D => n50, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => N341, D => n55, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => N341, D => n54, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => N341, D => n53, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => N341, D => n52, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => N341, D => n51, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => N341, D => n50, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => N342, D => n55, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => N342, D => n54, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => N342, D => n53, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => N342, D => n52, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => N342, D => n51, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => N342, D => n50, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => N343, D => n55, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => N343, D => n54, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => N343, D => n53, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => N343, D => n52, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => N343, D => n51, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => N343, D => n50, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => N324, D => n49, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => N325, D => n49, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => N326, D => n49, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => N327, D => n49, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => N328, D => n49, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => N329, D => n49, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => N330, D => n49, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => N331, D => n49, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => N332, D => n49, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => N333, D => n49, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => N334, D => n49, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => N335, D => n49, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => N336, D => n49, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => N337, D => n49, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => N338, D => n49, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => N339, D => n49, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => N340, D => n49, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => N341, D => n49, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => N342, D => n49, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => N343, D => n49, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => N344, D => n48, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => N344, D => n47, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => N344, D => n46, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => N344, D => n45, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => N344, D => n44, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => N344, D => n43, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => N344, D => n42, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => N344, D => n41, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => N344, D => n40, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => N345, D => n48, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => N345, D => n47, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => N345, D => n46, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => N345, D => n45, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => N345, D => n44, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => N345, D => n43, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => N345, D => n42, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => N345, D => n41, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => N345, D => n40, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => N346, D => n48, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => N346, D => n47, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => N346, D => n46, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => N346, D => n45, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => N346, D => n44, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => N346, D => n43, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => N346, D => n42, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => N346, D => n41, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => N346, D => n40, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => N347, D => n48, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => N347, D => n47, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => N347, D => n46, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => N347, D => n45, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => N347, D => n44, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => N347, D => n43, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => N347, D => n42, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => N347, D => n41, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => N347, D => n40, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => N348, D => n48, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => N348, D => n47, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => N348, D => n46, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => N348, D => n45, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => N348, D => n44, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => N348, D => n43, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => N348, D => n42, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => N348, D => n41, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => N348, D => n40, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => N349, D => n48, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => N349, D => n47, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => N349, D => n46, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => N349, D => n45, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => N349, D => n44, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => N349, D => n43, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => N349, D => n42, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => N349, D => n41, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => N349, D => n40, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => N350, D => n48, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => N350, D => n47, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => N350, D => n46, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => N350, D => n45, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => N350, D => n44, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => N350, D => n43, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => N350, D => n42, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => N350, D => n41, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => N350, D => n40, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => N351, D => n48, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => N351, D => n47, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => N351, D => n46, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => N351, D => n45, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => N351, D => n44, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => N351, D => n43, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => N351, D => n42, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => N351, D => n41, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => N351, D => n40, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => N352, D => n48, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => N352, D => n47, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => N352, D => n46, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => N352, D => n45, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => N352, D => n44, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => N352, D => n43, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => N352, D => n42, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => N352, D => n41, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => N352, D => n40, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => N353, D => n48, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => N353, D => n47, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => N353, D => n46, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => N353, D => n45, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N353, D => n44, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => N353, D => n43, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => N353, D => n42, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => N353, D => n41, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => N353, D => n40, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => N344, D => n38, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => N344, D => n37, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => N344, D => n36, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => N344, D => n35, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N344, D => n34, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => N344, D => n33, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N344, D => n32, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => N344, D => n31, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => N344, D => n30, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N344, D => n29, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => N344, D => n28, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => N345, D => n38, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => N345, D => n37, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => N345, D => n36, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => N345, D => n35, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => N345, D => n34, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N345, D => n33, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => N345, D => n32, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N345, D => n31, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N345, D => n30, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N345, D => n29, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => N345, D => n28, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => N346, D => n38, Q => 
                           REGISTERS_8_21_port);
   U3 : AND2_X1 port map( A1 => DATAIN(0), A2 => n1850, ZN => n1);
   U4 : AND2_X1 port map( A1 => n900, A2 => n1582, ZN => n2);
   U5 : AND2_X1 port map( A1 => n65, A2 => n747, ZN => n3);
   U6 : AND2_X1 port map( A1 => n66, A2 => n747, ZN => n4);
   U7 : AND2_X1 port map( A1 => n901, A2 => n1582, ZN => n5);
   U8 : BUF_X1 port map( A => n1849, Z => n1853);
   U9 : BUF_X1 port map( A => n1677, Z => n1678);
   U10 : BUF_X1 port map( A => n1659, Z => n1660);
   U11 : BUF_X1 port map( A => n1677, Z => n1679);
   U12 : BUF_X1 port map( A => n1659, Z => n1661);
   U13 : BUF_X1 port map( A => n1677, Z => n1680);
   U14 : BUF_X1 port map( A => n1659, Z => n1662);
   U15 : BUF_X1 port map( A => n842, Z => n843);
   U16 : BUF_X1 port map( A => n824, Z => n825);
   U17 : BUF_X1 port map( A => n842, Z => n844);
   U18 : BUF_X1 port map( A => n824, Z => n826);
   U19 : BUF_X1 port map( A => n842, Z => n845);
   U20 : BUF_X1 port map( A => n824, Z => n827);
   U21 : BUF_X1 port map( A => n6, Z => n1837);
   U22 : BUF_X1 port map( A => n7, Z => n1832);
   U23 : BUF_X1 port map( A => n28, Z => n1827);
   U24 : BUF_X1 port map( A => n29, Z => n1822);
   U25 : BUF_X1 port map( A => n30, Z => n1817);
   U26 : BUF_X1 port map( A => n31, Z => n1812);
   U27 : BUF_X1 port map( A => n32, Z => n1807);
   U28 : BUF_X1 port map( A => n33, Z => n1802);
   U29 : BUF_X1 port map( A => n34, Z => n1797);
   U30 : BUF_X1 port map( A => n35, Z => n1792);
   U31 : BUF_X1 port map( A => n36, Z => n1787);
   U32 : BUF_X1 port map( A => n37, Z => n1782);
   U33 : BUF_X1 port map( A => n38, Z => n1777);
   U34 : BUF_X1 port map( A => n39, Z => n1842);
   U66 : BUF_X1 port map( A => n1, Z => n1847);
   U67 : BUF_X1 port map( A => n40, Z => n1773);
   U68 : BUF_X1 port map( A => n41, Z => n1770);
   U69 : BUF_X1 port map( A => n42, Z => n1767);
   U70 : BUF_X1 port map( A => n43, Z => n1764);
   U71 : BUF_X1 port map( A => n44, Z => n1761);
   U72 : BUF_X1 port map( A => n45, Z => n1758);
   U73 : BUF_X1 port map( A => n46, Z => n1755);
   U74 : BUF_X1 port map( A => n47, Z => n1752);
   U75 : BUF_X1 port map( A => n48, Z => n1749);
   U76 : BUF_X1 port map( A => n2, Z => n1677);
   U77 : BUF_X1 port map( A => n5, Z => n1659);
   U78 : BUF_X1 port map( A => n3, Z => n842);
   U79 : BUF_X1 port map( A => n4, Z => n824);
   U80 : BUF_X1 port map( A => n1641, Z => n1642);
   U81 : BUF_X1 port map( A => n1623, Z => n1624);
   U82 : BUF_X1 port map( A => n1605, Z => n1606);
   U83 : BUF_X1 port map( A => n1587, Z => n1588);
   U84 : BUF_X1 port map( A => n1641, Z => n1643);
   U85 : BUF_X1 port map( A => n1623, Z => n1625);
   U86 : BUF_X1 port map( A => n1605, Z => n1607);
   U87 : BUF_X1 port map( A => n1587, Z => n1589);
   U88 : BUF_X1 port map( A => n1641, Z => n1644);
   U89 : BUF_X1 port map( A => n1623, Z => n1626);
   U90 : BUF_X1 port map( A => n1605, Z => n1608);
   U91 : BUF_X1 port map( A => n1587, Z => n1590);
   U92 : BUF_X1 port map( A => n806, Z => n807);
   U93 : BUF_X1 port map( A => n788, Z => n789);
   U94 : BUF_X1 port map( A => n770, Z => n771);
   U95 : BUF_X1 port map( A => n752, Z => n753);
   U96 : BUF_X1 port map( A => n806, Z => n808);
   U97 : BUF_X1 port map( A => n788, Z => n790);
   U98 : BUF_X1 port map( A => n770, Z => n772);
   U99 : BUF_X1 port map( A => n752, Z => n754);
   U100 : BUF_X1 port map( A => n806, Z => n809);
   U101 : BUF_X1 port map( A => n788, Z => n791);
   U102 : BUF_X1 port map( A => n770, Z => n773);
   U103 : BUF_X1 port map( A => n752, Z => n755);
   U104 : BUF_X1 port map( A => n1706, Z => n1707);
   U105 : BUF_X1 port map( A => n1706, Z => n1708);
   U106 : BUF_X1 port map( A => n1706, Z => n1709);
   U107 : BUF_X1 port map( A => n871, Z => n872);
   U108 : BUF_X1 port map( A => n871, Z => n873);
   U109 : BUF_X1 port map( A => n871, Z => n874);
   U110 : BUF_X1 port map( A => n1694, Z => n1697);
   U111 : BUF_X1 port map( A => n1694, Z => n1696);
   U112 : BUF_X1 port map( A => n859, Z => n862);
   U113 : BUF_X1 port map( A => n859, Z => n861);
   U114 : BUF_X1 port map( A => n1676, Z => n1681);
   U115 : BUF_X1 port map( A => n1658, Z => n1663);
   U116 : BUF_X1 port map( A => n841, Z => n846);
   U117 : BUF_X1 port map( A => n823, Z => n828);
   U118 : AND2_X1 port map( A1 => DATAIN(2), A2 => n1850, ZN => n6);
   U119 : AND2_X1 port map( A1 => DATAIN(10), A2 => n1850, ZN => n7);
   U120 : AND2_X1 port map( A1 => DATAIN(11), A2 => n1851, ZN => n28);
   U121 : AND2_X1 port map( A1 => DATAIN(12), A2 => n1851, ZN => n29);
   U122 : AND2_X1 port map( A1 => DATAIN(13), A2 => n1851, ZN => n30);
   U123 : AND2_X1 port map( A1 => DATAIN(14), A2 => n1851, ZN => n31);
   U124 : AND2_X1 port map( A1 => DATAIN(15), A2 => n1851, ZN => n32);
   U125 : AND2_X1 port map( A1 => DATAIN(16), A2 => n1851, ZN => n33);
   U126 : AND2_X1 port map( A1 => DATAIN(17), A2 => n1851, ZN => n34);
   U127 : AND2_X1 port map( A1 => DATAIN(18), A2 => n1851, ZN => n35);
   U128 : AND2_X1 port map( A1 => DATAIN(19), A2 => n1851, ZN => n36);
   U129 : AND2_X1 port map( A1 => DATAIN(20), A2 => n1851, ZN => n37);
   U130 : AND2_X1 port map( A1 => DATAIN(21), A2 => n1851, ZN => n38);
   U131 : AND2_X1 port map( A1 => DATAIN(1), A2 => n1850, ZN => n39);
   U132 : AND2_X1 port map( A1 => DATAIN(22), A2 => n1852, ZN => n40);
   U133 : AND2_X1 port map( A1 => DATAIN(23), A2 => n1852, ZN => n41);
   U134 : AND2_X1 port map( A1 => DATAIN(24), A2 => n1852, ZN => n42);
   U135 : AND2_X1 port map( A1 => DATAIN(25), A2 => n1852, ZN => n43);
   U136 : AND2_X1 port map( A1 => DATAIN(26), A2 => n1852, ZN => n44);
   U137 : AND2_X1 port map( A1 => DATAIN(27), A2 => n1852, ZN => n45);
   U138 : AND2_X1 port map( A1 => DATAIN(28), A2 => n1852, ZN => n46);
   U139 : AND2_X1 port map( A1 => DATAIN(29), A2 => n1852, ZN => n47);
   U140 : AND2_X1 port map( A1 => DATAIN(30), A2 => n1852, ZN => n48);
   U141 : AND2_X1 port map( A1 => DATAIN(9), A2 => n1850, ZN => n49);
   U142 : AND2_X1 port map( A1 => DATAIN(3), A2 => n1850, ZN => n50);
   U143 : AND2_X1 port map( A1 => DATAIN(4), A2 => n1850, ZN => n51);
   U144 : AND2_X1 port map( A1 => DATAIN(5), A2 => n1850, ZN => n52);
   U145 : AND2_X1 port map( A1 => DATAIN(6), A2 => n1850, ZN => n53);
   U146 : AND2_X1 port map( A1 => DATAIN(7), A2 => n1850, ZN => n54);
   U147 : AND2_X1 port map( A1 => DATAIN(8), A2 => n1850, ZN => n55);
   U148 : AND2_X1 port map( A1 => DATAIN(31), A2 => n1852, ZN => n56);
   U149 : BUF_X1 port map( A => n59, Z => n1641);
   U150 : BUF_X1 port map( A => n60, Z => n1623);
   U151 : BUF_X1 port map( A => n61, Z => n1605);
   U152 : BUF_X1 port map( A => n57, Z => n1587);
   U153 : BUF_X1 port map( A => n62, Z => n806);
   U154 : BUF_X1 port map( A => n63, Z => n788);
   U155 : BUF_X1 port map( A => n64, Z => n770);
   U156 : BUF_X1 port map( A => n58, Z => n752);
   U157 : BUF_X1 port map( A => n1568, Z => n1706);
   U158 : BUF_X1 port map( A => n1567, Z => n1694);
   U159 : BUF_X1 port map( A => n733, Z => n871);
   U160 : BUF_X1 port map( A => n732, Z => n859);
   U161 : BUF_X1 port map( A => n8, Z => n1743);
   U162 : BUF_X1 port map( A => n1640, Z => n1645);
   U163 : BUF_X1 port map( A => n1622, Z => n1627);
   U164 : BUF_X1 port map( A => n1604, Z => n1609);
   U165 : BUF_X1 port map( A => n1586, Z => n1591);
   U166 : BUF_X1 port map( A => n805, Z => n810);
   U167 : BUF_X1 port map( A => n787, Z => n792);
   U168 : BUF_X1 port map( A => n769, Z => n774);
   U169 : BUF_X1 port map( A => n751, Z => n756);
   U170 : BUF_X1 port map( A => n743, Z => n892);
   U171 : BUF_X1 port map( A => n745, Z => n896);
   U172 : BUF_X1 port map( A => n741, Z => n888);
   U173 : BUF_X1 port map( A => n739, Z => n884);
   U174 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n901, ZN => n57);
   U175 : BUF_X1 port map( A => n1576, Z => n1723);
   U176 : BUF_X1 port map( A => n1574, Z => n1719);
   U189 : BUF_X1 port map( A => n1578, Z => n1727);
   U190 : BUF_X1 port map( A => n1580, Z => n1731);
   U191 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n66, ZN => n58);
   U192 : AND2_X1 port map( A1 => n902, A2 => ADD_RD2(0), ZN => n59);
   U193 : AND2_X1 port map( A1 => n903, A2 => ADD_RD2(0), ZN => n60);
   U194 : AND2_X1 port map( A1 => n900, A2 => ADD_RD2(0), ZN => n61);
   U195 : AND2_X1 port map( A1 => n67, A2 => ADD_RD1(0), ZN => n62);
   U196 : AND2_X1 port map( A1 => n68, A2 => ADD_RD1(0), ZN => n63);
   U197 : AND2_X1 port map( A1 => n65, A2 => ADD_RD1(0), ZN => n64);
   U198 : BUF_X1 port map( A => n22, Z => n1742);
   U199 : BUF_X1 port map( A => n25, Z => n1738);
   U200 : INV_X1 port map( A => n1853, ZN => n1851);
   U201 : INV_X1 port map( A => n1853, ZN => n1850);
   U202 : INV_X1 port map( A => n1853, ZN => n1852);
   U203 : BUF_X1 port map( A => n1678, Z => n1693);
   U204 : BUF_X1 port map( A => n1679, Z => n1690);
   U205 : BUF_X1 port map( A => n1679, Z => n1689);
   U206 : BUF_X1 port map( A => n1680, Z => n1686);
   U207 : BUF_X1 port map( A => n1680, Z => n1685);
   U208 : BUF_X1 port map( A => n843, Z => n858);
   U209 : BUF_X1 port map( A => n844, Z => n855);
   U210 : BUF_X1 port map( A => n844, Z => n854);
   U211 : BUF_X1 port map( A => n845, Z => n851);
   U212 : BUF_X1 port map( A => n845, Z => n850);
   U213 : BUF_X1 port map( A => n1678, Z => n1692);
   U214 : BUF_X1 port map( A => n1678, Z => n1691);
   U215 : BUF_X1 port map( A => n1679, Z => n1688);
   U216 : BUF_X1 port map( A => n1680, Z => n1687);
   U217 : BUF_X1 port map( A => n843, Z => n857);
   U218 : BUF_X1 port map( A => n843, Z => n856);
   U219 : BUF_X1 port map( A => n844, Z => n853);
   U220 : BUF_X1 port map( A => n845, Z => n852);
   U221 : BUF_X1 port map( A => n1660, Z => n1675);
   U222 : BUF_X1 port map( A => n1661, Z => n1672);
   U223 : BUF_X1 port map( A => n1661, Z => n1671);
   U224 : BUF_X1 port map( A => n1662, Z => n1668);
   U225 : BUF_X1 port map( A => n1662, Z => n1667);
   U226 : BUF_X1 port map( A => n825, Z => n840);
   U227 : BUF_X1 port map( A => n826, Z => n837);
   U228 : BUF_X1 port map( A => n826, Z => n836);
   U229 : BUF_X1 port map( A => n827, Z => n833);
   U230 : BUF_X1 port map( A => n827, Z => n832);
   U231 : BUF_X1 port map( A => n1660, Z => n1674);
   U232 : BUF_X1 port map( A => n1660, Z => n1673);
   U233 : BUF_X1 port map( A => n1661, Z => n1670);
   U234 : BUF_X1 port map( A => n1662, Z => n1669);
   U235 : BUF_X1 port map( A => n825, Z => n839);
   U236 : BUF_X1 port map( A => n825, Z => n838);
   U237 : BUF_X1 port map( A => n826, Z => n835);
   U238 : BUF_X1 port map( A => n827, Z => n834);
   U239 : BUF_X1 port map( A => n1837, Z => n1836);
   U240 : BUF_X1 port map( A => n1832, Z => n1831);
   U241 : BUF_X1 port map( A => n1827, Z => n1826);
   U242 : BUF_X1 port map( A => n1822, Z => n1821);
   U243 : BUF_X1 port map( A => n1817, Z => n1816);
   U244 : BUF_X1 port map( A => n1812, Z => n1811);
   U245 : BUF_X1 port map( A => n1807, Z => n1806);
   U246 : BUF_X1 port map( A => n1802, Z => n1801);
   U247 : BUF_X1 port map( A => n1797, Z => n1796);
   U248 : BUF_X1 port map( A => n1792, Z => n1791);
   U249 : BUF_X1 port map( A => n1787, Z => n1786);
   U250 : BUF_X1 port map( A => n1782, Z => n1781);
   U251 : BUF_X1 port map( A => n1777, Z => n1776);
   U252 : BUF_X1 port map( A => n1773, Z => n1772);
   U253 : BUF_X1 port map( A => n1770, Z => n1769);
   U254 : BUF_X1 port map( A => n1767, Z => n1766);
   U255 : BUF_X1 port map( A => n1764, Z => n1763);
   U256 : BUF_X1 port map( A => n1761, Z => n1760);
   U257 : BUF_X1 port map( A => n1758, Z => n1757);
   U258 : BUF_X1 port map( A => n1755, Z => n1754);
   U259 : BUF_X1 port map( A => n1752, Z => n1751);
   U260 : BUF_X1 port map( A => n1749, Z => n1748);
   U261 : BUF_X1 port map( A => n1837, Z => n1835);
   U262 : BUF_X1 port map( A => n1832, Z => n1830);
   U263 : BUF_X1 port map( A => n1827, Z => n1825);
   U264 : BUF_X1 port map( A => n1822, Z => n1820);
   U265 : BUF_X1 port map( A => n1817, Z => n1815);
   U266 : BUF_X1 port map( A => n1812, Z => n1810);
   U267 : BUF_X1 port map( A => n1807, Z => n1805);
   U268 : BUF_X1 port map( A => n1802, Z => n1800);
   U269 : BUF_X1 port map( A => n1797, Z => n1795);
   U270 : BUF_X1 port map( A => n1792, Z => n1790);
   U271 : BUF_X1 port map( A => n1787, Z => n1785);
   U272 : BUF_X1 port map( A => n1782, Z => n1780);
   U273 : BUF_X1 port map( A => n1777, Z => n1775);
   U274 : BUF_X1 port map( A => n1773, Z => n1771);
   U275 : BUF_X1 port map( A => n1770, Z => n1768);
   U276 : BUF_X1 port map( A => n1767, Z => n1765);
   U277 : BUF_X1 port map( A => n1764, Z => n1762);
   U278 : BUF_X1 port map( A => n1761, Z => n1759);
   U279 : BUF_X1 port map( A => n1758, Z => n1756);
   U280 : BUF_X1 port map( A => n1755, Z => n1753);
   U281 : BUF_X1 port map( A => n1752, Z => n1750);
   U282 : BUF_X1 port map( A => n1749, Z => n1747);
   U283 : BUF_X1 port map( A => n1842, Z => n1841);
   U284 : BUF_X1 port map( A => n1842, Z => n1840);
   U285 : BUF_X1 port map( A => n1847, Z => n1846);
   U286 : BUF_X1 port map( A => n1847, Z => n1845);
   U287 : BUF_X1 port map( A => RESET, Z => n1849);
   U288 : BUF_X1 port map( A => n1695, Z => n1705);
   U289 : BUF_X1 port map( A => n1695, Z => n1704);
   U290 : BUF_X1 port map( A => n860, Z => n870);
   U291 : BUF_X1 port map( A => n860, Z => n869);
   U292 : BUF_X1 port map( A => n1697, Z => n1700);
   U293 : BUF_X1 port map( A => n862, Z => n865);
   U294 : BUF_X1 port map( A => n1696, Z => n1702);
   U295 : BUF_X1 port map( A => n1696, Z => n1701);
   U296 : BUF_X1 port map( A => n1697, Z => n1699);
   U297 : BUF_X1 port map( A => n861, Z => n867);
   U298 : BUF_X1 port map( A => n861, Z => n866);
   U299 : BUF_X1 port map( A => n862, Z => n864);
   U300 : BUF_X1 port map( A => n1696, Z => n1703);
   U301 : BUF_X1 port map( A => n861, Z => n868);
   U302 : BUF_X1 port map( A => n1642, Z => n1657);
   U303 : BUF_X1 port map( A => n1606, Z => n1621);
   U304 : BUF_X1 port map( A => n1707, Z => n1716);
   U305 : BUF_X1 port map( A => n1643, Z => n1654);
   U306 : BUF_X1 port map( A => n1607, Z => n1618);
   U307 : BUF_X1 port map( A => n1643, Z => n1653);
   U308 : BUF_X1 port map( A => n1607, Z => n1617);
   U309 : BUF_X1 port map( A => n1708, Z => n1713);
   U310 : BUF_X1 port map( A => n1644, Z => n1650);
   U311 : BUF_X1 port map( A => n1608, Z => n1614);
   U312 : BUF_X1 port map( A => n1644, Z => n1649);
   U313 : BUF_X1 port map( A => n1608, Z => n1613);
   U314 : BUF_X1 port map( A => n807, Z => n822);
   U315 : BUF_X1 port map( A => n771, Z => n786);
   U316 : BUF_X1 port map( A => n872, Z => n881);
   U317 : BUF_X1 port map( A => n808, Z => n819);
   U318 : BUF_X1 port map( A => n772, Z => n783);
   U319 : BUF_X1 port map( A => n808, Z => n818);
   U320 : BUF_X1 port map( A => n772, Z => n782);
   U321 : BUF_X1 port map( A => n873, Z => n878);
   U322 : BUF_X1 port map( A => n809, Z => n815);
   U323 : BUF_X1 port map( A => n773, Z => n779);
   U324 : BUF_X1 port map( A => n809, Z => n814);
   U325 : BUF_X1 port map( A => n773, Z => n778);
   U326 : BUF_X1 port map( A => n1707, Z => n1718);
   U327 : BUF_X1 port map( A => n1642, Z => n1656);
   U328 : BUF_X1 port map( A => n1606, Z => n1620);
   U329 : BUF_X1 port map( A => n1707, Z => n1717);
   U330 : BUF_X1 port map( A => n1642, Z => n1655);
   U331 : BUF_X1 port map( A => n1606, Z => n1619);
   U332 : BUF_X1 port map( A => n1708, Z => n1715);
   U333 : BUF_X1 port map( A => n1643, Z => n1652);
   U334 : BUF_X1 port map( A => n1607, Z => n1616);
   U335 : BUF_X1 port map( A => n1708, Z => n1714);
   U336 : BUF_X1 port map( A => n1644, Z => n1651);
   U337 : BUF_X1 port map( A => n1608, Z => n1615);
   U338 : BUF_X1 port map( A => n1709, Z => n1712);
   U339 : BUF_X1 port map( A => n1681, Z => n1684);
   U340 : BUF_X1 port map( A => n1709, Z => n1711);
   U341 : BUF_X1 port map( A => n1681, Z => n1683);
   U342 : BUF_X1 port map( A => n872, Z => n883);
   U343 : BUF_X1 port map( A => n807, Z => n821);
   U344 : BUF_X1 port map( A => n771, Z => n785);
   U345 : BUF_X1 port map( A => n872, Z => n882);
   U346 : BUF_X1 port map( A => n807, Z => n820);
   U347 : BUF_X1 port map( A => n771, Z => n784);
   U348 : BUF_X1 port map( A => n873, Z => n880);
   U349 : BUF_X1 port map( A => n808, Z => n817);
   U350 : BUF_X1 port map( A => n772, Z => n781);
   U351 : BUF_X1 port map( A => n873, Z => n879);
   U352 : BUF_X1 port map( A => n809, Z => n816);
   U353 : BUF_X1 port map( A => n773, Z => n780);
   U354 : BUF_X1 port map( A => n874, Z => n877);
   U355 : BUF_X1 port map( A => n846, Z => n849);
   U356 : BUF_X1 port map( A => n874, Z => n876);
   U357 : BUF_X1 port map( A => n846, Z => n848);
   U358 : BUF_X1 port map( A => n1624, Z => n1639);
   U359 : BUF_X1 port map( A => n1588, Z => n1603);
   U360 : BUF_X1 port map( A => n1625, Z => n1636);
   U361 : BUF_X1 port map( A => n1589, Z => n1600);
   U362 : BUF_X1 port map( A => n1625, Z => n1635);
   U363 : BUF_X1 port map( A => n1589, Z => n1599);
   U364 : BUF_X1 port map( A => n1626, Z => n1632);
   U365 : BUF_X1 port map( A => n1590, Z => n1596);
   U366 : BUF_X1 port map( A => n1626, Z => n1631);
   U367 : BUF_X1 port map( A => n1590, Z => n1595);
   U368 : BUF_X1 port map( A => n789, Z => n804);
   U369 : BUF_X1 port map( A => n753, Z => n768);
   U370 : BUF_X1 port map( A => n790, Z => n801);
   U371 : BUF_X1 port map( A => n754, Z => n765);
   U372 : BUF_X1 port map( A => n790, Z => n800);
   U373 : BUF_X1 port map( A => n754, Z => n764);
   U374 : BUF_X1 port map( A => n791, Z => n797);
   U375 : BUF_X1 port map( A => n755, Z => n761);
   U376 : BUF_X1 port map( A => n791, Z => n796);
   U377 : BUF_X1 port map( A => n755, Z => n760);
   U378 : BUF_X1 port map( A => n1624, Z => n1638);
   U379 : BUF_X1 port map( A => n1588, Z => n1602);
   U380 : BUF_X1 port map( A => n1624, Z => n1637);
   U381 : BUF_X1 port map( A => n1588, Z => n1601);
   U382 : BUF_X1 port map( A => n1625, Z => n1634);
   U383 : BUF_X1 port map( A => n1589, Z => n1598);
   U384 : BUF_X1 port map( A => n1626, Z => n1633);
   U385 : BUF_X1 port map( A => n1590, Z => n1597);
   U386 : BUF_X1 port map( A => n1663, Z => n1666);
   U387 : BUF_X1 port map( A => n1663, Z => n1665);
   U388 : BUF_X1 port map( A => n789, Z => n803);
   U389 : BUF_X1 port map( A => n753, Z => n767);
   U390 : BUF_X1 port map( A => n789, Z => n802);
   U391 : BUF_X1 port map( A => n753, Z => n766);
   U392 : BUF_X1 port map( A => n790, Z => n799);
   U393 : BUF_X1 port map( A => n754, Z => n763);
   U394 : BUF_X1 port map( A => n791, Z => n798);
   U395 : BUF_X1 port map( A => n755, Z => n762);
   U396 : BUF_X1 port map( A => n828, Z => n831);
   U397 : BUF_X1 port map( A => n828, Z => n830);
   U398 : BUF_X1 port map( A => n1697, Z => n1698);
   U399 : BUF_X1 port map( A => n862, Z => n863);
   U400 : BUF_X1 port map( A => n1709, Z => n1710);
   U401 : BUF_X1 port map( A => n874, Z => n875);
   U402 : BUF_X1 port map( A => n1681, Z => n1682);
   U403 : BUF_X1 port map( A => n846, Z => n847);
   U404 : BUF_X1 port map( A => n1663, Z => n1664);
   U405 : BUF_X1 port map( A => n828, Z => n829);
   U406 : BUF_X1 port map( A => n1838, Z => n1834);
   U407 : BUF_X1 port map( A => n6, Z => n1838);
   U408 : BUF_X1 port map( A => n1833, Z => n1829);
   U409 : BUF_X1 port map( A => n7, Z => n1833);
   U410 : BUF_X1 port map( A => n1828, Z => n1824);
   U411 : BUF_X1 port map( A => n28, Z => n1828);
   U412 : BUF_X1 port map( A => n1823, Z => n1819);
   U413 : BUF_X1 port map( A => n29, Z => n1823);
   U414 : BUF_X1 port map( A => n1818, Z => n1814);
   U415 : BUF_X1 port map( A => n30, Z => n1818);
   U416 : BUF_X1 port map( A => n1813, Z => n1809);
   U417 : BUF_X1 port map( A => n31, Z => n1813);
   U418 : BUF_X1 port map( A => n1808, Z => n1804);
   U419 : BUF_X1 port map( A => n32, Z => n1808);
   U420 : BUF_X1 port map( A => n1803, Z => n1799);
   U421 : BUF_X1 port map( A => n33, Z => n1803);
   U422 : BUF_X1 port map( A => n1798, Z => n1794);
   U423 : BUF_X1 port map( A => n34, Z => n1798);
   U424 : BUF_X1 port map( A => n1793, Z => n1789);
   U425 : BUF_X1 port map( A => n35, Z => n1793);
   U426 : BUF_X1 port map( A => n1788, Z => n1784);
   U427 : BUF_X1 port map( A => n36, Z => n1788);
   U428 : BUF_X1 port map( A => n1783, Z => n1779);
   U429 : BUF_X1 port map( A => n37, Z => n1783);
   U430 : BUF_X1 port map( A => n1778, Z => n1774);
   U431 : BUF_X1 port map( A => n38, Z => n1778);
   U432 : BUF_X1 port map( A => n1843, Z => n1839);
   U433 : BUF_X1 port map( A => n39, Z => n1843);
   U434 : BUF_X1 port map( A => n1848, Z => n1844);
   U435 : BUF_X1 port map( A => n1, Z => n1848);
   U436 : BUF_X1 port map( A => n2, Z => n1676);
   U437 : BUF_X1 port map( A => n5, Z => n1658);
   U438 : BUF_X1 port map( A => n3, Z => n841);
   U439 : BUF_X1 port map( A => n4, Z => n823);
   U440 : BUF_X1 port map( A => n1694, Z => n1695);
   U441 : BUF_X1 port map( A => n859, Z => n860);
   U442 : BUF_X1 port map( A => n1743, Z => n1744);
   U443 : BUF_X1 port map( A => n1743, Z => n1745);
   U444 : BUF_X1 port map( A => n1743, Z => n1746);
   U445 : BUF_X1 port map( A => n1645, Z => n1648);
   U446 : BUF_X1 port map( A => n1609, Z => n1612);
   U447 : BUF_X1 port map( A => n1645, Z => n1647);
   U448 : BUF_X1 port map( A => n1609, Z => n1611);
   U449 : BUF_X1 port map( A => n810, Z => n813);
   U450 : BUF_X1 port map( A => n774, Z => n777);
   U451 : BUF_X1 port map( A => n810, Z => n812);
   U452 : BUF_X1 port map( A => n774, Z => n776);
   U453 : BUF_X1 port map( A => n1627, Z => n1630);
   U454 : BUF_X1 port map( A => n1591, Z => n1594);
   U455 : BUF_X1 port map( A => n1627, Z => n1629);
   U456 : BUF_X1 port map( A => n1591, Z => n1593);
   U457 : BUF_X1 port map( A => n792, Z => n795);
   U458 : BUF_X1 port map( A => n756, Z => n759);
   U459 : BUF_X1 port map( A => n792, Z => n794);
   U460 : BUF_X1 port map( A => n756, Z => n758);
   U461 : BUF_X1 port map( A => n1645, Z => n1646);
   U462 : BUF_X1 port map( A => n1609, Z => n1610);
   U463 : BUF_X1 port map( A => n810, Z => n811);
   U464 : BUF_X1 port map( A => n774, Z => n775);
   U465 : BUF_X1 port map( A => n1627, Z => n1628);
   U466 : BUF_X1 port map( A => n1591, Z => n1592);
   U467 : BUF_X1 port map( A => n792, Z => n793);
   U468 : BUF_X1 port map( A => n756, Z => n757);
   U469 : NAND2_X1 port map( A1 => n1849, A2 => n1859, ZN => n8);
   U470 : BUF_X1 port map( A => n59, Z => n1640);
   U471 : BUF_X1 port map( A => n60, Z => n1622);
   U472 : BUF_X1 port map( A => n61, Z => n1604);
   U473 : BUF_X1 port map( A => n57, Z => n1586);
   U474 : BUF_X1 port map( A => n62, Z => n805);
   U475 : BUF_X1 port map( A => n63, Z => n787);
   U476 : BUF_X1 port map( A => n64, Z => n769);
   U477 : BUF_X1 port map( A => n58, Z => n751);
   U478 : AND2_X1 port map( A1 => N290, A2 => n1741, ZN => N291);
   U479 : AND2_X1 port map( A1 => N289, A2 => n1741, ZN => N292);
   U480 : AND2_X1 port map( A1 => N288, A2 => n1741, ZN => N293);
   U481 : AND2_X1 port map( A1 => N287, A2 => n1741, ZN => N294);
   U482 : AND2_X1 port map( A1 => N286, A2 => n1741, ZN => N295);
   U483 : AND2_X1 port map( A1 => N285, A2 => n1741, ZN => N296);
   U484 : AND2_X1 port map( A1 => N284, A2 => n1741, ZN => N297);
   U485 : AND2_X1 port map( A1 => N283, A2 => n1741, ZN => N298);
   U486 : AND2_X1 port map( A1 => N282, A2 => n1741, ZN => N299);
   U487 : AND2_X1 port map( A1 => N281, A2 => n1741, ZN => N300);
   U488 : AND2_X1 port map( A1 => N280, A2 => n1740, ZN => N301);
   U489 : AND2_X1 port map( A1 => N279, A2 => n1740, ZN => N302);
   U490 : AND2_X1 port map( A1 => N278, A2 => n1740, ZN => N303);
   U491 : AND2_X1 port map( A1 => N277, A2 => n1740, ZN => N304);
   U492 : AND2_X1 port map( A1 => N276, A2 => n1740, ZN => N305);
   U493 : AND2_X1 port map( A1 => N275, A2 => n1740, ZN => N306);
   U494 : AND2_X1 port map( A1 => N274, A2 => n1740, ZN => N307);
   U495 : AND2_X1 port map( A1 => N273, A2 => n1740, ZN => N308);
   U496 : AND2_X1 port map( A1 => N272, A2 => n1740, ZN => N309);
   U497 : AND2_X1 port map( A1 => N271, A2 => n1740, ZN => N310);
   U498 : AND2_X1 port map( A1 => N270, A2 => n1740, ZN => N311);
   U499 : AND2_X1 port map( A1 => N269, A2 => n1739, ZN => N312);
   U500 : AND2_X1 port map( A1 => N268, A2 => n1739, ZN => N313);
   U501 : AND2_X1 port map( A1 => N267, A2 => n1739, ZN => N314);
   U502 : AND2_X1 port map( A1 => N266, A2 => n1739, ZN => N315);
   U503 : AND2_X1 port map( A1 => N265, A2 => n1739, ZN => N316);
   U504 : AND2_X1 port map( A1 => N264, A2 => n1739, ZN => N317);
   U505 : AND2_X1 port map( A1 => N263, A2 => n1739, ZN => N318);
   U506 : AND2_X1 port map( A1 => N262, A2 => n1739, ZN => N319);
   U507 : AND2_X1 port map( A1 => N261, A2 => n1739, ZN => N320);
   U508 : AND2_X1 port map( A1 => N260, A2 => n1739, ZN => N321);
   U509 : AND2_X1 port map( A1 => N259, A2 => n1739, ZN => N322);
   U510 : AND2_X1 port map( A1 => N224, A2 => n1737, ZN => N225);
   U511 : AND2_X1 port map( A1 => N223, A2 => n1737, ZN => N226);
   U512 : AND2_X1 port map( A1 => N222, A2 => n1737, ZN => N227);
   U513 : AND2_X1 port map( A1 => N221, A2 => n1737, ZN => N228);
   U514 : AND2_X1 port map( A1 => N220, A2 => n1737, ZN => N229);
   U515 : AND2_X1 port map( A1 => N219, A2 => n1737, ZN => N230);
   U516 : AND2_X1 port map( A1 => N218, A2 => n1737, ZN => N231);
   U517 : AND2_X1 port map( A1 => N217, A2 => n1737, ZN => N232);
   U518 : AND2_X1 port map( A1 => N216, A2 => n1737, ZN => N233);
   U519 : AND2_X1 port map( A1 => N215, A2 => n1737, ZN => N234);
   U520 : AND2_X1 port map( A1 => N214, A2 => n1736, ZN => N235);
   U521 : AND2_X1 port map( A1 => N213, A2 => n1736, ZN => N236);
   U522 : AND2_X1 port map( A1 => N212, A2 => n1736, ZN => N237);
   U523 : AND2_X1 port map( A1 => N211, A2 => n1736, ZN => N238);
   U524 : AND2_X1 port map( A1 => N210, A2 => n1736, ZN => N239);
   U525 : AND2_X1 port map( A1 => N209, A2 => n1736, ZN => N240);
   U526 : AND2_X1 port map( A1 => N208, A2 => n1736, ZN => N241);
   U527 : AND2_X1 port map( A1 => N207, A2 => n1736, ZN => N242);
   U528 : AND2_X1 port map( A1 => N206, A2 => n1736, ZN => N243);
   U529 : AND2_X1 port map( A1 => N205, A2 => n1736, ZN => N244);
   U530 : AND2_X1 port map( A1 => N204, A2 => n1736, ZN => N245);
   U531 : AND2_X1 port map( A1 => N203, A2 => n1735, ZN => N246);
   U532 : AND2_X1 port map( A1 => N202, A2 => n1735, ZN => N247);
   U533 : AND2_X1 port map( A1 => N201, A2 => n1735, ZN => N248);
   U534 : AND2_X1 port map( A1 => N200, A2 => n1735, ZN => N249);
   U535 : AND2_X1 port map( A1 => N199, A2 => n1735, ZN => N250);
   U536 : AND2_X1 port map( A1 => N198, A2 => n1735, ZN => N251);
   U537 : AND2_X1 port map( A1 => N197, A2 => n1735, ZN => N252);
   U538 : AND2_X1 port map( A1 => N196, A2 => n1735, ZN => N253);
   U539 : AND2_X1 port map( A1 => N195, A2 => n1735, ZN => N254);
   U540 : AND2_X1 port map( A1 => N194, A2 => n1735, ZN => N255);
   U541 : AND2_X1 port map( A1 => N193, A2 => n1735, ZN => N256);
   U542 : BUF_X1 port map( A => n1723, Z => n1726);
   U543 : BUF_X1 port map( A => n1723, Z => n1725);
   U544 : BUF_X1 port map( A => n888, Z => n891);
   U545 : BUF_X1 port map( A => n888, Z => n890);
   U546 : BUF_X1 port map( A => n1742, Z => n1740);
   U547 : BUF_X1 port map( A => n1742, Z => n1739);
   U548 : BUF_X1 port map( A => n1738, Z => n1736);
   U549 : BUF_X1 port map( A => n1738, Z => n1735);
   U550 : BUF_X1 port map( A => n1719, Z => n1722);
   U551 : BUF_X1 port map( A => n1719, Z => n1721);
   U552 : BUF_X1 port map( A => n884, Z => n887);
   U553 : BUF_X1 port map( A => n884, Z => n886);
   U554 : BUF_X1 port map( A => n1731, Z => n1734);
   U555 : BUF_X1 port map( A => n1731, Z => n1733);
   U556 : BUF_X1 port map( A => n896, Z => n899);
   U557 : BUF_X1 port map( A => n896, Z => n898);
   U558 : BUF_X1 port map( A => n1727, Z => n1730);
   U559 : BUF_X1 port map( A => n892, Z => n895);
   U560 : BUF_X1 port map( A => n1727, Z => n1729);
   U561 : BUF_X1 port map( A => n892, Z => n894);
   U562 : BUF_X1 port map( A => n1723, Z => n1724);
   U563 : BUF_X1 port map( A => n888, Z => n889);
   U564 : BUF_X1 port map( A => n1742, Z => n1741);
   U565 : BUF_X1 port map( A => n1738, Z => n1737);
   U566 : BUF_X1 port map( A => n1719, Z => n1720);
   U567 : BUF_X1 port map( A => n884, Z => n885);
   U568 : BUF_X1 port map( A => n1731, Z => n1732);
   U569 : BUF_X1 port map( A => n896, Z => n897);
   U570 : BUF_X1 port map( A => n1727, Z => n1728);
   U571 : BUF_X1 port map( A => n892, Z => n893);
   U572 : NAND2_X1 port map( A1 => REGISTERS_2_31_port, A2 => n1703, ZN => 
                           n1563);
   U573 : NAND2_X1 port map( A1 => REGISTERS_2_31_port, A2 => n868, ZN => n728)
                           ;
   U574 : NAND2_X1 port map( A1 => REGISTERS_2_0_port, A2 => n1705, ZN => n912)
                           ;
   U575 : NAND2_X1 port map( A1 => REGISTERS_2_1_port, A2 => n1705, ZN => n933)
                           ;
   U576 : NAND2_X1 port map( A1 => REGISTERS_2_2_port, A2 => n1705, ZN => n954)
                           ;
   U577 : NAND2_X1 port map( A1 => REGISTERS_2_3_port, A2 => n1705, ZN => n975)
                           ;
   U578 : NAND2_X1 port map( A1 => REGISTERS_2_4_port, A2 => n1705, ZN => n996)
                           ;
   U579 : NAND2_X1 port map( A1 => REGISTERS_2_5_port, A2 => n1705, ZN => n1017
                           );
   U580 : NAND2_X1 port map( A1 => REGISTERS_2_6_port, A2 => n1705, ZN => n1038
                           );
   U581 : NAND2_X1 port map( A1 => REGISTERS_2_7_port, A2 => n1705, ZN => n1059
                           );
   U582 : NAND2_X1 port map( A1 => REGISTERS_2_8_port, A2 => n1705, ZN => n1080
                           );
   U583 : NAND2_X1 port map( A1 => REGISTERS_2_9_port, A2 => n1705, ZN => n1101
                           );
   U584 : NAND2_X1 port map( A1 => REGISTERS_2_10_port, A2 => n1705, ZN => 
                           n1122);
   U585 : NAND2_X1 port map( A1 => REGISTERS_2_11_port, A2 => n1705, ZN => 
                           n1143);
   U586 : NAND2_X1 port map( A1 => REGISTERS_2_12_port, A2 => n1704, ZN => 
                           n1164);
   U587 : NAND2_X1 port map( A1 => REGISTERS_2_13_port, A2 => n1704, ZN => 
                           n1185);
   U588 : NAND2_X1 port map( A1 => REGISTERS_2_14_port, A2 => n1704, ZN => 
                           n1206);
   U589 : NAND2_X1 port map( A1 => REGISTERS_2_15_port, A2 => n1704, ZN => 
                           n1227);
   U590 : NAND2_X1 port map( A1 => REGISTERS_2_16_port, A2 => n1704, ZN => 
                           n1248);
   U591 : NAND2_X1 port map( A1 => REGISTERS_2_17_port, A2 => n1704, ZN => 
                           n1269);
   U592 : NAND2_X1 port map( A1 => REGISTERS_2_18_port, A2 => n1704, ZN => 
                           n1290);
   U593 : NAND2_X1 port map( A1 => REGISTERS_2_19_port, A2 => n1704, ZN => 
                           n1311);
   U594 : NAND2_X1 port map( A1 => REGISTERS_2_20_port, A2 => n1704, ZN => 
                           n1332);
   U595 : NAND2_X1 port map( A1 => REGISTERS_2_21_port, A2 => n1704, ZN => 
                           n1353);
   U596 : NAND2_X1 port map( A1 => REGISTERS_2_22_port, A2 => n1704, ZN => 
                           n1374);
   U597 : NAND2_X1 port map( A1 => REGISTERS_2_23_port, A2 => n1704, ZN => 
                           n1395);
   U598 : NAND2_X1 port map( A1 => REGISTERS_2_24_port, A2 => n1703, ZN => 
                           n1416);
   U599 : NAND2_X1 port map( A1 => REGISTERS_2_25_port, A2 => n1703, ZN => 
                           n1437);
   U600 : NAND2_X1 port map( A1 => REGISTERS_2_26_port, A2 => n1703, ZN => 
                           n1458);
   U601 : NAND2_X1 port map( A1 => REGISTERS_2_27_port, A2 => n1703, ZN => 
                           n1479);
   U602 : NAND2_X1 port map( A1 => REGISTERS_2_28_port, A2 => n1703, ZN => 
                           n1500);
   U603 : NAND2_X1 port map( A1 => REGISTERS_2_29_port, A2 => n1703, ZN => 
                           n1521);
   U604 : NAND2_X1 port map( A1 => REGISTERS_2_30_port, A2 => n1703, ZN => 
                           n1542);
   U605 : NAND2_X1 port map( A1 => REGISTERS_2_0_port, A2 => n870, ZN => n77);
   U606 : NAND2_X1 port map( A1 => REGISTERS_2_1_port, A2 => n870, ZN => n98);
   U607 : NAND2_X1 port map( A1 => REGISTERS_2_2_port, A2 => n870, ZN => n119);
   U608 : NAND2_X1 port map( A1 => REGISTERS_2_3_port, A2 => n870, ZN => n140);
   U609 : NAND2_X1 port map( A1 => REGISTERS_2_4_port, A2 => n870, ZN => n161);
   U610 : NAND2_X1 port map( A1 => REGISTERS_2_5_port, A2 => n870, ZN => n182);
   U611 : NAND2_X1 port map( A1 => REGISTERS_2_6_port, A2 => n870, ZN => 
                           n203_port);
   U612 : NAND2_X1 port map( A1 => REGISTERS_2_7_port, A2 => n870, ZN => 
                           n224_port);
   U613 : NAND2_X1 port map( A1 => REGISTERS_2_8_port, A2 => n870, ZN => 
                           n245_port);
   U614 : NAND2_X1 port map( A1 => REGISTERS_2_9_port, A2 => n870, ZN => 
                           n266_port);
   U615 : NAND2_X1 port map( A1 => REGISTERS_2_10_port, A2 => n870, ZN => 
                           n287_port);
   U616 : NAND2_X1 port map( A1 => REGISTERS_2_11_port, A2 => n870, ZN => 
                           n308_port);
   U617 : NAND2_X1 port map( A1 => REGISTERS_2_12_port, A2 => n869, ZN => 
                           n329_port);
   U618 : NAND2_X1 port map( A1 => REGISTERS_2_13_port, A2 => n869, ZN => 
                           n350_port);
   U619 : NAND2_X1 port map( A1 => REGISTERS_2_14_port, A2 => n869, ZN => n371)
                           ;
   U620 : NAND2_X1 port map( A1 => REGISTERS_2_15_port, A2 => n869, ZN => n392)
                           ;
   U621 : NAND2_X1 port map( A1 => REGISTERS_2_16_port, A2 => n869, ZN => n413)
                           ;
   U622 : NAND2_X1 port map( A1 => REGISTERS_2_17_port, A2 => n869, ZN => n434)
                           ;
   U623 : NAND2_X1 port map( A1 => REGISTERS_2_18_port, A2 => n869, ZN => n455)
                           ;
   U624 : NAND2_X1 port map( A1 => REGISTERS_2_19_port, A2 => n869, ZN => n476)
                           ;
   U625 : NAND2_X1 port map( A1 => REGISTERS_2_20_port, A2 => n869, ZN => n497)
                           ;
   U626 : NAND2_X1 port map( A1 => REGISTERS_2_21_port, A2 => n869, ZN => n518)
                           ;
   U627 : NAND2_X1 port map( A1 => REGISTERS_2_22_port, A2 => n869, ZN => n539)
                           ;
   U628 : NAND2_X1 port map( A1 => REGISTERS_2_23_port, A2 => n869, ZN => n560)
                           ;
   U629 : NAND2_X1 port map( A1 => REGISTERS_2_24_port, A2 => n868, ZN => n581)
                           ;
   U630 : NAND2_X1 port map( A1 => REGISTERS_2_25_port, A2 => n868, ZN => n602)
                           ;
   U631 : NAND2_X1 port map( A1 => REGISTERS_2_26_port, A2 => n868, ZN => n623)
                           ;
   U632 : NAND2_X1 port map( A1 => REGISTERS_2_27_port, A2 => n868, ZN => n644)
                           ;
   U633 : NAND2_X1 port map( A1 => REGISTERS_2_28_port, A2 => n868, ZN => n665)
                           ;
   U634 : NAND2_X1 port map( A1 => REGISTERS_2_29_port, A2 => n868, ZN => n686)
                           ;
   U635 : NAND2_X1 port map( A1 => REGISTERS_2_30_port, A2 => n868, ZN => n707)
                           ;
   U636 : INV_X1 port map( A => ADD_RD2(0), ZN => n1582);
   U637 : INV_X1 port map( A => ADD_RD2(3), ZN => n1585);
   U638 : INV_X1 port map( A => ADD_RD2(2), ZN => n1584);
   U639 : INV_X1 port map( A => ADD_RD1(0), ZN => n747);
   U640 : INV_X1 port map( A => ADD_RD2(1), ZN => n1583);
   U641 : AND3_X1 port map( A1 => ENABLE, A2 => n1859, A3 => WR, ZN => n17);
   U642 : INV_X1 port map( A => ADD_RD1(3), ZN => n750);
   U643 : INV_X1 port map( A => ADD_RD1(2), ZN => n749);
   U644 : INV_X1 port map( A => ADD_RD1(1), ZN => n748);
   U645 : INV_X1 port map( A => ADD_WR(0), ZN => n1858);
   U646 : INV_X1 port map( A => ADD_WR(2), ZN => n1856);
   U647 : INV_X1 port map( A => ADD_WR(1), ZN => n1857);
   U648 : AND2_X1 port map( A1 => RD2, A2 => n23, ZN => n22);
   U649 : OR4_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => ADD_RD2(2)
                           , A4 => n24, ZN => n23);
   U650 : OR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), ZN => n24);
   U651 : AND2_X1 port map( A1 => RD1, A2 => n26, ZN => n25);
   U652 : OR4_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => ADD_RD1(2)
                           , A4 => n27, ZN => n26);
   U653 : OR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n27);
   U654 : INV_X1 port map( A => ADD_WR(4), ZN => n1854);
   U655 : INV_X1 port map( A => ADD_WR(3), ZN => n1855);
   U656 : INV_X1 port map( A => CLK, ZN => n1859);
   U657 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n750, ZN => n745);
   U658 : NOR2_X1 port map( A1 => n749, A2 => ADD_RD1(1), ZN => n65);
   U659 : NOR2_X1 port map( A1 => n749, A2 => n748, ZN => n66);
   U660 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n786, B1 => 
                           REGISTERS_23_0_port, B2 => n768, ZN => n72);
   U661 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n67);
   U662 : NOR2_X1 port map( A1 => n748, A2 => ADD_RD1(2), ZN => n68);
   U663 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n822, B1 => 
                           REGISTERS_19_0_port, B2 => n804, ZN => n71);
   U664 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n858, B1 => 
                           REGISTERS_22_0_port, B2 => n840, ZN => n70);
   U665 : AND2_X1 port map( A1 => n67, A2 => n747, ZN => n733);
   U666 : AND2_X1 port map( A1 => n68, A2 => n747, ZN => n732);
   U667 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n883, B1 => 
                           REGISTERS_18_0_port, B2 => n868, ZN => n69);
   U668 : AND4_X1 port map( A1 => n72, A2 => n71, A3 => n70, A4 => n69, ZN => 
                           n89);
   U669 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n743);
   U670 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n786, B1 => 
                           REGISTERS_31_0_port, B2 => n768, ZN => n76);
   U671 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n822, B1 => 
                           REGISTERS_27_0_port, B2 => n804, ZN => n75);
   U672 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n858, B1 => 
                           REGISTERS_30_0_port, B2 => n840, ZN => n74);
   U673 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n883, B1 => 
                           REGISTERS_26_0_port, B2 => n868, ZN => n73);
   U674 : AND4_X1 port map( A1 => n76, A2 => n75, A3 => n74, A4 => n73, ZN => 
                           n88);
   U675 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n786, B1 => 
                           REGISTERS_7_0_port, B2 => n768, ZN => n80);
   U676 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n822, B1 => 
                           REGISTERS_3_0_port, B2 => n804, ZN => n79);
   U677 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n858, B1 => 
                           REGISTERS_6_0_port, B2 => n840, ZN => n78);
   U678 : NAND4_X1 port map( A1 => n80, A2 => n79, A3 => n78, A4 => n77, ZN => 
                           n86);
   U679 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n741);
   U680 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n786, B1 => 
                           REGISTERS_15_0_port, B2 => n768, ZN => n84);
   U681 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n822, B1 => 
                           REGISTERS_11_0_port, B2 => n804, ZN => n83);
   U682 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n858, B1 => 
                           REGISTERS_14_0_port, B2 => n840, ZN => n82);
   U683 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n883, B1 => 
                           REGISTERS_10_0_port, B2 => n868, ZN => n81);
   U684 : NAND4_X1 port map( A1 => n84, A2 => n83, A3 => n82, A4 => n81, ZN => 
                           n85);
   U685 : NOR2_X1 port map( A1 => n750, A2 => ADD_RD1(4), ZN => n739);
   U686 : AOI22_X1 port map( A1 => n86, A2 => n891, B1 => n85, B2 => n887, ZN 
                           => n87);
   U687 : OAI221_X1 port map( B1 => n899, B2 => n89, C1 => n893, C2 => n88, A 
                           => n87, ZN => N224);
   U688 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n786, B1 => 
                           REGISTERS_23_1_port, B2 => n768, ZN => n93);
   U689 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n822, B1 => 
                           REGISTERS_19_1_port, B2 => n804, ZN => n92);
   U690 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n858, B1 => 
                           REGISTERS_22_1_port, B2 => n840, ZN => n91);
   U691 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n883, B1 => 
                           REGISTERS_18_1_port, B2 => n868, ZN => n90);
   U692 : AND4_X1 port map( A1 => n93, A2 => n92, A3 => n91, A4 => n90, ZN => 
                           n110);
   U693 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n786, B1 => 
                           REGISTERS_31_1_port, B2 => n768, ZN => n97);
   U694 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n822, B1 => 
                           REGISTERS_27_1_port, B2 => n804, ZN => n96);
   U695 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n858, B1 => 
                           REGISTERS_30_1_port, B2 => n840, ZN => n95);
   U696 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n883, B1 => 
                           REGISTERS_26_1_port, B2 => n868, ZN => n94);
   U697 : AND4_X1 port map( A1 => n97, A2 => n96, A3 => n95, A4 => n94, ZN => 
                           n109);
   U698 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n786, B1 => 
                           REGISTERS_7_1_port, B2 => n768, ZN => n101);
   U699 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n822, B1 => 
                           REGISTERS_3_1_port, B2 => n804, ZN => n100);
   U700 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n858, B1 => 
                           REGISTERS_6_1_port, B2 => n840, ZN => n99);
   U701 : NAND4_X1 port map( A1 => n101, A2 => n100, A3 => n99, A4 => n98, ZN 
                           => n107);
   U702 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n786, B1 => 
                           REGISTERS_15_1_port, B2 => n768, ZN => n105);
   U703 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n822, B1 => 
                           REGISTERS_11_1_port, B2 => n804, ZN => n104);
   U704 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n858, B1 => 
                           REGISTERS_14_1_port, B2 => n840, ZN => n103);
   U705 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n883, B1 => 
                           REGISTERS_10_1_port, B2 => n868, ZN => n102);
   U706 : NAND4_X1 port map( A1 => n105, A2 => n104, A3 => n103, A4 => n102, ZN
                           => n106);
   U707 : AOI22_X1 port map( A1 => n107, A2 => n891, B1 => n106, B2 => n887, ZN
                           => n108);
   U708 : OAI221_X1 port map( B1 => n899, B2 => n110, C1 => n893, C2 => n109, A
                           => n108, ZN => N223);
   U709 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n786, B1 => 
                           REGISTERS_23_2_port, B2 => n768, ZN => n114);
   U710 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n822, B1 => 
                           REGISTERS_19_2_port, B2 => n804, ZN => n113);
   U711 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n858, B1 => 
                           REGISTERS_22_2_port, B2 => n840, ZN => n112);
   U712 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n883, B1 => 
                           REGISTERS_18_2_port, B2 => n867, ZN => n111);
   U713 : AND4_X1 port map( A1 => n114, A2 => n113, A3 => n112, A4 => n111, ZN 
                           => n131);
   U714 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n786, B1 => 
                           REGISTERS_31_2_port, B2 => n768, ZN => n118);
   U715 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n822, B1 => 
                           REGISTERS_27_2_port, B2 => n804, ZN => n117);
   U716 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n858, B1 => 
                           REGISTERS_30_2_port, B2 => n840, ZN => n116);
   U717 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n883, B1 => 
                           REGISTERS_26_2_port, B2 => n867, ZN => n115);
   U718 : AND4_X1 port map( A1 => n118, A2 => n117, A3 => n116, A4 => n115, ZN 
                           => n130);
   U719 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n786, B1 => 
                           REGISTERS_7_2_port, B2 => n768, ZN => n122);
   U720 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n822, B1 => 
                           REGISTERS_3_2_port, B2 => n804, ZN => n121);
   U721 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n858, B1 => 
                           REGISTERS_6_2_port, B2 => n840, ZN => n120);
   U722 : NAND4_X1 port map( A1 => n122, A2 => n121, A3 => n120, A4 => n119, ZN
                           => n128);
   U723 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n785, B1 => 
                           REGISTERS_15_2_port, B2 => n767, ZN => n126);
   U724 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n821, B1 => 
                           REGISTERS_11_2_port, B2 => n803, ZN => n125);
   U725 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n857, B1 => 
                           REGISTERS_14_2_port, B2 => n839, ZN => n124);
   U726 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n883, B1 => 
                           REGISTERS_10_2_port, B2 => n867, ZN => n123);
   U727 : NAND4_X1 port map( A1 => n126, A2 => n125, A3 => n124, A4 => n123, ZN
                           => n127);
   U728 : AOI22_X1 port map( A1 => n128, A2 => n891, B1 => n127, B2 => n887, ZN
                           => n129);
   U729 : OAI221_X1 port map( B1 => n899, B2 => n131, C1 => n893, C2 => n130, A
                           => n129, ZN => N222);
   U730 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n785, B1 => 
                           REGISTERS_23_3_port, B2 => n767, ZN => n135);
   U731 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n821, B1 => 
                           REGISTERS_19_3_port, B2 => n803, ZN => n134);
   U732 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n857, B1 => 
                           REGISTERS_22_3_port, B2 => n839, ZN => n133);
   U733 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n883, B1 => 
                           REGISTERS_18_3_port, B2 => n867, ZN => n132);
   U734 : AND4_X1 port map( A1 => n135, A2 => n134, A3 => n133, A4 => n132, ZN 
                           => n152);
   U735 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n785, B1 => 
                           REGISTERS_31_3_port, B2 => n767, ZN => n139);
   U736 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n821, B1 => 
                           REGISTERS_27_3_port, B2 => n803, ZN => n138);
   U737 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n857, B1 => 
                           REGISTERS_30_3_port, B2 => n839, ZN => n137);
   U738 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n883, B1 => 
                           REGISTERS_26_3_port, B2 => n867, ZN => n136);
   U739 : AND4_X1 port map( A1 => n139, A2 => n138, A3 => n137, A4 => n136, ZN 
                           => n151);
   U740 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n785, B1 => 
                           REGISTERS_7_3_port, B2 => n767, ZN => n143);
   U741 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n821, B1 => 
                           REGISTERS_3_3_port, B2 => n803, ZN => n142);
   U742 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n857, B1 => 
                           REGISTERS_6_3_port, B2 => n839, ZN => n141);
   U743 : NAND4_X1 port map( A1 => n143, A2 => n142, A3 => n141, A4 => n140, ZN
                           => n149);
   U744 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n785, B1 => 
                           REGISTERS_15_3_port, B2 => n767, ZN => n147);
   U745 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n821, B1 => 
                           REGISTERS_11_3_port, B2 => n803, ZN => n146);
   U746 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n857, B1 => 
                           REGISTERS_14_3_port, B2 => n839, ZN => n145);
   U747 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n882, B1 => 
                           REGISTERS_10_3_port, B2 => n867, ZN => n144);
   U748 : NAND4_X1 port map( A1 => n147, A2 => n146, A3 => n145, A4 => n144, ZN
                           => n148);
   U749 : AOI22_X1 port map( A1 => n149, A2 => n891, B1 => n148, B2 => n887, ZN
                           => n150);
   U750 : OAI221_X1 port map( B1 => n899, B2 => n152, C1 => n893, C2 => n151, A
                           => n150, ZN => N221);
   U751 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n785, B1 => 
                           REGISTERS_23_4_port, B2 => n767, ZN => n156);
   U752 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n821, B1 => 
                           REGISTERS_19_4_port, B2 => n803, ZN => n155);
   U753 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n857, B1 => 
                           REGISTERS_22_4_port, B2 => n839, ZN => n154);
   U754 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n882, B1 => 
                           REGISTERS_18_4_port, B2 => n867, ZN => n153);
   U755 : AND4_X1 port map( A1 => n156, A2 => n155, A3 => n154, A4 => n153, ZN 
                           => n173);
   U756 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n785, B1 => 
                           REGISTERS_31_4_port, B2 => n767, ZN => n160);
   U757 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n821, B1 => 
                           REGISTERS_27_4_port, B2 => n803, ZN => n159);
   U758 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n857, B1 => 
                           REGISTERS_30_4_port, B2 => n839, ZN => n158);
   U759 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n882, B1 => 
                           REGISTERS_26_4_port, B2 => n867, ZN => n157);
   U760 : AND4_X1 port map( A1 => n160, A2 => n159, A3 => n158, A4 => n157, ZN 
                           => n172);
   U761 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n785, B1 => 
                           REGISTERS_7_4_port, B2 => n767, ZN => n164);
   U762 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n821, B1 => 
                           REGISTERS_3_4_port, B2 => n803, ZN => n163);
   U763 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n857, B1 => 
                           REGISTERS_6_4_port, B2 => n839, ZN => n162);
   U764 : NAND4_X1 port map( A1 => n164, A2 => n163, A3 => n162, A4 => n161, ZN
                           => n170);
   U765 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n785, B1 => 
                           REGISTERS_15_4_port, B2 => n767, ZN => n168);
   U766 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n821, B1 => 
                           REGISTERS_11_4_port, B2 => n803, ZN => n167);
   U767 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n857, B1 => 
                           REGISTERS_14_4_port, B2 => n839, ZN => n166);
   U768 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n882, B1 => 
                           REGISTERS_10_4_port, B2 => n867, ZN => n165);
   U769 : NAND4_X1 port map( A1 => n168, A2 => n167, A3 => n166, A4 => n165, ZN
                           => n169);
   U770 : AOI22_X1 port map( A1 => n170, A2 => n891, B1 => n169, B2 => n887, ZN
                           => n171);
   U771 : OAI221_X1 port map( B1 => n899, B2 => n173, C1 => n893, C2 => n172, A
                           => n171, ZN => N220);
   U772 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n785, B1 => 
                           REGISTERS_23_5_port, B2 => n767, ZN => n177);
   U773 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n821, B1 => 
                           REGISTERS_19_5_port, B2 => n803, ZN => n176);
   U774 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n857, B1 => 
                           REGISTERS_22_5_port, B2 => n839, ZN => n175);
   U775 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n882, B1 => 
                           REGISTERS_18_5_port, B2 => n867, ZN => n174);
   U776 : AND4_X1 port map( A1 => n177, A2 => n176, A3 => n175, A4 => n174, ZN 
                           => n194_port);
   U777 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n785, B1 => 
                           REGISTERS_31_5_port, B2 => n767, ZN => n181);
   U778 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n821, B1 => 
                           REGISTERS_27_5_port, B2 => n803, ZN => n180);
   U779 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n857, B1 => 
                           REGISTERS_30_5_port, B2 => n839, ZN => n179);
   U780 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n882, B1 => 
                           REGISTERS_26_5_port, B2 => n867, ZN => n178);
   U781 : AND4_X1 port map( A1 => n181, A2 => n180, A3 => n179, A4 => n178, ZN 
                           => n193_port);
   U782 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n784, B1 => 
                           REGISTERS_7_5_port, B2 => n766, ZN => n185);
   U783 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n820, B1 => 
                           REGISTERS_3_5_port, B2 => n802, ZN => n184);
   U784 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n856, B1 => 
                           REGISTERS_6_5_port, B2 => n838, ZN => n183);
   U785 : NAND4_X1 port map( A1 => n185, A2 => n184, A3 => n183, A4 => n182, ZN
                           => n191);
   U786 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n784, B1 => 
                           REGISTERS_15_5_port, B2 => n766, ZN => n189);
   U787 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n820, B1 => 
                           REGISTERS_11_5_port, B2 => n802, ZN => n188);
   U788 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n856, B1 => 
                           REGISTERS_14_5_port, B2 => n838, ZN => n187);
   U789 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n882, B1 => 
                           REGISTERS_10_5_port, B2 => n867, ZN => n186);
   U790 : NAND4_X1 port map( A1 => n189, A2 => n188, A3 => n187, A4 => n186, ZN
                           => n190);
   U791 : AOI22_X1 port map( A1 => n191, A2 => n891, B1 => n190, B2 => n887, ZN
                           => n192);
   U792 : OAI221_X1 port map( B1 => n899, B2 => n194_port, C1 => n893, C2 => 
                           n193_port, A => n192, ZN => N219);
   U793 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n784, B1 => 
                           REGISTERS_23_6_port, B2 => n766, ZN => n198_port);
   U794 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n820, B1 => 
                           REGISTERS_19_6_port, B2 => n802, ZN => n197_port);
   U795 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n856, B1 => 
                           REGISTERS_22_6_port, B2 => n838, ZN => n196_port);
   U796 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n882, B1 => 
                           REGISTERS_18_6_port, B2 => n867, ZN => n195_port);
   U797 : AND4_X1 port map( A1 => n198_port, A2 => n197_port, A3 => n196_port, 
                           A4 => n195_port, ZN => n215_port);
   U798 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n784, B1 => 
                           REGISTERS_31_6_port, B2 => n766, ZN => n202_port);
   U799 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n820, B1 => 
                           REGISTERS_27_6_port, B2 => n802, ZN => n201_port);
   U800 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n856, B1 => 
                           REGISTERS_30_6_port, B2 => n838, ZN => n200_port);
   U801 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n882, B1 => 
                           REGISTERS_26_6_port, B2 => n867, ZN => n199_port);
   U802 : AND4_X1 port map( A1 => n202_port, A2 => n201_port, A3 => n200_port, 
                           A4 => n199_port, ZN => n214_port);
   U803 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n784, B1 => 
                           REGISTERS_7_6_port, B2 => n766, ZN => n206_port);
   U804 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n820, B1 => 
                           REGISTERS_3_6_port, B2 => n802, ZN => n205_port);
   U805 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n856, B1 => 
                           REGISTERS_6_6_port, B2 => n838, ZN => n204_port);
   U806 : NAND4_X1 port map( A1 => n206_port, A2 => n205_port, A3 => n204_port,
                           A4 => n203_port, ZN => n212_port);
   U807 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n784, B1 => 
                           REGISTERS_15_6_port, B2 => n766, ZN => n210_port);
   U808 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n820, B1 => 
                           REGISTERS_11_6_port, B2 => n802, ZN => n209_port);
   U809 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n856, B1 => 
                           REGISTERS_14_6_port, B2 => n838, ZN => n208_port);
   U810 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n882, B1 => 
                           REGISTERS_10_6_port, B2 => n867, ZN => n207_port);
   U811 : NAND4_X1 port map( A1 => n210_port, A2 => n209_port, A3 => n208_port,
                           A4 => n207_port, ZN => n211_port);
   U812 : AOI22_X1 port map( A1 => n212_port, A2 => n891, B1 => n211_port, B2 
                           => n887, ZN => n213_port);
   U813 : OAI221_X1 port map( B1 => n899, B2 => n215_port, C1 => n893, C2 => 
                           n214_port, A => n213_port, ZN => N218);
   U814 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n784, B1 => 
                           REGISTERS_23_7_port, B2 => n766, ZN => n219_port);
   U815 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n820, B1 => 
                           REGISTERS_19_7_port, B2 => n802, ZN => n218_port);
   U816 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n856, B1 => 
                           REGISTERS_22_7_port, B2 => n838, ZN => n217_port);
   U817 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n882, B1 => 
                           REGISTERS_18_7_port, B2 => n867, ZN => n216_port);
   U818 : AND4_X1 port map( A1 => n219_port, A2 => n218_port, A3 => n217_port, 
                           A4 => n216_port, ZN => n236_port);
   U819 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n784, B1 => 
                           REGISTERS_31_7_port, B2 => n766, ZN => n223_port);
   U820 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n820, B1 => 
                           REGISTERS_27_7_port, B2 => n802, ZN => n222_port);
   U821 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n856, B1 => 
                           REGISTERS_30_7_port, B2 => n838, ZN => n221_port);
   U822 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n881, B1 => 
                           REGISTERS_26_7_port, B2 => n867, ZN => n220_port);
   U823 : AND4_X1 port map( A1 => n223_port, A2 => n222_port, A3 => n221_port, 
                           A4 => n220_port, ZN => n235_port);
   U824 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n784, B1 => 
                           REGISTERS_7_7_port, B2 => n766, ZN => n227_port);
   U825 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n820, B1 => 
                           REGISTERS_3_7_port, B2 => n802, ZN => n226_port);
   U826 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n856, B1 => 
                           REGISTERS_6_7_port, B2 => n838, ZN => n225_port);
   U827 : NAND4_X1 port map( A1 => n227_port, A2 => n226_port, A3 => n225_port,
                           A4 => n224_port, ZN => n233_port);
   U828 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n784, B1 => 
                           REGISTERS_15_7_port, B2 => n766, ZN => n231_port);
   U829 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n820, B1 => 
                           REGISTERS_11_7_port, B2 => n802, ZN => n230_port);
   U830 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n856, B1 => 
                           REGISTERS_14_7_port, B2 => n838, ZN => n229_port);
   U831 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n881, B1 => 
                           REGISTERS_10_7_port, B2 => n867, ZN => n228_port);
   U832 : NAND4_X1 port map( A1 => n231_port, A2 => n230_port, A3 => n229_port,
                           A4 => n228_port, ZN => n232_port);
   U833 : AOI22_X1 port map( A1 => n233_port, A2 => n891, B1 => n232_port, B2 
                           => n887, ZN => n234_port);
   U834 : OAI221_X1 port map( B1 => n899, B2 => n236_port, C1 => n893, C2 => 
                           n235_port, A => n234_port, ZN => N217);
   U835 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n784, B1 => 
                           REGISTERS_23_8_port, B2 => n766, ZN => n240_port);
   U836 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n820, B1 => 
                           REGISTERS_19_8_port, B2 => n802, ZN => n239_port);
   U837 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n856, B1 => 
                           REGISTERS_22_8_port, B2 => n838, ZN => n238_port);
   U838 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n881, B1 => 
                           REGISTERS_18_8_port, B2 => n867, ZN => n237_port);
   U839 : AND4_X1 port map( A1 => n240_port, A2 => n239_port, A3 => n238_port, 
                           A4 => n237_port, ZN => n257);
   U840 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n783, B1 => 
                           REGISTERS_31_8_port, B2 => n765, ZN => n244_port);
   U841 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n819, B1 => 
                           REGISTERS_27_8_port, B2 => n801, ZN => n243_port);
   U842 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n855, B1 => 
                           REGISTERS_30_8_port, B2 => n837, ZN => n242_port);
   U843 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n881, B1 => 
                           REGISTERS_26_8_port, B2 => n867, ZN => n241_port);
   U844 : AND4_X1 port map( A1 => n244_port, A2 => n243_port, A3 => n242_port, 
                           A4 => n241_port, ZN => n256_port);
   U845 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n783, B1 => 
                           REGISTERS_7_8_port, B2 => n765, ZN => n248_port);
   U846 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n819, B1 => 
                           REGISTERS_3_8_port, B2 => n801, ZN => n247_port);
   U847 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n855, B1 => 
                           REGISTERS_6_8_port, B2 => n837, ZN => n246_port);
   U848 : NAND4_X1 port map( A1 => n248_port, A2 => n247_port, A3 => n246_port,
                           A4 => n245_port, ZN => n254_port);
   U849 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n783, B1 => 
                           REGISTERS_15_8_port, B2 => n765, ZN => n252_port);
   U850 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n819, B1 => 
                           REGISTERS_11_8_port, B2 => n801, ZN => n251_port);
   U851 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n855, B1 => 
                           REGISTERS_14_8_port, B2 => n837, ZN => n250_port);
   U852 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n881, B1 => 
                           REGISTERS_10_8_port, B2 => n866, ZN => n249_port);
   U853 : NAND4_X1 port map( A1 => n252_port, A2 => n251_port, A3 => n250_port,
                           A4 => n249_port, ZN => n253_port);
   U854 : AOI22_X1 port map( A1 => n254_port, A2 => n891, B1 => n253_port, B2 
                           => n887, ZN => n255_port);
   U855 : OAI221_X1 port map( B1 => n899, B2 => n257, C1 => n893, C2 => 
                           n256_port, A => n255_port, ZN => N216);
   U856 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n783, B1 => 
                           REGISTERS_23_9_port, B2 => n765, ZN => n261_port);
   U857 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n819, B1 => 
                           REGISTERS_19_9_port, B2 => n801, ZN => n260_port);
   U858 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n855, B1 => 
                           REGISTERS_22_9_port, B2 => n837, ZN => n259_port);
   U859 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n881, B1 => 
                           REGISTERS_18_9_port, B2 => n866, ZN => n258);
   U860 : AND4_X1 port map( A1 => n261_port, A2 => n260_port, A3 => n259_port, 
                           A4 => n258, ZN => n278_port);
   U861 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n783, B1 => 
                           REGISTERS_31_9_port, B2 => n765, ZN => n265_port);
   U862 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n819, B1 => 
                           REGISTERS_27_9_port, B2 => n801, ZN => n264_port);
   U863 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n855, B1 => 
                           REGISTERS_30_9_port, B2 => n837, ZN => n263_port);
   U864 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n881, B1 => 
                           REGISTERS_26_9_port, B2 => n866, ZN => n262_port);
   U865 : AND4_X1 port map( A1 => n265_port, A2 => n264_port, A3 => n263_port, 
                           A4 => n262_port, ZN => n277_port);
   U866 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n783, B1 => 
                           REGISTERS_7_9_port, B2 => n765, ZN => n269_port);
   U867 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n819, B1 => 
                           REGISTERS_3_9_port, B2 => n801, ZN => n268_port);
   U868 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n855, B1 => 
                           REGISTERS_6_9_port, B2 => n837, ZN => n267_port);
   U869 : NAND4_X1 port map( A1 => n269_port, A2 => n268_port, A3 => n267_port,
                           A4 => n266_port, ZN => n275_port);
   U870 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n783, B1 => 
                           REGISTERS_15_9_port, B2 => n765, ZN => n273_port);
   U871 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n819, B1 => 
                           REGISTERS_11_9_port, B2 => n801, ZN => n272_port);
   U872 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n855, B1 => 
                           REGISTERS_14_9_port, B2 => n837, ZN => n271_port);
   U873 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n881, B1 => 
                           REGISTERS_10_9_port, B2 => n866, ZN => n270_port);
   U874 : NAND4_X1 port map( A1 => n273_port, A2 => n272_port, A3 => n271_port,
                           A4 => n270_port, ZN => n274_port);
   U875 : AOI22_X1 port map( A1 => n275_port, A2 => n891, B1 => n274_port, B2 
                           => n887, ZN => n276_port);
   U876 : OAI221_X1 port map( B1 => n899, B2 => n278_port, C1 => n893, C2 => 
                           n277_port, A => n276_port, ZN => N215);
   U877 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n783, B1 => 
                           REGISTERS_23_10_port, B2 => n765, ZN => n282_port);
   U878 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n819, B1 => 
                           REGISTERS_19_10_port, B2 => n801, ZN => n281_port);
   U879 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n855, B1 => 
                           REGISTERS_22_10_port, B2 => n837, ZN => n280_port);
   U880 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n881, B1 => 
                           REGISTERS_18_10_port, B2 => n866, ZN => n279_port);
   U881 : AND4_X1 port map( A1 => n282_port, A2 => n281_port, A3 => n280_port, 
                           A4 => n279_port, ZN => n299_port);
   U882 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n783, B1 => 
                           REGISTERS_31_10_port, B2 => n765, ZN => n286_port);
   U883 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n819, B1 => 
                           REGISTERS_27_10_port, B2 => n801, ZN => n285_port);
   U884 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n855, B1 => 
                           REGISTERS_30_10_port, B2 => n837, ZN => n284_port);
   U885 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n881, B1 => 
                           REGISTERS_26_10_port, B2 => n866, ZN => n283_port);
   U886 : AND4_X1 port map( A1 => n286_port, A2 => n285_port, A3 => n284_port, 
                           A4 => n283_port, ZN => n298_port);
   U887 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n783, B1 => 
                           REGISTERS_7_10_port, B2 => n765, ZN => n290_port);
   U888 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n819, B1 => 
                           REGISTERS_3_10_port, B2 => n801, ZN => n289_port);
   U889 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n855, B1 => 
                           REGISTERS_6_10_port, B2 => n837, ZN => n288_port);
   U890 : NAND4_X1 port map( A1 => n290_port, A2 => n289_port, A3 => n288_port,
                           A4 => n287_port, ZN => n296_port);
   U891 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n783, B1 => 
                           REGISTERS_15_10_port, B2 => n765, ZN => n294_port);
   U892 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n819, B1 => 
                           REGISTERS_11_10_port, B2 => n801, ZN => n293_port);
   U893 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n855, B1 => 
                           REGISTERS_14_10_port, B2 => n837, ZN => n292_port);
   U894 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n881, B1 => 
                           REGISTERS_10_10_port, B2 => n866, ZN => n291_port);
   U895 : NAND4_X1 port map( A1 => n294_port, A2 => n293_port, A3 => n292_port,
                           A4 => n291_port, ZN => n295_port);
   U896 : AOI22_X1 port map( A1 => n296_port, A2 => n891, B1 => n295_port, B2 
                           => n887, ZN => n297_port);
   U897 : OAI221_X1 port map( B1 => n899, B2 => n299_port, C1 => n894, C2 => 
                           n298_port, A => n297_port, ZN => N214);
   U898 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n782, B1 => 
                           REGISTERS_23_11_port, B2 => n764, ZN => n303_port);
   U899 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n818, B1 => 
                           REGISTERS_19_11_port, B2 => n800, ZN => n302_port);
   U900 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n854, B1 => 
                           REGISTERS_22_11_port, B2 => n836, ZN => n301_port);
   U901 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n880, B1 => 
                           REGISTERS_18_11_port, B2 => n866, ZN => n300_port);
   U902 : AND4_X1 port map( A1 => n303_port, A2 => n302_port, A3 => n301_port, 
                           A4 => n300_port, ZN => n320_port);
   U903 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n782, B1 => 
                           REGISTERS_31_11_port, B2 => n764, ZN => n307_port);
   U904 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n818, B1 => 
                           REGISTERS_27_11_port, B2 => n800, ZN => n306_port);
   U905 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n854, B1 => 
                           REGISTERS_30_11_port, B2 => n836, ZN => n305_port);
   U906 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n880, B1 => 
                           REGISTERS_26_11_port, B2 => n866, ZN => n304_port);
   U907 : AND4_X1 port map( A1 => n307_port, A2 => n306_port, A3 => n305_port, 
                           A4 => n304_port, ZN => n319_port);
   U908 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n782, B1 => 
                           REGISTERS_7_11_port, B2 => n764, ZN => n311_port);
   U909 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n818, B1 => 
                           REGISTERS_3_11_port, B2 => n800, ZN => n310_port);
   U910 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n854, B1 => 
                           REGISTERS_6_11_port, B2 => n836, ZN => n309_port);
   U911 : NAND4_X1 port map( A1 => n311_port, A2 => n310_port, A3 => n309_port,
                           A4 => n308_port, ZN => n317_port);
   U912 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n782, B1 => 
                           REGISTERS_15_11_port, B2 => n764, ZN => n315_port);
   U913 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n818, B1 => 
                           REGISTERS_11_11_port, B2 => n800, ZN => n314_port);
   U914 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n854, B1 => 
                           REGISTERS_14_11_port, B2 => n836, ZN => n313_port);
   U915 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n880, B1 => 
                           REGISTERS_10_11_port, B2 => n866, ZN => n312_port);
   U916 : NAND4_X1 port map( A1 => n315_port, A2 => n314_port, A3 => n313_port,
                           A4 => n312_port, ZN => n316_port);
   U917 : AOI22_X1 port map( A1 => n317_port, A2 => n890, B1 => n316_port, B2 
                           => n886, ZN => n318_port);
   U918 : OAI221_X1 port map( B1 => n898, B2 => n320_port, C1 => n894, C2 => 
                           n319_port, A => n318_port, ZN => N213);
   U919 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n782, B1 => 
                           REGISTERS_23_12_port, B2 => n764, ZN => n324_port);
   U920 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n818, B1 => 
                           REGISTERS_19_12_port, B2 => n800, ZN => n323_port);
   U921 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n854, B1 => 
                           REGISTERS_22_12_port, B2 => n836, ZN => n322_port);
   U922 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n880, B1 => 
                           REGISTERS_18_12_port, B2 => n866, ZN => n321_port);
   U923 : AND4_X1 port map( A1 => n324_port, A2 => n323_port, A3 => n322_port, 
                           A4 => n321_port, ZN => n341_port);
   U924 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n782, B1 => 
                           REGISTERS_31_12_port, B2 => n764, ZN => n328_port);
   U925 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n818, B1 => 
                           REGISTERS_27_12_port, B2 => n800, ZN => n327_port);
   U926 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n854, B1 => 
                           REGISTERS_30_12_port, B2 => n836, ZN => n326_port);
   U927 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n880, B1 => 
                           REGISTERS_26_12_port, B2 => n866, ZN => n325_port);
   U928 : AND4_X1 port map( A1 => n328_port, A2 => n327_port, A3 => n326_port, 
                           A4 => n325_port, ZN => n340_port);
   U929 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n782, B1 => 
                           REGISTERS_7_12_port, B2 => n764, ZN => n332_port);
   U930 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n818, B1 => 
                           REGISTERS_3_12_port, B2 => n800, ZN => n331_port);
   U931 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n854, B1 => 
                           REGISTERS_6_12_port, B2 => n836, ZN => n330_port);
   U932 : NAND4_X1 port map( A1 => n332_port, A2 => n331_port, A3 => n330_port,
                           A4 => n329_port, ZN => n338_port);
   U933 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n782, B1 => 
                           REGISTERS_15_12_port, B2 => n764, ZN => n336_port);
   U934 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n818, B1 => 
                           REGISTERS_11_12_port, B2 => n800, ZN => n335_port);
   U935 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n854, B1 => 
                           REGISTERS_14_12_port, B2 => n836, ZN => n334_port);
   U936 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n880, B1 => 
                           REGISTERS_10_12_port, B2 => n866, ZN => n333_port);
   U937 : NAND4_X1 port map( A1 => n336_port, A2 => n335_port, A3 => n334_port,
                           A4 => n333_port, ZN => n337_port);
   U938 : AOI22_X1 port map( A1 => n338_port, A2 => n890, B1 => n337_port, B2 
                           => n886, ZN => n339_port);
   U939 : OAI221_X1 port map( B1 => n898, B2 => n341_port, C1 => n894, C2 => 
                           n340_port, A => n339_port, ZN => N212);
   U940 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n782, B1 => 
                           REGISTERS_23_13_port, B2 => n764, ZN => n345_port);
   U941 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n818, B1 => 
                           REGISTERS_19_13_port, B2 => n800, ZN => n344_port);
   U942 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n854, B1 => 
                           REGISTERS_22_13_port, B2 => n836, ZN => n343_port);
   U943 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n880, B1 => 
                           REGISTERS_18_13_port, B2 => n866, ZN => n342_port);
   U944 : AND4_X1 port map( A1 => n345_port, A2 => n344_port, A3 => n343_port, 
                           A4 => n342_port, ZN => n362);
   U945 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n782, B1 => 
                           REGISTERS_31_13_port, B2 => n764, ZN => n349_port);
   U946 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n818, B1 => 
                           REGISTERS_27_13_port, B2 => n800, ZN => n348_port);
   U947 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n854, B1 => 
                           REGISTERS_30_13_port, B2 => n836, ZN => n347_port);
   U948 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n880, B1 => 
                           REGISTERS_26_13_port, B2 => n866, ZN => n346_port);
   U949 : AND4_X1 port map( A1 => n349_port, A2 => n348_port, A3 => n347_port, 
                           A4 => n346_port, ZN => n361);
   U950 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n782, B1 => 
                           REGISTERS_7_13_port, B2 => n764, ZN => n353_port);
   U951 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n818, B1 => 
                           REGISTERS_3_13_port, B2 => n800, ZN => n352_port);
   U952 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n854, B1 => 
                           REGISTERS_6_13_port, B2 => n836, ZN => n351_port);
   U953 : NAND4_X1 port map( A1 => n353_port, A2 => n352_port, A3 => n351_port,
                           A4 => n350_port, ZN => n359);
   U954 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n781, B1 => 
                           REGISTERS_15_13_port, B2 => n763, ZN => n357);
   U955 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n817, B1 => 
                           REGISTERS_11_13_port, B2 => n799, ZN => n356);
   U956 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n853, B1 => 
                           REGISTERS_14_13_port, B2 => n835, ZN => n355);
   U957 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n880, B1 => 
                           REGISTERS_10_13_port, B2 => n866, ZN => n354);
   U958 : NAND4_X1 port map( A1 => n357, A2 => n356, A3 => n355, A4 => n354, ZN
                           => n358);
   U959 : AOI22_X1 port map( A1 => n359, A2 => n890, B1 => n358, B2 => n886, ZN
                           => n360);
   U960 : OAI221_X1 port map( B1 => n898, B2 => n362, C1 => n894, C2 => n361, A
                           => n360, ZN => N211);
   U961 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n781, B1 => 
                           REGISTERS_23_14_port, B2 => n763, ZN => n366);
   U962 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n817, B1 => 
                           REGISTERS_19_14_port, B2 => n799, ZN => n365);
   U963 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n853, B1 => 
                           REGISTERS_22_14_port, B2 => n835, ZN => n364);
   U964 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n880, B1 => 
                           REGISTERS_18_14_port, B2 => n866, ZN => n363);
   U965 : AND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN 
                           => n383);
   U966 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n781, B1 => 
                           REGISTERS_31_14_port, B2 => n763, ZN => n370);
   U967 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n817, B1 => 
                           REGISTERS_27_14_port, B2 => n799, ZN => n369);
   U968 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n853, B1 => 
                           REGISTERS_30_14_port, B2 => n835, ZN => n368);
   U969 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n880, B1 => 
                           REGISTERS_26_14_port, B2 => n866, ZN => n367);
   U970 : AND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN 
                           => n382);
   U971 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n781, B1 => 
                           REGISTERS_7_14_port, B2 => n763, ZN => n374);
   U972 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n817, B1 => 
                           REGISTERS_3_14_port, B2 => n799, ZN => n373);
   U973 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n853, B1 => 
                           REGISTERS_6_14_port, B2 => n835, ZN => n372);
   U974 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => n380);
   U975 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n781, B1 => 
                           REGISTERS_15_14_port, B2 => n763, ZN => n378);
   U976 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n817, B1 => 
                           REGISTERS_11_14_port, B2 => n799, ZN => n377);
   U977 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n853, B1 => 
                           REGISTERS_14_14_port, B2 => n835, ZN => n376);
   U978 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n879, B1 => 
                           REGISTERS_10_14_port, B2 => n866, ZN => n375);
   U979 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => n379);
   U980 : AOI22_X1 port map( A1 => n380, A2 => n890, B1 => n379, B2 => n886, ZN
                           => n381);
   U981 : OAI221_X1 port map( B1 => n898, B2 => n383, C1 => n894, C2 => n382, A
                           => n381, ZN => N210);
   U982 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n781, B1 => 
                           REGISTERS_23_15_port, B2 => n763, ZN => n387);
   U983 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n817, B1 => 
                           REGISTERS_19_15_port, B2 => n799, ZN => n386);
   U984 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n853, B1 => 
                           REGISTERS_22_15_port, B2 => n835, ZN => n385);
   U985 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n879, B1 => 
                           REGISTERS_18_15_port, B2 => n866, ZN => n384);
   U986 : AND4_X1 port map( A1 => n387, A2 => n386, A3 => n385, A4 => n384, ZN 
                           => n404);
   U987 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n781, B1 => 
                           REGISTERS_31_15_port, B2 => n763, ZN => n391);
   U988 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n817, B1 => 
                           REGISTERS_27_15_port, B2 => n799, ZN => n390);
   U989 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n853, B1 => 
                           REGISTERS_30_15_port, B2 => n835, ZN => n389);
   U990 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n879, B1 => 
                           REGISTERS_26_15_port, B2 => n865, ZN => n388);
   U991 : AND4_X1 port map( A1 => n391, A2 => n390, A3 => n389, A4 => n388, ZN 
                           => n403);
   U992 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n781, B1 => 
                           REGISTERS_7_15_port, B2 => n763, ZN => n395);
   U993 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n817, B1 => 
                           REGISTERS_3_15_port, B2 => n799, ZN => n394);
   U994 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n853, B1 => 
                           REGISTERS_6_15_port, B2 => n835, ZN => n393);
   U995 : NAND4_X1 port map( A1 => n395, A2 => n394, A3 => n393, A4 => n392, ZN
                           => n401);
   U996 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n781, B1 => 
                           REGISTERS_15_15_port, B2 => n763, ZN => n399);
   U997 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n817, B1 => 
                           REGISTERS_11_15_port, B2 => n799, ZN => n398);
   U998 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n853, B1 => 
                           REGISTERS_14_15_port, B2 => n835, ZN => n397);
   U999 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n879, B1 => 
                           REGISTERS_10_15_port, B2 => n865, ZN => n396);
   U1000 : NAND4_X1 port map( A1 => n399, A2 => n398, A3 => n397, A4 => n396, 
                           ZN => n400);
   U1001 : AOI22_X1 port map( A1 => n401, A2 => n890, B1 => n400, B2 => n886, 
                           ZN => n402);
   U1002 : OAI221_X1 port map( B1 => n898, B2 => n404, C1 => n894, C2 => n403, 
                           A => n402, ZN => N209);
   U1003 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n781, B1 => 
                           REGISTERS_23_16_port, B2 => n763, ZN => n408);
   U1004 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n817, B1 => 
                           REGISTERS_19_16_port, B2 => n799, ZN => n407);
   U1005 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n853, B1 => 
                           REGISTERS_22_16_port, B2 => n835, ZN => n406);
   U1006 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n879, B1 => 
                           REGISTERS_18_16_port, B2 => n865, ZN => n405);
   U1007 : AND4_X1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, ZN
                           => n425);
   U1008 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n781, B1 => 
                           REGISTERS_31_16_port, B2 => n763, ZN => n412);
   U1009 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n817, B1 => 
                           REGISTERS_27_16_port, B2 => n799, ZN => n411);
   U1010 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n853, B1 => 
                           REGISTERS_30_16_port, B2 => n835, ZN => n410);
   U1011 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n879, B1 => 
                           REGISTERS_26_16_port, B2 => n865, ZN => n409);
   U1012 : AND4_X1 port map( A1 => n412, A2 => n411, A3 => n410, A4 => n409, ZN
                           => n424);
   U1013 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n780, B1 => 
                           REGISTERS_7_16_port, B2 => n762, ZN => n416);
   U1014 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n816, B1 => 
                           REGISTERS_3_16_port, B2 => n798, ZN => n415);
   U1015 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n852, B1 => 
                           REGISTERS_6_16_port, B2 => n834, ZN => n414);
   U1016 : NAND4_X1 port map( A1 => n416, A2 => n415, A3 => n414, A4 => n413, 
                           ZN => n422);
   U1017 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n780, B1 => 
                           REGISTERS_15_16_port, B2 => n762, ZN => n420);
   U1018 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n816, B1 => 
                           REGISTERS_11_16_port, B2 => n798, ZN => n419);
   U1019 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n852, B1 => 
                           REGISTERS_14_16_port, B2 => n834, ZN => n418);
   U1020 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n879, B1 => 
                           REGISTERS_10_16_port, B2 => n865, ZN => n417);
   U1021 : NAND4_X1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, 
                           ZN => n421);
   U1022 : AOI22_X1 port map( A1 => n422, A2 => n890, B1 => n421, B2 => n886, 
                           ZN => n423);
   U1023 : OAI221_X1 port map( B1 => n898, B2 => n425, C1 => n894, C2 => n424, 
                           A => n423, ZN => N208);
   U1024 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n780, B1 => 
                           REGISTERS_23_17_port, B2 => n762, ZN => n429);
   U1025 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n816, B1 => 
                           REGISTERS_19_17_port, B2 => n798, ZN => n428);
   U1026 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n852, B1 => 
                           REGISTERS_22_17_port, B2 => n834, ZN => n427);
   U1027 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n879, B1 => 
                           REGISTERS_18_17_port, B2 => n865, ZN => n426);
   U1028 : AND4_X1 port map( A1 => n429, A2 => n428, A3 => n427, A4 => n426, ZN
                           => n446);
   U1029 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n780, B1 => 
                           REGISTERS_31_17_port, B2 => n762, ZN => n433);
   U1030 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n816, B1 => 
                           REGISTERS_27_17_port, B2 => n798, ZN => n432);
   U1031 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n852, B1 => 
                           REGISTERS_30_17_port, B2 => n834, ZN => n431);
   U1032 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n879, B1 => 
                           REGISTERS_26_17_port, B2 => n865, ZN => n430);
   U1033 : AND4_X1 port map( A1 => n433, A2 => n432, A3 => n431, A4 => n430, ZN
                           => n445);
   U1034 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n780, B1 => 
                           REGISTERS_7_17_port, B2 => n762, ZN => n437);
   U1035 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n816, B1 => 
                           REGISTERS_3_17_port, B2 => n798, ZN => n436);
   U1036 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n852, B1 => 
                           REGISTERS_6_17_port, B2 => n834, ZN => n435);
   U1037 : NAND4_X1 port map( A1 => n437, A2 => n436, A3 => n435, A4 => n434, 
                           ZN => n443);
   U1038 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n780, B1 => 
                           REGISTERS_15_17_port, B2 => n762, ZN => n441);
   U1039 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n816, B1 => 
                           REGISTERS_11_17_port, B2 => n798, ZN => n440);
   U1040 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n852, B1 => 
                           REGISTERS_14_17_port, B2 => n834, ZN => n439);
   U1041 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n879, B1 => 
                           REGISTERS_10_17_port, B2 => n865, ZN => n438);
   U1042 : NAND4_X1 port map( A1 => n441, A2 => n440, A3 => n439, A4 => n438, 
                           ZN => n442);
   U1043 : AOI22_X1 port map( A1 => n443, A2 => n890, B1 => n442, B2 => n886, 
                           ZN => n444);
   U1044 : OAI221_X1 port map( B1 => n898, B2 => n446, C1 => n894, C2 => n445, 
                           A => n444, ZN => N207);
   U1045 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n780, B1 => 
                           REGISTERS_23_18_port, B2 => n762, ZN => n450);
   U1046 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n816, B1 => 
                           REGISTERS_19_18_port, B2 => n798, ZN => n449);
   U1047 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n852, B1 => 
                           REGISTERS_22_18_port, B2 => n834, ZN => n448);
   U1048 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n879, B1 => 
                           REGISTERS_18_18_port, B2 => n865, ZN => n447);
   U1049 : AND4_X1 port map( A1 => n450, A2 => n449, A3 => n448, A4 => n447, ZN
                           => n467);
   U1050 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n780, B1 => 
                           REGISTERS_31_18_port, B2 => n762, ZN => n454);
   U1051 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n816, B1 => 
                           REGISTERS_27_18_port, B2 => n798, ZN => n453);
   U1052 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n852, B1 => 
                           REGISTERS_30_18_port, B2 => n834, ZN => n452);
   U1053 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n878, B1 => 
                           REGISTERS_26_18_port, B2 => n865, ZN => n451);
   U1054 : AND4_X1 port map( A1 => n454, A2 => n453, A3 => n452, A4 => n451, ZN
                           => n466);
   U1055 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n780, B1 => 
                           REGISTERS_7_18_port, B2 => n762, ZN => n458);
   U1056 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n816, B1 => 
                           REGISTERS_3_18_port, B2 => n798, ZN => n457);
   U1057 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n852, B1 => 
                           REGISTERS_6_18_port, B2 => n834, ZN => n456);
   U1058 : NAND4_X1 port map( A1 => n458, A2 => n457, A3 => n456, A4 => n455, 
                           ZN => n464);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n780, B1 => 
                           REGISTERS_15_18_port, B2 => n762, ZN => n462);
   U1060 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n816, B1 => 
                           REGISTERS_11_18_port, B2 => n798, ZN => n461);
   U1061 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n852, B1 => 
                           REGISTERS_14_18_port, B2 => n834, ZN => n460);
   U1062 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n878, B1 => 
                           REGISTERS_10_18_port, B2 => n865, ZN => n459);
   U1063 : NAND4_X1 port map( A1 => n462, A2 => n461, A3 => n460, A4 => n459, 
                           ZN => n463);
   U1064 : AOI22_X1 port map( A1 => n464, A2 => n890, B1 => n463, B2 => n886, 
                           ZN => n465);
   U1065 : OAI221_X1 port map( B1 => n898, B2 => n467, C1 => n894, C2 => n466, 
                           A => n465, ZN => N206);
   U1066 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n780, B1 => 
                           REGISTERS_23_19_port, B2 => n762, ZN => n471);
   U1067 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n816, B1 => 
                           REGISTERS_19_19_port, B2 => n798, ZN => n470);
   U1068 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n852, B1 => 
                           REGISTERS_22_19_port, B2 => n834, ZN => n469);
   U1069 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n878, B1 => 
                           REGISTERS_18_19_port, B2 => n865, ZN => n468);
   U1070 : AND4_X1 port map( A1 => n471, A2 => n470, A3 => n469, A4 => n468, ZN
                           => n488);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n779, B1 => 
                           REGISTERS_31_19_port, B2 => n761, ZN => n475);
   U1072 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n815, B1 => 
                           REGISTERS_27_19_port, B2 => n797, ZN => n474);
   U1073 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n851, B1 => 
                           REGISTERS_30_19_port, B2 => n833, ZN => n473);
   U1074 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n878, B1 => 
                           REGISTERS_26_19_port, B2 => n865, ZN => n472);
   U1075 : AND4_X1 port map( A1 => n475, A2 => n474, A3 => n473, A4 => n472, ZN
                           => n487);
   U1076 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n779, B1 => 
                           REGISTERS_7_19_port, B2 => n761, ZN => n479);
   U1077 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n815, B1 => 
                           REGISTERS_3_19_port, B2 => n797, ZN => n478);
   U1078 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n851, B1 => 
                           REGISTERS_6_19_port, B2 => n833, ZN => n477);
   U1079 : NAND4_X1 port map( A1 => n479, A2 => n478, A3 => n477, A4 => n476, 
                           ZN => n485);
   U1080 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n779, B1 => 
                           REGISTERS_15_19_port, B2 => n761, ZN => n483);
   U1081 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n815, B1 => 
                           REGISTERS_11_19_port, B2 => n797, ZN => n482);
   U1082 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n851, B1 => 
                           REGISTERS_14_19_port, B2 => n833, ZN => n481);
   U1083 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n878, B1 => 
                           REGISTERS_10_19_port, B2 => n865, ZN => n480);
   U1084 : NAND4_X1 port map( A1 => n483, A2 => n482, A3 => n481, A4 => n480, 
                           ZN => n484);
   U1085 : AOI22_X1 port map( A1 => n485, A2 => n890, B1 => n484, B2 => n886, 
                           ZN => n486);
   U1086 : OAI221_X1 port map( B1 => n898, B2 => n488, C1 => n894, C2 => n487, 
                           A => n486, ZN => N205);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n779, B1 => 
                           REGISTERS_23_20_port, B2 => n761, ZN => n492);
   U1088 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n815, B1 => 
                           REGISTERS_19_20_port, B2 => n797, ZN => n491);
   U1089 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n851, B1 => 
                           REGISTERS_22_20_port, B2 => n833, ZN => n490);
   U1090 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n878, B1 => 
                           REGISTERS_18_20_port, B2 => n865, ZN => n489);
   U1091 : AND4_X1 port map( A1 => n492, A2 => n491, A3 => n490, A4 => n489, ZN
                           => n509);
   U1092 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n779, B1 => 
                           REGISTERS_31_20_port, B2 => n761, ZN => n496);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n815, B1 => 
                           REGISTERS_27_20_port, B2 => n797, ZN => n495);
   U1094 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n851, B1 => 
                           REGISTERS_30_20_port, B2 => n833, ZN => n494);
   U1095 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n878, B1 => 
                           REGISTERS_26_20_port, B2 => n865, ZN => n493);
   U1096 : AND4_X1 port map( A1 => n496, A2 => n495, A3 => n494, A4 => n493, ZN
                           => n508);
   U1097 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n779, B1 => 
                           REGISTERS_7_20_port, B2 => n761, ZN => n500);
   U1098 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n815, B1 => 
                           REGISTERS_3_20_port, B2 => n797, ZN => n499);
   U1099 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n851, B1 => 
                           REGISTERS_6_20_port, B2 => n833, ZN => n498);
   U1100 : NAND4_X1 port map( A1 => n500, A2 => n499, A3 => n498, A4 => n497, 
                           ZN => n506);
   U1101 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n779, B1 => 
                           REGISTERS_15_20_port, B2 => n761, ZN => n504);
   U1102 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n815, B1 => 
                           REGISTERS_11_20_port, B2 => n797, ZN => n503);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n851, B1 => 
                           REGISTERS_14_20_port, B2 => n833, ZN => n502);
   U1104 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n878, B1 => 
                           REGISTERS_10_20_port, B2 => n865, ZN => n501);
   U1105 : NAND4_X1 port map( A1 => n504, A2 => n503, A3 => n502, A4 => n501, 
                           ZN => n505);
   U1106 : AOI22_X1 port map( A1 => n506, A2 => n890, B1 => n505, B2 => n886, 
                           ZN => n507);
   U1107 : OAI221_X1 port map( B1 => n898, B2 => n509, C1 => n894, C2 => n508, 
                           A => n507, ZN => N204);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n779, B1 => 
                           REGISTERS_23_21_port, B2 => n761, ZN => n513);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n815, B1 => 
                           REGISTERS_19_21_port, B2 => n797, ZN => n512);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n851, B1 => 
                           REGISTERS_22_21_port, B2 => n833, ZN => n511);
   U1111 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n878, B1 => 
                           REGISTERS_18_21_port, B2 => n865, ZN => n510);
   U1112 : AND4_X1 port map( A1 => n513, A2 => n512, A3 => n511, A4 => n510, ZN
                           => n530);
   U1113 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n779, B1 => 
                           REGISTERS_31_21_port, B2 => n761, ZN => n517);
   U1114 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n815, B1 => 
                           REGISTERS_27_21_port, B2 => n797, ZN => n516);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n851, B1 => 
                           REGISTERS_30_21_port, B2 => n833, ZN => n515);
   U1116 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n878, B1 => 
                           REGISTERS_26_21_port, B2 => n865, ZN => n514);
   U1117 : AND4_X1 port map( A1 => n517, A2 => n516, A3 => n515, A4 => n514, ZN
                           => n529);
   U1118 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n779, B1 => 
                           REGISTERS_7_21_port, B2 => n761, ZN => n521);
   U1119 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n815, B1 => 
                           REGISTERS_3_21_port, B2 => n797, ZN => n520);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n851, B1 => 
                           REGISTERS_6_21_port, B2 => n833, ZN => n519);
   U1121 : NAND4_X1 port map( A1 => n521, A2 => n520, A3 => n519, A4 => n518, 
                           ZN => n527);
   U1122 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n779, B1 => 
                           REGISTERS_15_21_port, B2 => n761, ZN => n525);
   U1123 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n815, B1 => 
                           REGISTERS_11_21_port, B2 => n797, ZN => n524);
   U1124 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n851, B1 => 
                           REGISTERS_14_21_port, B2 => n833, ZN => n523);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n878, B1 => 
                           REGISTERS_10_21_port, B2 => n865, ZN => n522);
   U1126 : NAND4_X1 port map( A1 => n525, A2 => n524, A3 => n523, A4 => n522, 
                           ZN => n526);
   U1127 : AOI22_X1 port map( A1 => n527, A2 => n890, B1 => n526, B2 => n886, 
                           ZN => n528);
   U1128 : OAI221_X1 port map( B1 => n898, B2 => n530, C1 => n895, C2 => n529, 
                           A => n528, ZN => N203);
   U1129 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n778, B1 => 
                           REGISTERS_23_22_port, B2 => n760, ZN => n534);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n814, B1 => 
                           REGISTERS_19_22_port, B2 => n796, ZN => n533);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n850, B1 => 
                           REGISTERS_22_22_port, B2 => n832, ZN => n532);
   U1132 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n877, B1 => 
                           REGISTERS_18_22_port, B2 => n864, ZN => n531);
   U1133 : AND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => n551);
   U1134 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n778, B1 => 
                           REGISTERS_31_22_port, B2 => n760, ZN => n538);
   U1135 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n814, B1 => 
                           REGISTERS_27_22_port, B2 => n796, ZN => n537);
   U1136 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n850, B1 => 
                           REGISTERS_30_22_port, B2 => n832, ZN => n536);
   U1137 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n877, B1 => 
                           REGISTERS_26_22_port, B2 => n864, ZN => n535);
   U1138 : AND4_X1 port map( A1 => n538, A2 => n537, A3 => n536, A4 => n535, ZN
                           => n550);
   U1139 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n778, B1 => 
                           REGISTERS_7_22_port, B2 => n760, ZN => n542);
   U1140 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n814, B1 => 
                           REGISTERS_3_22_port, B2 => n796, ZN => n541);
   U1141 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n850, B1 => 
                           REGISTERS_6_22_port, B2 => n832, ZN => n540);
   U1142 : NAND4_X1 port map( A1 => n542, A2 => n541, A3 => n540, A4 => n539, 
                           ZN => n548);
   U1143 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n778, B1 => 
                           REGISTERS_15_22_port, B2 => n760, ZN => n546);
   U1144 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n814, B1 => 
                           REGISTERS_11_22_port, B2 => n796, ZN => n545);
   U1145 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n850, B1 => 
                           REGISTERS_14_22_port, B2 => n832, ZN => n544);
   U1146 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n877, B1 => 
                           REGISTERS_10_22_port, B2 => n864, ZN => n543);
   U1147 : NAND4_X1 port map( A1 => n546, A2 => n545, A3 => n544, A4 => n543, 
                           ZN => n547);
   U1148 : AOI22_X1 port map( A1 => n548, A2 => n889, B1 => n547, B2 => n885, 
                           ZN => n549);
   U1149 : OAI221_X1 port map( B1 => n897, B2 => n551, C1 => n895, C2 => n550, 
                           A => n549, ZN => N202);
   U1150 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n778, B1 => 
                           REGISTERS_23_23_port, B2 => n760, ZN => n555);
   U1151 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n814, B1 => 
                           REGISTERS_19_23_port, B2 => n796, ZN => n554);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n850, B1 => 
                           REGISTERS_22_23_port, B2 => n832, ZN => n553);
   U1153 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n877, B1 => 
                           REGISTERS_18_23_port, B2 => n864, ZN => n552);
   U1154 : AND4_X1 port map( A1 => n555, A2 => n554, A3 => n553, A4 => n552, ZN
                           => n572);
   U1155 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n778, B1 => 
                           REGISTERS_31_23_port, B2 => n760, ZN => n559);
   U1156 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n814, B1 => 
                           REGISTERS_27_23_port, B2 => n796, ZN => n558);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n850, B1 => 
                           REGISTERS_30_23_port, B2 => n832, ZN => n557);
   U1158 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n877, B1 => 
                           REGISTERS_26_23_port, B2 => n864, ZN => n556);
   U1159 : AND4_X1 port map( A1 => n559, A2 => n558, A3 => n557, A4 => n556, ZN
                           => n571);
   U1160 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n778, B1 => 
                           REGISTERS_7_23_port, B2 => n760, ZN => n563);
   U1161 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n814, B1 => 
                           REGISTERS_3_23_port, B2 => n796, ZN => n562);
   U1162 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n850, B1 => 
                           REGISTERS_6_23_port, B2 => n832, ZN => n561);
   U1163 : NAND4_X1 port map( A1 => n563, A2 => n562, A3 => n561, A4 => n560, 
                           ZN => n569);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n778, B1 => 
                           REGISTERS_15_23_port, B2 => n760, ZN => n567);
   U1165 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n814, B1 => 
                           REGISTERS_11_23_port, B2 => n796, ZN => n566);
   U1166 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n850, B1 => 
                           REGISTERS_14_23_port, B2 => n832, ZN => n565);
   U1167 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n877, B1 => 
                           REGISTERS_10_23_port, B2 => n864, ZN => n564);
   U1168 : NAND4_X1 port map( A1 => n567, A2 => n566, A3 => n565, A4 => n564, 
                           ZN => n568);
   U1169 : AOI22_X1 port map( A1 => n569, A2 => n889, B1 => n568, B2 => n885, 
                           ZN => n570);
   U1170 : OAI221_X1 port map( B1 => n897, B2 => n572, C1 => n895, C2 => n571, 
                           A => n570, ZN => N201);
   U1171 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n778, B1 => 
                           REGISTERS_23_24_port, B2 => n760, ZN => n576);
   U1172 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n814, B1 => 
                           REGISTERS_19_24_port, B2 => n796, ZN => n575);
   U1173 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n850, B1 => 
                           REGISTERS_22_24_port, B2 => n832, ZN => n574);
   U1174 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n877, B1 => 
                           REGISTERS_18_24_port, B2 => n864, ZN => n573);
   U1175 : AND4_X1 port map( A1 => n576, A2 => n575, A3 => n574, A4 => n573, ZN
                           => n593);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n778, B1 => 
                           REGISTERS_31_24_port, B2 => n760, ZN => n580);
   U1177 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n814, B1 => 
                           REGISTERS_27_24_port, B2 => n796, ZN => n579);
   U1178 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n850, B1 => 
                           REGISTERS_30_24_port, B2 => n832, ZN => n578);
   U1179 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n877, B1 => 
                           REGISTERS_26_24_port, B2 => n864, ZN => n577);
   U1180 : AND4_X1 port map( A1 => n580, A2 => n579, A3 => n578, A4 => n577, ZN
                           => n592);
   U1181 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n778, B1 => 
                           REGISTERS_7_24_port, B2 => n760, ZN => n584);
   U1182 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n814, B1 => 
                           REGISTERS_3_24_port, B2 => n796, ZN => n583);
   U1183 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n850, B1 => 
                           REGISTERS_6_24_port, B2 => n832, ZN => n582);
   U1184 : NAND4_X1 port map( A1 => n584, A2 => n583, A3 => n582, A4 => n581, 
                           ZN => n590);
   U1185 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n777, B1 => 
                           REGISTERS_15_24_port, B2 => n759, ZN => n588);
   U1186 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n813, B1 => 
                           REGISTERS_11_24_port, B2 => n795, ZN => n587);
   U1187 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n849, B1 => 
                           REGISTERS_14_24_port, B2 => n831, ZN => n586);
   U1188 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n877, B1 => 
                           REGISTERS_10_24_port, B2 => n864, ZN => n585);
   U1189 : NAND4_X1 port map( A1 => n588, A2 => n587, A3 => n586, A4 => n585, 
                           ZN => n589);
   U1190 : AOI22_X1 port map( A1 => n590, A2 => n889, B1 => n589, B2 => n885, 
                           ZN => n591);
   U1191 : OAI221_X1 port map( B1 => n897, B2 => n593, C1 => n895, C2 => n592, 
                           A => n591, ZN => N200);
   U1192 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n777, B1 => 
                           REGISTERS_23_25_port, B2 => n759, ZN => n597);
   U1193 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n813, B1 => 
                           REGISTERS_19_25_port, B2 => n795, ZN => n596);
   U1194 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n849, B1 => 
                           REGISTERS_22_25_port, B2 => n831, ZN => n595);
   U1195 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n877, B1 => 
                           REGISTERS_18_25_port, B2 => n864, ZN => n594);
   U1196 : AND4_X1 port map( A1 => n597, A2 => n596, A3 => n595, A4 => n594, ZN
                           => n614);
   U1197 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n777, B1 => 
                           REGISTERS_31_25_port, B2 => n759, ZN => n601);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n813, B1 => 
                           REGISTERS_27_25_port, B2 => n795, ZN => n600);
   U1199 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n849, B1 => 
                           REGISTERS_30_25_port, B2 => n831, ZN => n599);
   U1200 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n877, B1 => 
                           REGISTERS_26_25_port, B2 => n864, ZN => n598);
   U1201 : AND4_X1 port map( A1 => n601, A2 => n600, A3 => n599, A4 => n598, ZN
                           => n613);
   U1202 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n777, B1 => 
                           REGISTERS_7_25_port, B2 => n759, ZN => n605);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n813, B1 => 
                           REGISTERS_3_25_port, B2 => n795, ZN => n604);
   U1204 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n849, B1 => 
                           REGISTERS_6_25_port, B2 => n831, ZN => n603);
   U1205 : NAND4_X1 port map( A1 => n605, A2 => n604, A3 => n603, A4 => n602, 
                           ZN => n611);
   U1206 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n777, B1 => 
                           REGISTERS_15_25_port, B2 => n759, ZN => n609);
   U1207 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n813, B1 => 
                           REGISTERS_11_25_port, B2 => n795, ZN => n608);
   U1208 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n849, B1 => 
                           REGISTERS_14_25_port, B2 => n831, ZN => n607);
   U1209 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n876, B1 => 
                           REGISTERS_10_25_port, B2 => n864, ZN => n606);
   U1210 : NAND4_X1 port map( A1 => n609, A2 => n608, A3 => n607, A4 => n606, 
                           ZN => n610);
   U1211 : AOI22_X1 port map( A1 => n611, A2 => n889, B1 => n610, B2 => n885, 
                           ZN => n612);
   U1212 : OAI221_X1 port map( B1 => n897, B2 => n614, C1 => n895, C2 => n613, 
                           A => n612, ZN => N199);
   U1213 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n777, B1 => 
                           REGISTERS_23_26_port, B2 => n759, ZN => n618);
   U1214 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n813, B1 => 
                           REGISTERS_19_26_port, B2 => n795, ZN => n617);
   U1215 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n849, B1 => 
                           REGISTERS_22_26_port, B2 => n831, ZN => n616);
   U1216 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n876, B1 => 
                           REGISTERS_18_26_port, B2 => n864, ZN => n615);
   U1217 : AND4_X1 port map( A1 => n618, A2 => n617, A3 => n616, A4 => n615, ZN
                           => n635);
   U1218 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n777, B1 => 
                           REGISTERS_31_26_port, B2 => n759, ZN => n622);
   U1219 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n813, B1 => 
                           REGISTERS_27_26_port, B2 => n795, ZN => n621);
   U1220 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n849, B1 => 
                           REGISTERS_30_26_port, B2 => n831, ZN => n620);
   U1221 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n876, B1 => 
                           REGISTERS_26_26_port, B2 => n864, ZN => n619);
   U1222 : AND4_X1 port map( A1 => n622, A2 => n621, A3 => n620, A4 => n619, ZN
                           => n634);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n777, B1 => 
                           REGISTERS_7_26_port, B2 => n759, ZN => n626);
   U1224 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n813, B1 => 
                           REGISTERS_3_26_port, B2 => n795, ZN => n625);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n849, B1 => 
                           REGISTERS_6_26_port, B2 => n831, ZN => n624);
   U1226 : NAND4_X1 port map( A1 => n626, A2 => n625, A3 => n624, A4 => n623, 
                           ZN => n632);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n777, B1 => 
                           REGISTERS_15_26_port, B2 => n759, ZN => n630);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n813, B1 => 
                           REGISTERS_11_26_port, B2 => n795, ZN => n629);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n849, B1 => 
                           REGISTERS_14_26_port, B2 => n831, ZN => n628);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n876, B1 => 
                           REGISTERS_10_26_port, B2 => n864, ZN => n627);
   U1231 : NAND4_X1 port map( A1 => n630, A2 => n629, A3 => n628, A4 => n627, 
                           ZN => n631);
   U1232 : AOI22_X1 port map( A1 => n632, A2 => n889, B1 => n631, B2 => n885, 
                           ZN => n633);
   U1233 : OAI221_X1 port map( B1 => n897, B2 => n635, C1 => n895, C2 => n634, 
                           A => n633, ZN => N198);
   U1234 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n777, B1 => 
                           REGISTERS_23_27_port, B2 => n759, ZN => n639);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n813, B1 => 
                           REGISTERS_19_27_port, B2 => n795, ZN => n638);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n849, B1 => 
                           REGISTERS_22_27_port, B2 => n831, ZN => n637);
   U1237 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n876, B1 => 
                           REGISTERS_18_27_port, B2 => n864, ZN => n636);
   U1238 : AND4_X1 port map( A1 => n639, A2 => n638, A3 => n637, A4 => n636, ZN
                           => n656);
   U1239 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n777, B1 => 
                           REGISTERS_31_27_port, B2 => n759, ZN => n643);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n813, B1 => 
                           REGISTERS_27_27_port, B2 => n795, ZN => n642);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n849, B1 => 
                           REGISTERS_30_27_port, B2 => n831, ZN => n641);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n876, B1 => 
                           REGISTERS_26_27_port, B2 => n864, ZN => n640);
   U1243 : AND4_X1 port map( A1 => n643, A2 => n642, A3 => n641, A4 => n640, ZN
                           => n655);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n776, B1 => 
                           REGISTERS_7_27_port, B2 => n758, ZN => n647);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n812, B1 => 
                           REGISTERS_3_27_port, B2 => n794, ZN => n646);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n848, B1 => 
                           REGISTERS_6_27_port, B2 => n830, ZN => n645);
   U1247 : NAND4_X1 port map( A1 => n647, A2 => n646, A3 => n645, A4 => n644, 
                           ZN => n653);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n776, B1 => 
                           REGISTERS_15_27_port, B2 => n758, ZN => n651);
   U1249 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n812, B1 => 
                           REGISTERS_11_27_port, B2 => n794, ZN => n650);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n848, B1 => 
                           REGISTERS_14_27_port, B2 => n830, ZN => n649);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n876, B1 => 
                           REGISTERS_10_27_port, B2 => n864, ZN => n648);
   U1252 : NAND4_X1 port map( A1 => n651, A2 => n650, A3 => n649, A4 => n648, 
                           ZN => n652);
   U1253 : AOI22_X1 port map( A1 => n653, A2 => n889, B1 => n652, B2 => n885, 
                           ZN => n654);
   U1254 : OAI221_X1 port map( B1 => n897, B2 => n656, C1 => n895, C2 => n655, 
                           A => n654, ZN => N197);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n776, B1 => 
                           REGISTERS_23_28_port, B2 => n758, ZN => n660);
   U1256 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n812, B1 => 
                           REGISTERS_19_28_port, B2 => n794, ZN => n659);
   U1257 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n848, B1 => 
                           REGISTERS_22_28_port, B2 => n830, ZN => n658);
   U1258 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n876, B1 => 
                           REGISTERS_18_28_port, B2 => n864, ZN => n657);
   U1259 : AND4_X1 port map( A1 => n660, A2 => n659, A3 => n658, A4 => n657, ZN
                           => n677);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n776, B1 => 
                           REGISTERS_31_28_port, B2 => n758, ZN => n664);
   U1261 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n812, B1 => 
                           REGISTERS_27_28_port, B2 => n794, ZN => n663);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n848, B1 => 
                           REGISTERS_30_28_port, B2 => n830, ZN => n662);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n876, B1 => 
                           REGISTERS_26_28_port, B2 => n864, ZN => n661);
   U1264 : AND4_X1 port map( A1 => n664, A2 => n663, A3 => n662, A4 => n661, ZN
                           => n676);
   U1265 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n776, B1 => 
                           REGISTERS_7_28_port, B2 => n758, ZN => n668);
   U1266 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n812, B1 => 
                           REGISTERS_3_28_port, B2 => n794, ZN => n667);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n848, B1 => 
                           REGISTERS_6_28_port, B2 => n830, ZN => n666);
   U1268 : NAND4_X1 port map( A1 => n668, A2 => n667, A3 => n666, A4 => n665, 
                           ZN => n674);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n776, B1 => 
                           REGISTERS_15_28_port, B2 => n758, ZN => n672);
   U1270 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n812, B1 => 
                           REGISTERS_11_28_port, B2 => n794, ZN => n671);
   U1271 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n848, B1 => 
                           REGISTERS_14_28_port, B2 => n830, ZN => n670);
   U1272 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n876, B1 => 
                           REGISTERS_10_28_port, B2 => n863, ZN => n669);
   U1273 : NAND4_X1 port map( A1 => n672, A2 => n671, A3 => n670, A4 => n669, 
                           ZN => n673);
   U1274 : AOI22_X1 port map( A1 => n674, A2 => n889, B1 => n673, B2 => n885, 
                           ZN => n675);
   U1275 : OAI221_X1 port map( B1 => n897, B2 => n677, C1 => n895, C2 => n676, 
                           A => n675, ZN => N196);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n776, B1 => 
                           REGISTERS_23_29_port, B2 => n758, ZN => n681);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n812, B1 => 
                           REGISTERS_19_29_port, B2 => n794, ZN => n680);
   U1278 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n848, B1 => 
                           REGISTERS_22_29_port, B2 => n830, ZN => n679);
   U1279 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n876, B1 => 
                           REGISTERS_18_29_port, B2 => n863, ZN => n678);
   U1280 : AND4_X1 port map( A1 => n681, A2 => n680, A3 => n679, A4 => n678, ZN
                           => n698);
   U1281 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n776, B1 => 
                           REGISTERS_31_29_port, B2 => n758, ZN => n685);
   U1282 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n812, B1 => 
                           REGISTERS_27_29_port, B2 => n794, ZN => n684);
   U1283 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n848, B1 => 
                           REGISTERS_30_29_port, B2 => n830, ZN => n683);
   U1284 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n875, B1 => 
                           REGISTERS_26_29_port, B2 => n863, ZN => n682);
   U1285 : AND4_X1 port map( A1 => n685, A2 => n684, A3 => n683, A4 => n682, ZN
                           => n697);
   U1286 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n776, B1 => 
                           REGISTERS_7_29_port, B2 => n758, ZN => n689);
   U1287 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n812, B1 => 
                           REGISTERS_3_29_port, B2 => n794, ZN => n688);
   U1288 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n848, B1 => 
                           REGISTERS_6_29_port, B2 => n830, ZN => n687);
   U1289 : NAND4_X1 port map( A1 => n689, A2 => n688, A3 => n687, A4 => n686, 
                           ZN => n695);
   U1290 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n776, B1 => 
                           REGISTERS_15_29_port, B2 => n758, ZN => n693);
   U1291 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n812, B1 => 
                           REGISTERS_11_29_port, B2 => n794, ZN => n692);
   U1292 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n848, B1 => 
                           REGISTERS_14_29_port, B2 => n830, ZN => n691);
   U1293 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n875, B1 => 
                           REGISTERS_10_29_port, B2 => n863, ZN => n690);
   U1294 : NAND4_X1 port map( A1 => n693, A2 => n692, A3 => n691, A4 => n690, 
                           ZN => n694);
   U1295 : AOI22_X1 port map( A1 => n695, A2 => n889, B1 => n694, B2 => n885, 
                           ZN => n696);
   U1296 : OAI221_X1 port map( B1 => n897, B2 => n698, C1 => n895, C2 => n697, 
                           A => n696, ZN => N195);
   U1297 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n776, B1 => 
                           REGISTERS_23_30_port, B2 => n758, ZN => n702);
   U1298 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n812, B1 => 
                           REGISTERS_19_30_port, B2 => n794, ZN => n701);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n848, B1 => 
                           REGISTERS_22_30_port, B2 => n830, ZN => n700);
   U1300 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n875, B1 => 
                           REGISTERS_18_30_port, B2 => n863, ZN => n699);
   U1301 : AND4_X1 port map( A1 => n702, A2 => n701, A3 => n700, A4 => n699, ZN
                           => n719);
   U1302 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n775, B1 => 
                           REGISTERS_31_30_port, B2 => n757, ZN => n706);
   U1303 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n811, B1 => 
                           REGISTERS_27_30_port, B2 => n793, ZN => n705);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n847, B1 => 
                           REGISTERS_30_30_port, B2 => n829, ZN => n704);
   U1305 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n875, B1 => 
                           REGISTERS_26_30_port, B2 => n863, ZN => n703);
   U1306 : AND4_X1 port map( A1 => n706, A2 => n705, A3 => n704, A4 => n703, ZN
                           => n718);
   U1307 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n775, B1 => 
                           REGISTERS_7_30_port, B2 => n757, ZN => n710);
   U1308 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n811, B1 => 
                           REGISTERS_3_30_port, B2 => n793, ZN => n709);
   U1309 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n847, B1 => 
                           REGISTERS_6_30_port, B2 => n829, ZN => n708);
   U1310 : NAND4_X1 port map( A1 => n710, A2 => n709, A3 => n708, A4 => n707, 
                           ZN => n716);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n775, B1 => 
                           REGISTERS_15_30_port, B2 => n757, ZN => n714);
   U1312 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n811, B1 => 
                           REGISTERS_11_30_port, B2 => n793, ZN => n713);
   U1313 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n847, B1 => 
                           REGISTERS_14_30_port, B2 => n829, ZN => n712);
   U1314 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n875, B1 => 
                           REGISTERS_10_30_port, B2 => n863, ZN => n711);
   U1315 : NAND4_X1 port map( A1 => n714, A2 => n713, A3 => n712, A4 => n711, 
                           ZN => n715);
   U1316 : AOI22_X1 port map( A1 => n716, A2 => n889, B1 => n715, B2 => n885, 
                           ZN => n717);
   U1317 : OAI221_X1 port map( B1 => n897, B2 => n719, C1 => n895, C2 => n718, 
                           A => n717, ZN => N194);
   U1318 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n775, B1 => 
                           REGISTERS_23_31_port, B2 => n757, ZN => n723);
   U1319 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n811, B1 => 
                           REGISTERS_19_31_port, B2 => n793, ZN => n722);
   U1320 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n847, B1 => 
                           REGISTERS_22_31_port, B2 => n829, ZN => n721);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n875, B1 => 
                           REGISTERS_18_31_port, B2 => n863, ZN => n720);
   U1322 : AND4_X1 port map( A1 => n723, A2 => n722, A3 => n721, A4 => n720, ZN
                           => n746);
   U1323 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n775, B1 => 
                           REGISTERS_31_31_port, B2 => n757, ZN => n727);
   U1324 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n811, B1 => 
                           REGISTERS_27_31_port, B2 => n793, ZN => n726);
   U1325 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n847, B1 => 
                           REGISTERS_30_31_port, B2 => n829, ZN => n725);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n875, B1 => 
                           REGISTERS_26_31_port, B2 => n863, ZN => n724);
   U1327 : AND4_X1 port map( A1 => n727, A2 => n726, A3 => n725, A4 => n724, ZN
                           => n744);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n775, B1 => 
                           REGISTERS_7_31_port, B2 => n757, ZN => n731);
   U1329 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n811, B1 => 
                           REGISTERS_3_31_port, B2 => n793, ZN => n730);
   U1330 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n847, B1 => 
                           REGISTERS_6_31_port, B2 => n829, ZN => n729);
   U1331 : NAND4_X1 port map( A1 => n731, A2 => n730, A3 => n729, A4 => n728, 
                           ZN => n740);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n775, B1 => 
                           REGISTERS_15_31_port, B2 => n757, ZN => n737);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n811, B1 => 
                           REGISTERS_11_31_port, B2 => n793, ZN => n736);
   U1334 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n847, B1 => 
                           REGISTERS_14_31_port, B2 => n829, ZN => n735);
   U1335 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n875, B1 => 
                           REGISTERS_10_31_port, B2 => n863, ZN => n734);
   U1336 : NAND4_X1 port map( A1 => n737, A2 => n736, A3 => n735, A4 => n734, 
                           ZN => n738);
   U1337 : AOI22_X1 port map( A1 => n889, A2 => n740, B1 => n885, B2 => n738, 
                           ZN => n742);
   U1338 : OAI221_X1 port map( B1 => n746, B2 => n897, C1 => n744, C2 => n895, 
                           A => n742, ZN => N193);
   U1339 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n1585, ZN => n1580);
   U1340 : NOR2_X1 port map( A1 => n1584, A2 => ADD_RD2(1), ZN => n900);
   U1341 : NOR2_X1 port map( A1 => n1584, A2 => n1583, ZN => n901);
   U1342 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n1621, B1 => 
                           REGISTERS_23_0_port, B2 => n1603, ZN => n907);
   U1343 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n902);
   U1344 : NOR2_X1 port map( A1 => n1583, A2 => ADD_RD2(2), ZN => n903);
   U1345 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n1657, B1 => 
                           REGISTERS_19_0_port, B2 => n1639, ZN => n906);
   U1346 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n1693, B1 => 
                           REGISTERS_22_0_port, B2 => n1675, ZN => n905);
   U1347 : AND2_X1 port map( A1 => n902, A2 => n1582, ZN => n1568);
   U1348 : AND2_X1 port map( A1 => n903, A2 => n1582, ZN => n1567);
   U1349 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n1718, B1 => 
                           REGISTERS_18_0_port, B2 => n1703, ZN => n904);
   U1350 : AND4_X1 port map( A1 => n907, A2 => n906, A3 => n905, A4 => n904, ZN
                           => n924);
   U1351 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1578);
   U1352 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n1621, B1 => 
                           REGISTERS_31_0_port, B2 => n1603, ZN => n911);
   U1353 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n1657, B1 => 
                           REGISTERS_27_0_port, B2 => n1639, ZN => n910);
   U1354 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n1693, B1 => 
                           REGISTERS_30_0_port, B2 => n1675, ZN => n909);
   U1355 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n1718, B1 => 
                           REGISTERS_26_0_port, B2 => n1703, ZN => n908);
   U1356 : AND4_X1 port map( A1 => n911, A2 => n910, A3 => n909, A4 => n908, ZN
                           => n923);
   U1357 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n1621, B1 => 
                           REGISTERS_7_0_port, B2 => n1603, ZN => n915);
   U1358 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n1657, B1 => 
                           REGISTERS_3_0_port, B2 => n1639, ZN => n914);
   U1359 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n1693, B1 => 
                           REGISTERS_6_0_port, B2 => n1675, ZN => n913);
   U1360 : NAND4_X1 port map( A1 => n915, A2 => n914, A3 => n913, A4 => n912, 
                           ZN => n921);
   U1361 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1576);
   U1362 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n1621, B1 => 
                           REGISTERS_15_0_port, B2 => n1603, ZN => n919);
   U1363 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n1657, B1 => 
                           REGISTERS_11_0_port, B2 => n1639, ZN => n918);
   U1364 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n1693, B1 => 
                           REGISTERS_14_0_port, B2 => n1675, ZN => n917);
   U1365 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n1718, B1 => 
                           REGISTERS_10_0_port, B2 => n1703, ZN => n916);
   U1366 : NAND4_X1 port map( A1 => n919, A2 => n918, A3 => n917, A4 => n916, 
                           ZN => n920);
   U1367 : NOR2_X1 port map( A1 => n1585, A2 => ADD_RD2(4), ZN => n1574);
   U1368 : AOI22_X1 port map( A1 => n921, A2 => n1726, B1 => n920, B2 => n1722,
                           ZN => n922);
   U1369 : OAI221_X1 port map( B1 => n1734, B2 => n924, C1 => n1728, C2 => n923
                           , A => n922, ZN => N290);
   U1370 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n1621, B1 => 
                           REGISTERS_23_1_port, B2 => n1603, ZN => n928);
   U1371 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n1657, B1 => 
                           REGISTERS_19_1_port, B2 => n1639, ZN => n927);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n1693, B1 => 
                           REGISTERS_22_1_port, B2 => n1675, ZN => n926);
   U1373 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n1718, B1 => 
                           REGISTERS_18_1_port, B2 => n1703, ZN => n925);
   U1374 : AND4_X1 port map( A1 => n928, A2 => n927, A3 => n926, A4 => n925, ZN
                           => n945);
   U1375 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n1621, B1 => 
                           REGISTERS_31_1_port, B2 => n1603, ZN => n932);
   U1376 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n1657, B1 => 
                           REGISTERS_27_1_port, B2 => n1639, ZN => n931);
   U1377 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n1693, B1 => 
                           REGISTERS_30_1_port, B2 => n1675, ZN => n930);
   U1378 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n1718, B1 => 
                           REGISTERS_26_1_port, B2 => n1703, ZN => n929);
   U1379 : AND4_X1 port map( A1 => n932, A2 => n931, A3 => n930, A4 => n929, ZN
                           => n944);
   U1380 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n1621, B1 => 
                           REGISTERS_7_1_port, B2 => n1603, ZN => n936);
   U1381 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n1657, B1 => 
                           REGISTERS_3_1_port, B2 => n1639, ZN => n935);
   U1382 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n1693, B1 => 
                           REGISTERS_6_1_port, B2 => n1675, ZN => n934);
   U1383 : NAND4_X1 port map( A1 => n936, A2 => n935, A3 => n934, A4 => n933, 
                           ZN => n942);
   U1384 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n1621, B1 => 
                           REGISTERS_15_1_port, B2 => n1603, ZN => n940);
   U1385 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n1657, B1 => 
                           REGISTERS_11_1_port, B2 => n1639, ZN => n939);
   U1386 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n1693, B1 => 
                           REGISTERS_14_1_port, B2 => n1675, ZN => n938);
   U1387 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n1718, B1 => 
                           REGISTERS_10_1_port, B2 => n1703, ZN => n937);
   U1388 : NAND4_X1 port map( A1 => n940, A2 => n939, A3 => n938, A4 => n937, 
                           ZN => n941);
   U1389 : AOI22_X1 port map( A1 => n942, A2 => n1726, B1 => n941, B2 => n1722,
                           ZN => n943);
   U1390 : OAI221_X1 port map( B1 => n1734, B2 => n945, C1 => n1728, C2 => n944
                           , A => n943, ZN => N289);
   U1391 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n1621, B1 => 
                           REGISTERS_23_2_port, B2 => n1603, ZN => n949);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n1657, B1 => 
                           REGISTERS_19_2_port, B2 => n1639, ZN => n948);
   U1393 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n1693, B1 => 
                           REGISTERS_22_2_port, B2 => n1675, ZN => n947);
   U1394 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n1718, B1 => 
                           REGISTERS_18_2_port, B2 => n1702, ZN => n946);
   U1395 : AND4_X1 port map( A1 => n949, A2 => n948, A3 => n947, A4 => n946, ZN
                           => n966);
   U1396 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n1621, B1 => 
                           REGISTERS_31_2_port, B2 => n1603, ZN => n953);
   U1397 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n1657, B1 => 
                           REGISTERS_27_2_port, B2 => n1639, ZN => n952);
   U1398 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n1693, B1 => 
                           REGISTERS_30_2_port, B2 => n1675, ZN => n951);
   U1399 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n1718, B1 => 
                           REGISTERS_26_2_port, B2 => n1702, ZN => n950);
   U1400 : AND4_X1 port map( A1 => n953, A2 => n952, A3 => n951, A4 => n950, ZN
                           => n965);
   U1401 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n1621, B1 => 
                           REGISTERS_7_2_port, B2 => n1603, ZN => n957);
   U1402 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n1657, B1 => 
                           REGISTERS_3_2_port, B2 => n1639, ZN => n956);
   U1403 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n1693, B1 => 
                           REGISTERS_6_2_port, B2 => n1675, ZN => n955);
   U1404 : NAND4_X1 port map( A1 => n957, A2 => n956, A3 => n955, A4 => n954, 
                           ZN => n963);
   U1405 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n1620, B1 => 
                           REGISTERS_15_2_port, B2 => n1602, ZN => n961);
   U1406 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n1656, B1 => 
                           REGISTERS_11_2_port, B2 => n1638, ZN => n960);
   U1407 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n1692, B1 => 
                           REGISTERS_14_2_port, B2 => n1674, ZN => n959);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n1718, B1 => 
                           REGISTERS_10_2_port, B2 => n1702, ZN => n958);
   U1409 : NAND4_X1 port map( A1 => n961, A2 => n960, A3 => n959, A4 => n958, 
                           ZN => n962);
   U1410 : AOI22_X1 port map( A1 => n963, A2 => n1726, B1 => n962, B2 => n1722,
                           ZN => n964);
   U1411 : OAI221_X1 port map( B1 => n1734, B2 => n966, C1 => n1728, C2 => n965
                           , A => n964, ZN => N288);
   U1412 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n1620, B1 => 
                           REGISTERS_23_3_port, B2 => n1602, ZN => n970);
   U1413 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n1656, B1 => 
                           REGISTERS_19_3_port, B2 => n1638, ZN => n969);
   U1414 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n1692, B1 => 
                           REGISTERS_22_3_port, B2 => n1674, ZN => n968);
   U1415 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n1718, B1 => 
                           REGISTERS_18_3_port, B2 => n1702, ZN => n967);
   U1416 : AND4_X1 port map( A1 => n970, A2 => n969, A3 => n968, A4 => n967, ZN
                           => n987);
   U1417 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n1620, B1 => 
                           REGISTERS_31_3_port, B2 => n1602, ZN => n974);
   U1418 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n1656, B1 => 
                           REGISTERS_27_3_port, B2 => n1638, ZN => n973);
   U1419 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n1692, B1 => 
                           REGISTERS_30_3_port, B2 => n1674, ZN => n972);
   U1420 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n1718, B1 => 
                           REGISTERS_26_3_port, B2 => n1702, ZN => n971);
   U1421 : AND4_X1 port map( A1 => n974, A2 => n973, A3 => n972, A4 => n971, ZN
                           => n986);
   U1422 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n1620, B1 => 
                           REGISTERS_7_3_port, B2 => n1602, ZN => n978);
   U1423 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n1656, B1 => 
                           REGISTERS_3_3_port, B2 => n1638, ZN => n977);
   U1424 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n1692, B1 => 
                           REGISTERS_6_3_port, B2 => n1674, ZN => n976);
   U1425 : NAND4_X1 port map( A1 => n978, A2 => n977, A3 => n976, A4 => n975, 
                           ZN => n984);
   U1426 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n1620, B1 => 
                           REGISTERS_15_3_port, B2 => n1602, ZN => n982);
   U1427 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n1656, B1 => 
                           REGISTERS_11_3_port, B2 => n1638, ZN => n981);
   U1428 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n1692, B1 => 
                           REGISTERS_14_3_port, B2 => n1674, ZN => n980);
   U1429 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n1717, B1 => 
                           REGISTERS_10_3_port, B2 => n1702, ZN => n979);
   U1430 : NAND4_X1 port map( A1 => n982, A2 => n981, A3 => n980, A4 => n979, 
                           ZN => n983);
   U1431 : AOI22_X1 port map( A1 => n984, A2 => n1726, B1 => n983, B2 => n1722,
                           ZN => n985);
   U1432 : OAI221_X1 port map( B1 => n1734, B2 => n987, C1 => n1728, C2 => n986
                           , A => n985, ZN => N287);
   U1433 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n1620, B1 => 
                           REGISTERS_23_4_port, B2 => n1602, ZN => n991);
   U1434 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n1656, B1 => 
                           REGISTERS_19_4_port, B2 => n1638, ZN => n990);
   U1435 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n1692, B1 => 
                           REGISTERS_22_4_port, B2 => n1674, ZN => n989);
   U1436 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n1717, B1 => 
                           REGISTERS_18_4_port, B2 => n1702, ZN => n988);
   U1437 : AND4_X1 port map( A1 => n991, A2 => n990, A3 => n989, A4 => n988, ZN
                           => n1008);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n1620, B1 => 
                           REGISTERS_31_4_port, B2 => n1602, ZN => n995);
   U1439 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n1656, B1 => 
                           REGISTERS_27_4_port, B2 => n1638, ZN => n994);
   U1440 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n1692, B1 => 
                           REGISTERS_30_4_port, B2 => n1674, ZN => n993);
   U1441 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n1717, B1 => 
                           REGISTERS_26_4_port, B2 => n1702, ZN => n992);
   U1442 : AND4_X1 port map( A1 => n995, A2 => n994, A3 => n993, A4 => n992, ZN
                           => n1007);
   U1443 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n1620, B1 => 
                           REGISTERS_7_4_port, B2 => n1602, ZN => n999);
   U1444 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n1656, B1 => 
                           REGISTERS_3_4_port, B2 => n1638, ZN => n998);
   U1445 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n1692, B1 => 
                           REGISTERS_6_4_port, B2 => n1674, ZN => n997);
   U1446 : NAND4_X1 port map( A1 => n999, A2 => n998, A3 => n997, A4 => n996, 
                           ZN => n1005);
   U1447 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n1620, B1 => 
                           REGISTERS_15_4_port, B2 => n1602, ZN => n1003);
   U1448 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n1656, B1 => 
                           REGISTERS_11_4_port, B2 => n1638, ZN => n1002);
   U1449 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n1692, B1 => 
                           REGISTERS_14_4_port, B2 => n1674, ZN => n1001);
   U1450 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n1717, B1 => 
                           REGISTERS_10_4_port, B2 => n1702, ZN => n1000);
   U1451 : NAND4_X1 port map( A1 => n1003, A2 => n1002, A3 => n1001, A4 => 
                           n1000, ZN => n1004);
   U1452 : AOI22_X1 port map( A1 => n1005, A2 => n1726, B1 => n1004, B2 => 
                           n1722, ZN => n1006);
   U1453 : OAI221_X1 port map( B1 => n1734, B2 => n1008, C1 => n1728, C2 => 
                           n1007, A => n1006, ZN => N286);
   U1454 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n1620, B1 => 
                           REGISTERS_23_5_port, B2 => n1602, ZN => n1012);
   U1455 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n1656, B1 => 
                           REGISTERS_19_5_port, B2 => n1638, ZN => n1011);
   U1456 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n1692, B1 => 
                           REGISTERS_22_5_port, B2 => n1674, ZN => n1010);
   U1457 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n1717, B1 => 
                           REGISTERS_18_5_port, B2 => n1702, ZN => n1009);
   U1458 : AND4_X1 port map( A1 => n1012, A2 => n1011, A3 => n1010, A4 => n1009
                           , ZN => n1029);
   U1459 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n1620, B1 => 
                           REGISTERS_31_5_port, B2 => n1602, ZN => n1016);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n1656, B1 => 
                           REGISTERS_27_5_port, B2 => n1638, ZN => n1015);
   U1461 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n1692, B1 => 
                           REGISTERS_30_5_port, B2 => n1674, ZN => n1014);
   U1462 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n1717, B1 => 
                           REGISTERS_26_5_port, B2 => n1702, ZN => n1013);
   U1463 : AND4_X1 port map( A1 => n1016, A2 => n1015, A3 => n1014, A4 => n1013
                           , ZN => n1028);
   U1464 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n1619, B1 => 
                           REGISTERS_7_5_port, B2 => n1601, ZN => n1020);
   U1465 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n1655, B1 => 
                           REGISTERS_3_5_port, B2 => n1637, ZN => n1019);
   U1466 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n1691, B1 => 
                           REGISTERS_6_5_port, B2 => n1673, ZN => n1018);
   U1467 : NAND4_X1 port map( A1 => n1020, A2 => n1019, A3 => n1018, A4 => 
                           n1017, ZN => n1026);
   U1468 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n1619, B1 => 
                           REGISTERS_15_5_port, B2 => n1601, ZN => n1024);
   U1469 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n1655, B1 => 
                           REGISTERS_11_5_port, B2 => n1637, ZN => n1023);
   U1470 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n1691, B1 => 
                           REGISTERS_14_5_port, B2 => n1673, ZN => n1022);
   U1471 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n1717, B1 => 
                           REGISTERS_10_5_port, B2 => n1702, ZN => n1021);
   U1472 : NAND4_X1 port map( A1 => n1024, A2 => n1023, A3 => n1022, A4 => 
                           n1021, ZN => n1025);
   U1473 : AOI22_X1 port map( A1 => n1026, A2 => n1726, B1 => n1025, B2 => 
                           n1722, ZN => n1027);
   U1474 : OAI221_X1 port map( B1 => n1734, B2 => n1029, C1 => n1728, C2 => 
                           n1028, A => n1027, ZN => N285);
   U1475 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n1619, B1 => 
                           REGISTERS_23_6_port, B2 => n1601, ZN => n1033);
   U1476 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n1655, B1 => 
                           REGISTERS_19_6_port, B2 => n1637, ZN => n1032);
   U1477 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n1691, B1 => 
                           REGISTERS_22_6_port, B2 => n1673, ZN => n1031);
   U1478 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n1717, B1 => 
                           REGISTERS_18_6_port, B2 => n1702, ZN => n1030);
   U1479 : AND4_X1 port map( A1 => n1033, A2 => n1032, A3 => n1031, A4 => n1030
                           , ZN => n1050);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n1619, B1 => 
                           REGISTERS_31_6_port, B2 => n1601, ZN => n1037);
   U1481 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n1655, B1 => 
                           REGISTERS_27_6_port, B2 => n1637, ZN => n1036);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n1691, B1 => 
                           REGISTERS_30_6_port, B2 => n1673, ZN => n1035);
   U1483 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n1717, B1 => 
                           REGISTERS_26_6_port, B2 => n1702, ZN => n1034);
   U1484 : AND4_X1 port map( A1 => n1037, A2 => n1036, A3 => n1035, A4 => n1034
                           , ZN => n1049);
   U1485 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n1619, B1 => 
                           REGISTERS_7_6_port, B2 => n1601, ZN => n1041);
   U1486 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n1655, B1 => 
                           REGISTERS_3_6_port, B2 => n1637, ZN => n1040);
   U1487 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n1691, B1 => 
                           REGISTERS_6_6_port, B2 => n1673, ZN => n1039);
   U1488 : NAND4_X1 port map( A1 => n1041, A2 => n1040, A3 => n1039, A4 => 
                           n1038, ZN => n1047);
   U1489 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n1619, B1 => 
                           REGISTERS_15_6_port, B2 => n1601, ZN => n1045);
   U1490 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n1655, B1 => 
                           REGISTERS_11_6_port, B2 => n1637, ZN => n1044);
   U1491 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n1691, B1 => 
                           REGISTERS_14_6_port, B2 => n1673, ZN => n1043);
   U1492 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n1717, B1 => 
                           REGISTERS_10_6_port, B2 => n1702, ZN => n1042);
   U1493 : NAND4_X1 port map( A1 => n1045, A2 => n1044, A3 => n1043, A4 => 
                           n1042, ZN => n1046);
   U1494 : AOI22_X1 port map( A1 => n1047, A2 => n1726, B1 => n1046, B2 => 
                           n1722, ZN => n1048);
   U1495 : OAI221_X1 port map( B1 => n1734, B2 => n1050, C1 => n1728, C2 => 
                           n1049, A => n1048, ZN => N284);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n1619, B1 => 
                           REGISTERS_23_7_port, B2 => n1601, ZN => n1054);
   U1497 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n1655, B1 => 
                           REGISTERS_19_7_port, B2 => n1637, ZN => n1053);
   U1498 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n1691, B1 => 
                           REGISTERS_22_7_port, B2 => n1673, ZN => n1052);
   U1499 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n1717, B1 => 
                           REGISTERS_18_7_port, B2 => n1702, ZN => n1051);
   U1500 : AND4_X1 port map( A1 => n1054, A2 => n1053, A3 => n1052, A4 => n1051
                           , ZN => n1071);
   U1501 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n1619, B1 => 
                           REGISTERS_31_7_port, B2 => n1601, ZN => n1058);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n1655, B1 => 
                           REGISTERS_27_7_port, B2 => n1637, ZN => n1057);
   U1503 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n1691, B1 => 
                           REGISTERS_30_7_port, B2 => n1673, ZN => n1056);
   U1504 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n1716, B1 => 
                           REGISTERS_26_7_port, B2 => n1702, ZN => n1055);
   U1505 : AND4_X1 port map( A1 => n1058, A2 => n1057, A3 => n1056, A4 => n1055
                           , ZN => n1070);
   U1506 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n1619, B1 => 
                           REGISTERS_7_7_port, B2 => n1601, ZN => n1062);
   U1507 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n1655, B1 => 
                           REGISTERS_3_7_port, B2 => n1637, ZN => n1061);
   U1508 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n1691, B1 => 
                           REGISTERS_6_7_port, B2 => n1673, ZN => n1060);
   U1509 : NAND4_X1 port map( A1 => n1062, A2 => n1061, A3 => n1060, A4 => 
                           n1059, ZN => n1068);
   U1510 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n1619, B1 => 
                           REGISTERS_15_7_port, B2 => n1601, ZN => n1066);
   U1511 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n1655, B1 => 
                           REGISTERS_11_7_port, B2 => n1637, ZN => n1065);
   U1512 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n1691, B1 => 
                           REGISTERS_14_7_port, B2 => n1673, ZN => n1064);
   U1513 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n1716, B1 => 
                           REGISTERS_10_7_port, B2 => n1702, ZN => n1063);
   U1514 : NAND4_X1 port map( A1 => n1066, A2 => n1065, A3 => n1064, A4 => 
                           n1063, ZN => n1067);
   U1515 : AOI22_X1 port map( A1 => n1068, A2 => n1726, B1 => n1067, B2 => 
                           n1722, ZN => n1069);
   U1516 : OAI221_X1 port map( B1 => n1734, B2 => n1071, C1 => n1728, C2 => 
                           n1070, A => n1069, ZN => N283);
   U1517 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n1619, B1 => 
                           REGISTERS_23_8_port, B2 => n1601, ZN => n1075);
   U1518 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n1655, B1 => 
                           REGISTERS_19_8_port, B2 => n1637, ZN => n1074);
   U1519 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n1691, B1 => 
                           REGISTERS_22_8_port, B2 => n1673, ZN => n1073);
   U1520 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n1716, B1 => 
                           REGISTERS_18_8_port, B2 => n1702, ZN => n1072);
   U1521 : AND4_X1 port map( A1 => n1075, A2 => n1074, A3 => n1073, A4 => n1072
                           , ZN => n1092);
   U1522 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n1618, B1 => 
                           REGISTERS_31_8_port, B2 => n1600, ZN => n1079);
   U1523 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n1654, B1 => 
                           REGISTERS_27_8_port, B2 => n1636, ZN => n1078);
   U1524 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n1690, B1 => 
                           REGISTERS_30_8_port, B2 => n1672, ZN => n1077);
   U1525 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n1716, B1 => 
                           REGISTERS_26_8_port, B2 => n1702, ZN => n1076);
   U1526 : AND4_X1 port map( A1 => n1079, A2 => n1078, A3 => n1077, A4 => n1076
                           , ZN => n1091);
   U1527 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n1618, B1 => 
                           REGISTERS_7_8_port, B2 => n1600, ZN => n1083);
   U1528 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n1654, B1 => 
                           REGISTERS_3_8_port, B2 => n1636, ZN => n1082);
   U1529 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n1690, B1 => 
                           REGISTERS_6_8_port, B2 => n1672, ZN => n1081);
   U1530 : NAND4_X1 port map( A1 => n1083, A2 => n1082, A3 => n1081, A4 => 
                           n1080, ZN => n1089);
   U1531 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n1618, B1 => 
                           REGISTERS_15_8_port, B2 => n1600, ZN => n1087);
   U1532 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n1654, B1 => 
                           REGISTERS_11_8_port, B2 => n1636, ZN => n1086);
   U1533 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n1690, B1 => 
                           REGISTERS_14_8_port, B2 => n1672, ZN => n1085);
   U1534 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n1716, B1 => 
                           REGISTERS_10_8_port, B2 => n1701, ZN => n1084);
   U1535 : NAND4_X1 port map( A1 => n1087, A2 => n1086, A3 => n1085, A4 => 
                           n1084, ZN => n1088);
   U1536 : AOI22_X1 port map( A1 => n1089, A2 => n1726, B1 => n1088, B2 => 
                           n1722, ZN => n1090);
   U1537 : OAI221_X1 port map( B1 => n1734, B2 => n1092, C1 => n1728, C2 => 
                           n1091, A => n1090, ZN => N282);
   U1538 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n1618, B1 => 
                           REGISTERS_23_9_port, B2 => n1600, ZN => n1096);
   U1539 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n1654, B1 => 
                           REGISTERS_19_9_port, B2 => n1636, ZN => n1095);
   U1540 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n1690, B1 => 
                           REGISTERS_22_9_port, B2 => n1672, ZN => n1094);
   U1541 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n1716, B1 => 
                           REGISTERS_18_9_port, B2 => n1701, ZN => n1093);
   U1542 : AND4_X1 port map( A1 => n1096, A2 => n1095, A3 => n1094, A4 => n1093
                           , ZN => n1113);
   U1543 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n1618, B1 => 
                           REGISTERS_31_9_port, B2 => n1600, ZN => n1100);
   U1544 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n1654, B1 => 
                           REGISTERS_27_9_port, B2 => n1636, ZN => n1099);
   U1545 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n1690, B1 => 
                           REGISTERS_30_9_port, B2 => n1672, ZN => n1098);
   U1546 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n1716, B1 => 
                           REGISTERS_26_9_port, B2 => n1701, ZN => n1097);
   U1547 : AND4_X1 port map( A1 => n1100, A2 => n1099, A3 => n1098, A4 => n1097
                           , ZN => n1112);
   U1548 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n1618, B1 => 
                           REGISTERS_7_9_port, B2 => n1600, ZN => n1104);
   U1549 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n1654, B1 => 
                           REGISTERS_3_9_port, B2 => n1636, ZN => n1103);
   U1550 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n1690, B1 => 
                           REGISTERS_6_9_port, B2 => n1672, ZN => n1102);
   U1551 : NAND4_X1 port map( A1 => n1104, A2 => n1103, A3 => n1102, A4 => 
                           n1101, ZN => n1110);
   U1552 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n1618, B1 => 
                           REGISTERS_15_9_port, B2 => n1600, ZN => n1108);
   U1553 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n1654, B1 => 
                           REGISTERS_11_9_port, B2 => n1636, ZN => n1107);
   U1554 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n1690, B1 => 
                           REGISTERS_14_9_port, B2 => n1672, ZN => n1106);
   U1555 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n1716, B1 => 
                           REGISTERS_10_9_port, B2 => n1701, ZN => n1105);
   U1556 : NAND4_X1 port map( A1 => n1108, A2 => n1107, A3 => n1106, A4 => 
                           n1105, ZN => n1109);
   U1557 : AOI22_X1 port map( A1 => n1110, A2 => n1726, B1 => n1109, B2 => 
                           n1722, ZN => n1111);
   U1558 : OAI221_X1 port map( B1 => n1734, B2 => n1113, C1 => n1728, C2 => 
                           n1112, A => n1111, ZN => N281);
   U1559 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n1618, B1 => 
                           REGISTERS_23_10_port, B2 => n1600, ZN => n1117);
   U1560 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n1654, B1 => 
                           REGISTERS_19_10_port, B2 => n1636, ZN => n1116);
   U1561 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n1690, B1 => 
                           REGISTERS_22_10_port, B2 => n1672, ZN => n1115);
   U1562 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n1716, B1 => 
                           REGISTERS_18_10_port, B2 => n1701, ZN => n1114);
   U1563 : AND4_X1 port map( A1 => n1117, A2 => n1116, A3 => n1115, A4 => n1114
                           , ZN => n1134);
   U1564 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n1618, B1 => 
                           REGISTERS_31_10_port, B2 => n1600, ZN => n1121);
   U1565 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n1654, B1 => 
                           REGISTERS_27_10_port, B2 => n1636, ZN => n1120);
   U1566 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n1690, B1 => 
                           REGISTERS_30_10_port, B2 => n1672, ZN => n1119);
   U1567 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n1716, B1 => 
                           REGISTERS_26_10_port, B2 => n1701, ZN => n1118);
   U1568 : AND4_X1 port map( A1 => n1121, A2 => n1120, A3 => n1119, A4 => n1118
                           , ZN => n1133);
   U1569 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n1618, B1 => 
                           REGISTERS_7_10_port, B2 => n1600, ZN => n1125);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n1654, B1 => 
                           REGISTERS_3_10_port, B2 => n1636, ZN => n1124);
   U1571 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n1690, B1 => 
                           REGISTERS_6_10_port, B2 => n1672, ZN => n1123);
   U1572 : NAND4_X1 port map( A1 => n1125, A2 => n1124, A3 => n1123, A4 => 
                           n1122, ZN => n1131);
   U1573 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n1618, B1 => 
                           REGISTERS_15_10_port, B2 => n1600, ZN => n1129);
   U1574 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n1654, B1 => 
                           REGISTERS_11_10_port, B2 => n1636, ZN => n1128);
   U1575 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n1690, B1 => 
                           REGISTERS_14_10_port, B2 => n1672, ZN => n1127);
   U1576 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n1716, B1 => 
                           REGISTERS_10_10_port, B2 => n1701, ZN => n1126);
   U1577 : NAND4_X1 port map( A1 => n1129, A2 => n1128, A3 => n1127, A4 => 
                           n1126, ZN => n1130);
   U1578 : AOI22_X1 port map( A1 => n1131, A2 => n1726, B1 => n1130, B2 => 
                           n1722, ZN => n1132);
   U1579 : OAI221_X1 port map( B1 => n1734, B2 => n1134, C1 => n1729, C2 => 
                           n1133, A => n1132, ZN => N280);
   U1580 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n1617, B1 => 
                           REGISTERS_23_11_port, B2 => n1599, ZN => n1138);
   U1581 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n1653, B1 => 
                           REGISTERS_19_11_port, B2 => n1635, ZN => n1137);
   U1582 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n1689, B1 => 
                           REGISTERS_22_11_port, B2 => n1671, ZN => n1136);
   U1583 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n1715, B1 => 
                           REGISTERS_18_11_port, B2 => n1701, ZN => n1135);
   U1584 : AND4_X1 port map( A1 => n1138, A2 => n1137, A3 => n1136, A4 => n1135
                           , ZN => n1155);
   U1585 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n1617, B1 => 
                           REGISTERS_31_11_port, B2 => n1599, ZN => n1142);
   U1586 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n1653, B1 => 
                           REGISTERS_27_11_port, B2 => n1635, ZN => n1141);
   U1587 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n1689, B1 => 
                           REGISTERS_30_11_port, B2 => n1671, ZN => n1140);
   U1588 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n1715, B1 => 
                           REGISTERS_26_11_port, B2 => n1701, ZN => n1139);
   U1589 : AND4_X1 port map( A1 => n1142, A2 => n1141, A3 => n1140, A4 => n1139
                           , ZN => n1154);
   U1590 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n1617, B1 => 
                           REGISTERS_7_11_port, B2 => n1599, ZN => n1146);
   U1591 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n1653, B1 => 
                           REGISTERS_3_11_port, B2 => n1635, ZN => n1145);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n1689, B1 => 
                           REGISTERS_6_11_port, B2 => n1671, ZN => n1144);
   U1593 : NAND4_X1 port map( A1 => n1146, A2 => n1145, A3 => n1144, A4 => 
                           n1143, ZN => n1152);
   U1594 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n1617, B1 => 
                           REGISTERS_15_11_port, B2 => n1599, ZN => n1150);
   U1595 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n1653, B1 => 
                           REGISTERS_11_11_port, B2 => n1635, ZN => n1149);
   U1596 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n1689, B1 => 
                           REGISTERS_14_11_port, B2 => n1671, ZN => n1148);
   U1597 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n1715, B1 => 
                           REGISTERS_10_11_port, B2 => n1701, ZN => n1147);
   U1598 : NAND4_X1 port map( A1 => n1150, A2 => n1149, A3 => n1148, A4 => 
                           n1147, ZN => n1151);
   U1599 : AOI22_X1 port map( A1 => n1152, A2 => n1725, B1 => n1151, B2 => 
                           n1721, ZN => n1153);
   U1600 : OAI221_X1 port map( B1 => n1733, B2 => n1155, C1 => n1729, C2 => 
                           n1154, A => n1153, ZN => N279);
   U1601 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n1617, B1 => 
                           REGISTERS_23_12_port, B2 => n1599, ZN => n1159);
   U1602 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n1653, B1 => 
                           REGISTERS_19_12_port, B2 => n1635, ZN => n1158);
   U1603 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n1689, B1 => 
                           REGISTERS_22_12_port, B2 => n1671, ZN => n1157);
   U1604 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n1715, B1 => 
                           REGISTERS_18_12_port, B2 => n1701, ZN => n1156);
   U1605 : AND4_X1 port map( A1 => n1159, A2 => n1158, A3 => n1157, A4 => n1156
                           , ZN => n1176);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n1617, B1 => 
                           REGISTERS_31_12_port, B2 => n1599, ZN => n1163);
   U1607 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n1653, B1 => 
                           REGISTERS_27_12_port, B2 => n1635, ZN => n1162);
   U1608 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n1689, B1 => 
                           REGISTERS_30_12_port, B2 => n1671, ZN => n1161);
   U1609 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n1715, B1 => 
                           REGISTERS_26_12_port, B2 => n1701, ZN => n1160);
   U1610 : AND4_X1 port map( A1 => n1163, A2 => n1162, A3 => n1161, A4 => n1160
                           , ZN => n1175);
   U1611 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n1617, B1 => 
                           REGISTERS_7_12_port, B2 => n1599, ZN => n1167);
   U1612 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n1653, B1 => 
                           REGISTERS_3_12_port, B2 => n1635, ZN => n1166);
   U1613 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n1689, B1 => 
                           REGISTERS_6_12_port, B2 => n1671, ZN => n1165);
   U1614 : NAND4_X1 port map( A1 => n1167, A2 => n1166, A3 => n1165, A4 => 
                           n1164, ZN => n1173);
   U1615 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n1617, B1 => 
                           REGISTERS_15_12_port, B2 => n1599, ZN => n1171);
   U1616 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n1653, B1 => 
                           REGISTERS_11_12_port, B2 => n1635, ZN => n1170);
   U1617 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n1689, B1 => 
                           REGISTERS_14_12_port, B2 => n1671, ZN => n1169);
   U1618 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n1715, B1 => 
                           REGISTERS_10_12_port, B2 => n1701, ZN => n1168);
   U1619 : NAND4_X1 port map( A1 => n1171, A2 => n1170, A3 => n1169, A4 => 
                           n1168, ZN => n1172);
   U1620 : AOI22_X1 port map( A1 => n1173, A2 => n1725, B1 => n1172, B2 => 
                           n1721, ZN => n1174);
   U1621 : OAI221_X1 port map( B1 => n1733, B2 => n1176, C1 => n1729, C2 => 
                           n1175, A => n1174, ZN => N278);
   U1622 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n1617, B1 => 
                           REGISTERS_23_13_port, B2 => n1599, ZN => n1180);
   U1623 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n1653, B1 => 
                           REGISTERS_19_13_port, B2 => n1635, ZN => n1179);
   U1624 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n1689, B1 => 
                           REGISTERS_22_13_port, B2 => n1671, ZN => n1178);
   U1625 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n1715, B1 => 
                           REGISTERS_18_13_port, B2 => n1701, ZN => n1177);
   U1626 : AND4_X1 port map( A1 => n1180, A2 => n1179, A3 => n1178, A4 => n1177
                           , ZN => n1197);
   U1627 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n1617, B1 => 
                           REGISTERS_31_13_port, B2 => n1599, ZN => n1184);
   U1628 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n1653, B1 => 
                           REGISTERS_27_13_port, B2 => n1635, ZN => n1183);
   U1629 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n1689, B1 => 
                           REGISTERS_30_13_port, B2 => n1671, ZN => n1182);
   U1630 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n1715, B1 => 
                           REGISTERS_26_13_port, B2 => n1701, ZN => n1181);
   U1631 : AND4_X1 port map( A1 => n1184, A2 => n1183, A3 => n1182, A4 => n1181
                           , ZN => n1196);
   U1632 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n1617, B1 => 
                           REGISTERS_7_13_port, B2 => n1599, ZN => n1188);
   U1633 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n1653, B1 => 
                           REGISTERS_3_13_port, B2 => n1635, ZN => n1187);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n1689, B1 => 
                           REGISTERS_6_13_port, B2 => n1671, ZN => n1186);
   U1635 : NAND4_X1 port map( A1 => n1188, A2 => n1187, A3 => n1186, A4 => 
                           n1185, ZN => n1194);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n1616, B1 => 
                           REGISTERS_15_13_port, B2 => n1598, ZN => n1192);
   U1637 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n1652, B1 => 
                           REGISTERS_11_13_port, B2 => n1634, ZN => n1191);
   U1638 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n1688, B1 => 
                           REGISTERS_14_13_port, B2 => n1670, ZN => n1190);
   U1639 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n1715, B1 => 
                           REGISTERS_10_13_port, B2 => n1701, ZN => n1189);
   U1640 : NAND4_X1 port map( A1 => n1192, A2 => n1191, A3 => n1190, A4 => 
                           n1189, ZN => n1193);
   U1641 : AOI22_X1 port map( A1 => n1194, A2 => n1725, B1 => n1193, B2 => 
                           n1721, ZN => n1195);
   U1642 : OAI221_X1 port map( B1 => n1733, B2 => n1197, C1 => n1729, C2 => 
                           n1196, A => n1195, ZN => N277);
   U1643 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n1616, B1 => 
                           REGISTERS_23_14_port, B2 => n1598, ZN => n1201);
   U1644 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n1652, B1 => 
                           REGISTERS_19_14_port, B2 => n1634, ZN => n1200);
   U1645 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n1688, B1 => 
                           REGISTERS_22_14_port, B2 => n1670, ZN => n1199);
   U1646 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n1715, B1 => 
                           REGISTERS_18_14_port, B2 => n1701, ZN => n1198);
   U1647 : AND4_X1 port map( A1 => n1201, A2 => n1200, A3 => n1199, A4 => n1198
                           , ZN => n1218);
   U1648 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n1616, B1 => 
                           REGISTERS_31_14_port, B2 => n1598, ZN => n1205);
   U1649 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n1652, B1 => 
                           REGISTERS_27_14_port, B2 => n1634, ZN => n1204);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n1688, B1 => 
                           REGISTERS_30_14_port, B2 => n1670, ZN => n1203);
   U1651 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n1715, B1 => 
                           REGISTERS_26_14_port, B2 => n1701, ZN => n1202);
   U1652 : AND4_X1 port map( A1 => n1205, A2 => n1204, A3 => n1203, A4 => n1202
                           , ZN => n1217);
   U1653 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n1616, B1 => 
                           REGISTERS_7_14_port, B2 => n1598, ZN => n1209);
   U1654 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n1652, B1 => 
                           REGISTERS_3_14_port, B2 => n1634, ZN => n1208);
   U1655 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n1688, B1 => 
                           REGISTERS_6_14_port, B2 => n1670, ZN => n1207);
   U1656 : NAND4_X1 port map( A1 => n1209, A2 => n1208, A3 => n1207, A4 => 
                           n1206, ZN => n1215);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n1616, B1 => 
                           REGISTERS_15_14_port, B2 => n1598, ZN => n1213);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n1652, B1 => 
                           REGISTERS_11_14_port, B2 => n1634, ZN => n1212);
   U1659 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n1688, B1 => 
                           REGISTERS_14_14_port, B2 => n1670, ZN => n1211);
   U1660 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n1714, B1 => 
                           REGISTERS_10_14_port, B2 => n1701, ZN => n1210);
   U1661 : NAND4_X1 port map( A1 => n1213, A2 => n1212, A3 => n1211, A4 => 
                           n1210, ZN => n1214);
   U1662 : AOI22_X1 port map( A1 => n1215, A2 => n1725, B1 => n1214, B2 => 
                           n1721, ZN => n1216);
   U1663 : OAI221_X1 port map( B1 => n1733, B2 => n1218, C1 => n1729, C2 => 
                           n1217, A => n1216, ZN => N276);
   U1664 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n1616, B1 => 
                           REGISTERS_23_15_port, B2 => n1598, ZN => n1222);
   U1665 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n1652, B1 => 
                           REGISTERS_19_15_port, B2 => n1634, ZN => n1221);
   U1666 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n1688, B1 => 
                           REGISTERS_22_15_port, B2 => n1670, ZN => n1220);
   U1667 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n1714, B1 => 
                           REGISTERS_18_15_port, B2 => n1701, ZN => n1219);
   U1668 : AND4_X1 port map( A1 => n1222, A2 => n1221, A3 => n1220, A4 => n1219
                           , ZN => n1239);
   U1669 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n1616, B1 => 
                           REGISTERS_31_15_port, B2 => n1598, ZN => n1226);
   U1670 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n1652, B1 => 
                           REGISTERS_27_15_port, B2 => n1634, ZN => n1225);
   U1671 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n1688, B1 => 
                           REGISTERS_30_15_port, B2 => n1670, ZN => n1224);
   U1672 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n1714, B1 => 
                           REGISTERS_26_15_port, B2 => n1700, ZN => n1223);
   U1673 : AND4_X1 port map( A1 => n1226, A2 => n1225, A3 => n1224, A4 => n1223
                           , ZN => n1238);
   U1674 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n1616, B1 => 
                           REGISTERS_7_15_port, B2 => n1598, ZN => n1230);
   U1675 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n1652, B1 => 
                           REGISTERS_3_15_port, B2 => n1634, ZN => n1229);
   U1676 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n1688, B1 => 
                           REGISTERS_6_15_port, B2 => n1670, ZN => n1228);
   U1677 : NAND4_X1 port map( A1 => n1230, A2 => n1229, A3 => n1228, A4 => 
                           n1227, ZN => n1236);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n1616, B1 => 
                           REGISTERS_15_15_port, B2 => n1598, ZN => n1234);
   U1679 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n1652, B1 => 
                           REGISTERS_11_15_port, B2 => n1634, ZN => n1233);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n1688, B1 => 
                           REGISTERS_14_15_port, B2 => n1670, ZN => n1232);
   U1681 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n1714, B1 => 
                           REGISTERS_10_15_port, B2 => n1700, ZN => n1231);
   U1682 : NAND4_X1 port map( A1 => n1234, A2 => n1233, A3 => n1232, A4 => 
                           n1231, ZN => n1235);
   U1683 : AOI22_X1 port map( A1 => n1236, A2 => n1725, B1 => n1235, B2 => 
                           n1721, ZN => n1237);
   U1684 : OAI221_X1 port map( B1 => n1733, B2 => n1239, C1 => n1729, C2 => 
                           n1238, A => n1237, ZN => N275);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n1616, B1 => 
                           REGISTERS_23_16_port, B2 => n1598, ZN => n1243);
   U1686 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n1652, B1 => 
                           REGISTERS_19_16_port, B2 => n1634, ZN => n1242);
   U1687 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n1688, B1 => 
                           REGISTERS_22_16_port, B2 => n1670, ZN => n1241);
   U1688 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n1714, B1 => 
                           REGISTERS_18_16_port, B2 => n1700, ZN => n1240);
   U1689 : AND4_X1 port map( A1 => n1243, A2 => n1242, A3 => n1241, A4 => n1240
                           , ZN => n1260);
   U1690 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n1616, B1 => 
                           REGISTERS_31_16_port, B2 => n1598, ZN => n1247);
   U1691 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n1652, B1 => 
                           REGISTERS_27_16_port, B2 => n1634, ZN => n1246);
   U1692 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n1688, B1 => 
                           REGISTERS_30_16_port, B2 => n1670, ZN => n1245);
   U1693 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n1714, B1 => 
                           REGISTERS_26_16_port, B2 => n1700, ZN => n1244);
   U1694 : AND4_X1 port map( A1 => n1247, A2 => n1246, A3 => n1245, A4 => n1244
                           , ZN => n1259);
   U1695 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n1615, B1 => 
                           REGISTERS_7_16_port, B2 => n1597, ZN => n1251);
   U1696 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n1651, B1 => 
                           REGISTERS_3_16_port, B2 => n1633, ZN => n1250);
   U1697 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n1687, B1 => 
                           REGISTERS_6_16_port, B2 => n1669, ZN => n1249);
   U1698 : NAND4_X1 port map( A1 => n1251, A2 => n1250, A3 => n1249, A4 => 
                           n1248, ZN => n1257);
   U1699 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n1615, B1 => 
                           REGISTERS_15_16_port, B2 => n1597, ZN => n1255);
   U1700 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n1651, B1 => 
                           REGISTERS_11_16_port, B2 => n1633, ZN => n1254);
   U1701 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n1687, B1 => 
                           REGISTERS_14_16_port, B2 => n1669, ZN => n1253);
   U1702 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n1714, B1 => 
                           REGISTERS_10_16_port, B2 => n1700, ZN => n1252);
   U1703 : NAND4_X1 port map( A1 => n1255, A2 => n1254, A3 => n1253, A4 => 
                           n1252, ZN => n1256);
   U1704 : AOI22_X1 port map( A1 => n1257, A2 => n1725, B1 => n1256, B2 => 
                           n1721, ZN => n1258);
   U1705 : OAI221_X1 port map( B1 => n1733, B2 => n1260, C1 => n1729, C2 => 
                           n1259, A => n1258, ZN => N274);
   U1706 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n1615, B1 => 
                           REGISTERS_23_17_port, B2 => n1597, ZN => n1264);
   U1707 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n1651, B1 => 
                           REGISTERS_19_17_port, B2 => n1633, ZN => n1263);
   U1708 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n1687, B1 => 
                           REGISTERS_22_17_port, B2 => n1669, ZN => n1262);
   U1709 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n1714, B1 => 
                           REGISTERS_18_17_port, B2 => n1700, ZN => n1261);
   U1710 : AND4_X1 port map( A1 => n1264, A2 => n1263, A3 => n1262, A4 => n1261
                           , ZN => n1281);
   U1711 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n1615, B1 => 
                           REGISTERS_31_17_port, B2 => n1597, ZN => n1268);
   U1712 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n1651, B1 => 
                           REGISTERS_27_17_port, B2 => n1633, ZN => n1267);
   U1713 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n1687, B1 => 
                           REGISTERS_30_17_port, B2 => n1669, ZN => n1266);
   U1714 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n1714, B1 => 
                           REGISTERS_26_17_port, B2 => n1700, ZN => n1265);
   U1715 : AND4_X1 port map( A1 => n1268, A2 => n1267, A3 => n1266, A4 => n1265
                           , ZN => n1280);
   U1716 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n1615, B1 => 
                           REGISTERS_7_17_port, B2 => n1597, ZN => n1272);
   U1717 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n1651, B1 => 
                           REGISTERS_3_17_port, B2 => n1633, ZN => n1271);
   U1718 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n1687, B1 => 
                           REGISTERS_6_17_port, B2 => n1669, ZN => n1270);
   U1719 : NAND4_X1 port map( A1 => n1272, A2 => n1271, A3 => n1270, A4 => 
                           n1269, ZN => n1278);
   U1720 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n1615, B1 => 
                           REGISTERS_15_17_port, B2 => n1597, ZN => n1276);
   U1721 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n1651, B1 => 
                           REGISTERS_11_17_port, B2 => n1633, ZN => n1275);
   U1722 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n1687, B1 => 
                           REGISTERS_14_17_port, B2 => n1669, ZN => n1274);
   U1723 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n1714, B1 => 
                           REGISTERS_10_17_port, B2 => n1700, ZN => n1273);
   U1724 : NAND4_X1 port map( A1 => n1276, A2 => n1275, A3 => n1274, A4 => 
                           n1273, ZN => n1277);
   U1725 : AOI22_X1 port map( A1 => n1278, A2 => n1725, B1 => n1277, B2 => 
                           n1721, ZN => n1279);
   U1726 : OAI221_X1 port map( B1 => n1733, B2 => n1281, C1 => n1729, C2 => 
                           n1280, A => n1279, ZN => N273);
   U1727 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n1615, B1 => 
                           REGISTERS_23_18_port, B2 => n1597, ZN => n1285);
   U1728 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n1651, B1 => 
                           REGISTERS_19_18_port, B2 => n1633, ZN => n1284);
   U1729 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n1687, B1 => 
                           REGISTERS_22_18_port, B2 => n1669, ZN => n1283);
   U1730 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n1714, B1 => 
                           REGISTERS_18_18_port, B2 => n1700, ZN => n1282);
   U1731 : AND4_X1 port map( A1 => n1285, A2 => n1284, A3 => n1283, A4 => n1282
                           , ZN => n1302);
   U1732 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n1615, B1 => 
                           REGISTERS_31_18_port, B2 => n1597, ZN => n1289);
   U1733 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n1651, B1 => 
                           REGISTERS_27_18_port, B2 => n1633, ZN => n1288);
   U1734 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n1687, B1 => 
                           REGISTERS_30_18_port, B2 => n1669, ZN => n1287);
   U1735 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n1713, B1 => 
                           REGISTERS_26_18_port, B2 => n1700, ZN => n1286);
   U1736 : AND4_X1 port map( A1 => n1289, A2 => n1288, A3 => n1287, A4 => n1286
                           , ZN => n1301);
   U1737 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n1615, B1 => 
                           REGISTERS_7_18_port, B2 => n1597, ZN => n1293);
   U1738 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n1651, B1 => 
                           REGISTERS_3_18_port, B2 => n1633, ZN => n1292);
   U1739 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n1687, B1 => 
                           REGISTERS_6_18_port, B2 => n1669, ZN => n1291);
   U1740 : NAND4_X1 port map( A1 => n1293, A2 => n1292, A3 => n1291, A4 => 
                           n1290, ZN => n1299);
   U1741 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n1615, B1 => 
                           REGISTERS_15_18_port, B2 => n1597, ZN => n1297);
   U1742 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n1651, B1 => 
                           REGISTERS_11_18_port, B2 => n1633, ZN => n1296);
   U1743 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n1687, B1 => 
                           REGISTERS_14_18_port, B2 => n1669, ZN => n1295);
   U1744 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n1713, B1 => 
                           REGISTERS_10_18_port, B2 => n1700, ZN => n1294);
   U1745 : NAND4_X1 port map( A1 => n1297, A2 => n1296, A3 => n1295, A4 => 
                           n1294, ZN => n1298);
   U1746 : AOI22_X1 port map( A1 => n1299, A2 => n1725, B1 => n1298, B2 => 
                           n1721, ZN => n1300);
   U1747 : OAI221_X1 port map( B1 => n1733, B2 => n1302, C1 => n1729, C2 => 
                           n1301, A => n1300, ZN => N272);
   U1748 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n1615, B1 => 
                           REGISTERS_23_19_port, B2 => n1597, ZN => n1306);
   U1749 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n1651, B1 => 
                           REGISTERS_19_19_port, B2 => n1633, ZN => n1305);
   U1750 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n1687, B1 => 
                           REGISTERS_22_19_port, B2 => n1669, ZN => n1304);
   U1751 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n1713, B1 => 
                           REGISTERS_18_19_port, B2 => n1700, ZN => n1303);
   U1752 : AND4_X1 port map( A1 => n1306, A2 => n1305, A3 => n1304, A4 => n1303
                           , ZN => n1323);
   U1753 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n1614, B1 => 
                           REGISTERS_31_19_port, B2 => n1596, ZN => n1310);
   U1754 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n1650, B1 => 
                           REGISTERS_27_19_port, B2 => n1632, ZN => n1309);
   U1755 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n1686, B1 => 
                           REGISTERS_30_19_port, B2 => n1668, ZN => n1308);
   U1756 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n1713, B1 => 
                           REGISTERS_26_19_port, B2 => n1700, ZN => n1307);
   U1757 : AND4_X1 port map( A1 => n1310, A2 => n1309, A3 => n1308, A4 => n1307
                           , ZN => n1322);
   U1758 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n1614, B1 => 
                           REGISTERS_7_19_port, B2 => n1596, ZN => n1314);
   U1759 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n1650, B1 => 
                           REGISTERS_3_19_port, B2 => n1632, ZN => n1313);
   U1760 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n1686, B1 => 
                           REGISTERS_6_19_port, B2 => n1668, ZN => n1312);
   U1761 : NAND4_X1 port map( A1 => n1314, A2 => n1313, A3 => n1312, A4 => 
                           n1311, ZN => n1320);
   U1762 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n1614, B1 => 
                           REGISTERS_15_19_port, B2 => n1596, ZN => n1318);
   U1763 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n1650, B1 => 
                           REGISTERS_11_19_port, B2 => n1632, ZN => n1317);
   U1764 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n1686, B1 => 
                           REGISTERS_14_19_port, B2 => n1668, ZN => n1316);
   U1765 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n1713, B1 => 
                           REGISTERS_10_19_port, B2 => n1700, ZN => n1315);
   U1766 : NAND4_X1 port map( A1 => n1318, A2 => n1317, A3 => n1316, A4 => 
                           n1315, ZN => n1319);
   U1767 : AOI22_X1 port map( A1 => n1320, A2 => n1725, B1 => n1319, B2 => 
                           n1721, ZN => n1321);
   U1768 : OAI221_X1 port map( B1 => n1733, B2 => n1323, C1 => n1729, C2 => 
                           n1322, A => n1321, ZN => N271);
   U1769 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n1614, B1 => 
                           REGISTERS_23_20_port, B2 => n1596, ZN => n1327);
   U1770 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n1650, B1 => 
                           REGISTERS_19_20_port, B2 => n1632, ZN => n1326);
   U1771 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n1686, B1 => 
                           REGISTERS_22_20_port, B2 => n1668, ZN => n1325);
   U1772 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n1713, B1 => 
                           REGISTERS_18_20_port, B2 => n1700, ZN => n1324);
   U1773 : AND4_X1 port map( A1 => n1327, A2 => n1326, A3 => n1325, A4 => n1324
                           , ZN => n1344);
   U1774 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n1614, B1 => 
                           REGISTERS_31_20_port, B2 => n1596, ZN => n1331);
   U1775 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n1650, B1 => 
                           REGISTERS_27_20_port, B2 => n1632, ZN => n1330);
   U1776 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n1686, B1 => 
                           REGISTERS_30_20_port, B2 => n1668, ZN => n1329);
   U1777 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n1713, B1 => 
                           REGISTERS_26_20_port, B2 => n1700, ZN => n1328);
   U1778 : AND4_X1 port map( A1 => n1331, A2 => n1330, A3 => n1329, A4 => n1328
                           , ZN => n1343);
   U1779 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n1614, B1 => 
                           REGISTERS_7_20_port, B2 => n1596, ZN => n1335);
   U1780 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n1650, B1 => 
                           REGISTERS_3_20_port, B2 => n1632, ZN => n1334);
   U1781 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n1686, B1 => 
                           REGISTERS_6_20_port, B2 => n1668, ZN => n1333);
   U1782 : NAND4_X1 port map( A1 => n1335, A2 => n1334, A3 => n1333, A4 => 
                           n1332, ZN => n1341);
   U1783 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n1614, B1 => 
                           REGISTERS_15_20_port, B2 => n1596, ZN => n1339);
   U1784 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n1650, B1 => 
                           REGISTERS_11_20_port, B2 => n1632, ZN => n1338);
   U1785 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n1686, B1 => 
                           REGISTERS_14_20_port, B2 => n1668, ZN => n1337);
   U1786 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n1713, B1 => 
                           REGISTERS_10_20_port, B2 => n1700, ZN => n1336);
   U1787 : NAND4_X1 port map( A1 => n1339, A2 => n1338, A3 => n1337, A4 => 
                           n1336, ZN => n1340);
   U1788 : AOI22_X1 port map( A1 => n1341, A2 => n1725, B1 => n1340, B2 => 
                           n1721, ZN => n1342);
   U1789 : OAI221_X1 port map( B1 => n1733, B2 => n1344, C1 => n1729, C2 => 
                           n1343, A => n1342, ZN => N270);
   U1790 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n1614, B1 => 
                           REGISTERS_23_21_port, B2 => n1596, ZN => n1348);
   U1791 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n1650, B1 => 
                           REGISTERS_19_21_port, B2 => n1632, ZN => n1347);
   U1792 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n1686, B1 => 
                           REGISTERS_22_21_port, B2 => n1668, ZN => n1346);
   U1793 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n1713, B1 => 
                           REGISTERS_18_21_port, B2 => n1700, ZN => n1345);
   U1794 : AND4_X1 port map( A1 => n1348, A2 => n1347, A3 => n1346, A4 => n1345
                           , ZN => n1365);
   U1795 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n1614, B1 => 
                           REGISTERS_31_21_port, B2 => n1596, ZN => n1352);
   U1796 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n1650, B1 => 
                           REGISTERS_27_21_port, B2 => n1632, ZN => n1351);
   U1797 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n1686, B1 => 
                           REGISTERS_30_21_port, B2 => n1668, ZN => n1350);
   U1798 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n1713, B1 => 
                           REGISTERS_26_21_port, B2 => n1700, ZN => n1349);
   U1799 : AND4_X1 port map( A1 => n1352, A2 => n1351, A3 => n1350, A4 => n1349
                           , ZN => n1364);
   U1800 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n1614, B1 => 
                           REGISTERS_7_21_port, B2 => n1596, ZN => n1356);
   U1801 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n1650, B1 => 
                           REGISTERS_3_21_port, B2 => n1632, ZN => n1355);
   U1802 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n1686, B1 => 
                           REGISTERS_6_21_port, B2 => n1668, ZN => n1354);
   U1803 : NAND4_X1 port map( A1 => n1356, A2 => n1355, A3 => n1354, A4 => 
                           n1353, ZN => n1362);
   U1804 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n1614, B1 => 
                           REGISTERS_15_21_port, B2 => n1596, ZN => n1360);
   U1805 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n1650, B1 => 
                           REGISTERS_11_21_port, B2 => n1632, ZN => n1359);
   U1806 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n1686, B1 => 
                           REGISTERS_14_21_port, B2 => n1668, ZN => n1358);
   U1807 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n1713, B1 => 
                           REGISTERS_10_21_port, B2 => n1700, ZN => n1357);
   U1808 : NAND4_X1 port map( A1 => n1360, A2 => n1359, A3 => n1358, A4 => 
                           n1357, ZN => n1361);
   U1809 : AOI22_X1 port map( A1 => n1362, A2 => n1725, B1 => n1361, B2 => 
                           n1721, ZN => n1363);
   U1810 : OAI221_X1 port map( B1 => n1733, B2 => n1365, C1 => n1730, C2 => 
                           n1364, A => n1363, ZN => N269);
   U1811 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n1613, B1 => 
                           REGISTERS_23_22_port, B2 => n1595, ZN => n1369);
   U1812 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n1649, B1 => 
                           REGISTERS_19_22_port, B2 => n1631, ZN => n1368);
   U1813 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n1685, B1 => 
                           REGISTERS_22_22_port, B2 => n1667, ZN => n1367);
   U1814 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n1712, B1 => 
                           REGISTERS_18_22_port, B2 => n1699, ZN => n1366);
   U1815 : AND4_X1 port map( A1 => n1369, A2 => n1368, A3 => n1367, A4 => n1366
                           , ZN => n1386);
   U1816 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n1613, B1 => 
                           REGISTERS_31_22_port, B2 => n1595, ZN => n1373);
   U1817 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n1649, B1 => 
                           REGISTERS_27_22_port, B2 => n1631, ZN => n1372);
   U1818 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n1685, B1 => 
                           REGISTERS_30_22_port, B2 => n1667, ZN => n1371);
   U1819 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n1712, B1 => 
                           REGISTERS_26_22_port, B2 => n1699, ZN => n1370);
   U1820 : AND4_X1 port map( A1 => n1373, A2 => n1372, A3 => n1371, A4 => n1370
                           , ZN => n1385);
   U1821 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n1613, B1 => 
                           REGISTERS_7_22_port, B2 => n1595, ZN => n1377);
   U1822 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n1649, B1 => 
                           REGISTERS_3_22_port, B2 => n1631, ZN => n1376);
   U1823 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n1685, B1 => 
                           REGISTERS_6_22_port, B2 => n1667, ZN => n1375);
   U1824 : NAND4_X1 port map( A1 => n1377, A2 => n1376, A3 => n1375, A4 => 
                           n1374, ZN => n1383);
   U1825 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n1613, B1 => 
                           REGISTERS_15_22_port, B2 => n1595, ZN => n1381);
   U1826 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n1649, B1 => 
                           REGISTERS_11_22_port, B2 => n1631, ZN => n1380);
   U1827 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n1685, B1 => 
                           REGISTERS_14_22_port, B2 => n1667, ZN => n1379);
   U1828 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n1712, B1 => 
                           REGISTERS_10_22_port, B2 => n1699, ZN => n1378);
   U1829 : NAND4_X1 port map( A1 => n1381, A2 => n1380, A3 => n1379, A4 => 
                           n1378, ZN => n1382);
   U1830 : AOI22_X1 port map( A1 => n1383, A2 => n1724, B1 => n1382, B2 => 
                           n1720, ZN => n1384);
   U1831 : OAI221_X1 port map( B1 => n1732, B2 => n1386, C1 => n1730, C2 => 
                           n1385, A => n1384, ZN => N268);
   U1832 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n1613, B1 => 
                           REGISTERS_23_23_port, B2 => n1595, ZN => n1390);
   U1833 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n1649, B1 => 
                           REGISTERS_19_23_port, B2 => n1631, ZN => n1389);
   U1834 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n1685, B1 => 
                           REGISTERS_22_23_port, B2 => n1667, ZN => n1388);
   U1835 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n1712, B1 => 
                           REGISTERS_18_23_port, B2 => n1699, ZN => n1387);
   U1836 : AND4_X1 port map( A1 => n1390, A2 => n1389, A3 => n1388, A4 => n1387
                           , ZN => n1407);
   U1837 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n1613, B1 => 
                           REGISTERS_31_23_port, B2 => n1595, ZN => n1394);
   U1838 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n1649, B1 => 
                           REGISTERS_27_23_port, B2 => n1631, ZN => n1393);
   U1839 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n1685, B1 => 
                           REGISTERS_30_23_port, B2 => n1667, ZN => n1392);
   U1840 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n1712, B1 => 
                           REGISTERS_26_23_port, B2 => n1699, ZN => n1391);
   U1841 : AND4_X1 port map( A1 => n1394, A2 => n1393, A3 => n1392, A4 => n1391
                           , ZN => n1406);
   U1842 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n1613, B1 => 
                           REGISTERS_7_23_port, B2 => n1595, ZN => n1398);
   U1843 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n1649, B1 => 
                           REGISTERS_3_23_port, B2 => n1631, ZN => n1397);
   U1844 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n1685, B1 => 
                           REGISTERS_6_23_port, B2 => n1667, ZN => n1396);
   U1845 : NAND4_X1 port map( A1 => n1398, A2 => n1397, A3 => n1396, A4 => 
                           n1395, ZN => n1404);
   U1846 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n1613, B1 => 
                           REGISTERS_15_23_port, B2 => n1595, ZN => n1402);
   U1847 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n1649, B1 => 
                           REGISTERS_11_23_port, B2 => n1631, ZN => n1401);
   U1848 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n1685, B1 => 
                           REGISTERS_14_23_port, B2 => n1667, ZN => n1400);
   U1849 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n1712, B1 => 
                           REGISTERS_10_23_port, B2 => n1699, ZN => n1399);
   U1850 : NAND4_X1 port map( A1 => n1402, A2 => n1401, A3 => n1400, A4 => 
                           n1399, ZN => n1403);
   U1851 : AOI22_X1 port map( A1 => n1404, A2 => n1724, B1 => n1403, B2 => 
                           n1720, ZN => n1405);
   U1852 : OAI221_X1 port map( B1 => n1732, B2 => n1407, C1 => n1730, C2 => 
                           n1406, A => n1405, ZN => N267);
   U1853 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n1613, B1 => 
                           REGISTERS_23_24_port, B2 => n1595, ZN => n1411);
   U1854 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n1649, B1 => 
                           REGISTERS_19_24_port, B2 => n1631, ZN => n1410);
   U1855 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n1685, B1 => 
                           REGISTERS_22_24_port, B2 => n1667, ZN => n1409);
   U1856 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n1712, B1 => 
                           REGISTERS_18_24_port, B2 => n1699, ZN => n1408);
   U1857 : AND4_X1 port map( A1 => n1411, A2 => n1410, A3 => n1409, A4 => n1408
                           , ZN => n1428);
   U1858 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n1613, B1 => 
                           REGISTERS_31_24_port, B2 => n1595, ZN => n1415);
   U1859 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n1649, B1 => 
                           REGISTERS_27_24_port, B2 => n1631, ZN => n1414);
   U1860 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n1685, B1 => 
                           REGISTERS_30_24_port, B2 => n1667, ZN => n1413);
   U1861 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n1712, B1 => 
                           REGISTERS_26_24_port, B2 => n1699, ZN => n1412);
   U1862 : AND4_X1 port map( A1 => n1415, A2 => n1414, A3 => n1413, A4 => n1412
                           , ZN => n1427);
   U1863 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n1613, B1 => 
                           REGISTERS_7_24_port, B2 => n1595, ZN => n1419);
   U1864 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n1649, B1 => 
                           REGISTERS_3_24_port, B2 => n1631, ZN => n1418);
   U1865 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n1685, B1 => 
                           REGISTERS_6_24_port, B2 => n1667, ZN => n1417);
   U1866 : NAND4_X1 port map( A1 => n1419, A2 => n1418, A3 => n1417, A4 => 
                           n1416, ZN => n1425);
   U1867 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n1612, B1 => 
                           REGISTERS_15_24_port, B2 => n1594, ZN => n1423);
   U1868 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n1648, B1 => 
                           REGISTERS_11_24_port, B2 => n1630, ZN => n1422);
   U1869 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n1684, B1 => 
                           REGISTERS_14_24_port, B2 => n1666, ZN => n1421);
   U1870 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n1712, B1 => 
                           REGISTERS_10_24_port, B2 => n1699, ZN => n1420);
   U1871 : NAND4_X1 port map( A1 => n1423, A2 => n1422, A3 => n1421, A4 => 
                           n1420, ZN => n1424);
   U1872 : AOI22_X1 port map( A1 => n1425, A2 => n1724, B1 => n1424, B2 => 
                           n1720, ZN => n1426);
   U1873 : OAI221_X1 port map( B1 => n1732, B2 => n1428, C1 => n1730, C2 => 
                           n1427, A => n1426, ZN => N266);
   U1874 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n1612, B1 => 
                           REGISTERS_23_25_port, B2 => n1594, ZN => n1432);
   U1875 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n1648, B1 => 
                           REGISTERS_19_25_port, B2 => n1630, ZN => n1431);
   U1876 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n1684, B1 => 
                           REGISTERS_22_25_port, B2 => n1666, ZN => n1430);
   U1877 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n1712, B1 => 
                           REGISTERS_18_25_port, B2 => n1699, ZN => n1429);
   U1878 : AND4_X1 port map( A1 => n1432, A2 => n1431, A3 => n1430, A4 => n1429
                           , ZN => n1449);
   U1879 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n1612, B1 => 
                           REGISTERS_31_25_port, B2 => n1594, ZN => n1436);
   U1880 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n1648, B1 => 
                           REGISTERS_27_25_port, B2 => n1630, ZN => n1435);
   U1881 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n1684, B1 => 
                           REGISTERS_30_25_port, B2 => n1666, ZN => n1434);
   U1882 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n1712, B1 => 
                           REGISTERS_26_25_port, B2 => n1699, ZN => n1433);
   U1883 : AND4_X1 port map( A1 => n1436, A2 => n1435, A3 => n1434, A4 => n1433
                           , ZN => n1448);
   U1884 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n1612, B1 => 
                           REGISTERS_7_25_port, B2 => n1594, ZN => n1440);
   U1885 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n1648, B1 => 
                           REGISTERS_3_25_port, B2 => n1630, ZN => n1439);
   U1886 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n1684, B1 => 
                           REGISTERS_6_25_port, B2 => n1666, ZN => n1438);
   U1887 : NAND4_X1 port map( A1 => n1440, A2 => n1439, A3 => n1438, A4 => 
                           n1437, ZN => n1446);
   U1888 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n1612, B1 => 
                           REGISTERS_15_25_port, B2 => n1594, ZN => n1444);
   U1889 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n1648, B1 => 
                           REGISTERS_11_25_port, B2 => n1630, ZN => n1443);
   U1890 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n1684, B1 => 
                           REGISTERS_14_25_port, B2 => n1666, ZN => n1442);
   U1891 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n1711, B1 => 
                           REGISTERS_10_25_port, B2 => n1699, ZN => n1441);
   U1892 : NAND4_X1 port map( A1 => n1444, A2 => n1443, A3 => n1442, A4 => 
                           n1441, ZN => n1445);
   U1893 : AOI22_X1 port map( A1 => n1446, A2 => n1724, B1 => n1445, B2 => 
                           n1720, ZN => n1447);
   U1894 : OAI221_X1 port map( B1 => n1732, B2 => n1449, C1 => n1730, C2 => 
                           n1448, A => n1447, ZN => N265);
   U1895 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n1612, B1 => 
                           REGISTERS_23_26_port, B2 => n1594, ZN => n1453);
   U1896 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n1648, B1 => 
                           REGISTERS_19_26_port, B2 => n1630, ZN => n1452);
   U1897 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n1684, B1 => 
                           REGISTERS_22_26_port, B2 => n1666, ZN => n1451);
   U1898 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n1711, B1 => 
                           REGISTERS_18_26_port, B2 => n1699, ZN => n1450);
   U1899 : AND4_X1 port map( A1 => n1453, A2 => n1452, A3 => n1451, A4 => n1450
                           , ZN => n1470);
   U1900 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n1612, B1 => 
                           REGISTERS_31_26_port, B2 => n1594, ZN => n1457);
   U1901 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n1648, B1 => 
                           REGISTERS_27_26_port, B2 => n1630, ZN => n1456);
   U1902 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n1684, B1 => 
                           REGISTERS_30_26_port, B2 => n1666, ZN => n1455);
   U1903 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n1711, B1 => 
                           REGISTERS_26_26_port, B2 => n1699, ZN => n1454);
   U1904 : AND4_X1 port map( A1 => n1457, A2 => n1456, A3 => n1455, A4 => n1454
                           , ZN => n1469);
   U1905 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n1612, B1 => 
                           REGISTERS_7_26_port, B2 => n1594, ZN => n1461);
   U1906 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n1648, B1 => 
                           REGISTERS_3_26_port, B2 => n1630, ZN => n1460);
   U1907 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n1684, B1 => 
                           REGISTERS_6_26_port, B2 => n1666, ZN => n1459);
   U1908 : NAND4_X1 port map( A1 => n1461, A2 => n1460, A3 => n1459, A4 => 
                           n1458, ZN => n1467);
   U1909 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n1612, B1 => 
                           REGISTERS_15_26_port, B2 => n1594, ZN => n1465);
   U1910 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n1648, B1 => 
                           REGISTERS_11_26_port, B2 => n1630, ZN => n1464);
   U1911 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n1684, B1 => 
                           REGISTERS_14_26_port, B2 => n1666, ZN => n1463);
   U1912 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n1711, B1 => 
                           REGISTERS_10_26_port, B2 => n1699, ZN => n1462);
   U1913 : NAND4_X1 port map( A1 => n1465, A2 => n1464, A3 => n1463, A4 => 
                           n1462, ZN => n1466);
   U1914 : AOI22_X1 port map( A1 => n1467, A2 => n1724, B1 => n1466, B2 => 
                           n1720, ZN => n1468);
   U1915 : OAI221_X1 port map( B1 => n1732, B2 => n1470, C1 => n1730, C2 => 
                           n1469, A => n1468, ZN => N264);
   U1916 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n1612, B1 => 
                           REGISTERS_23_27_port, B2 => n1594, ZN => n1474);
   U1917 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n1648, B1 => 
                           REGISTERS_19_27_port, B2 => n1630, ZN => n1473);
   U1918 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n1684, B1 => 
                           REGISTERS_22_27_port, B2 => n1666, ZN => n1472);
   U1919 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n1711, B1 => 
                           REGISTERS_18_27_port, B2 => n1699, ZN => n1471);
   U1920 : AND4_X1 port map( A1 => n1474, A2 => n1473, A3 => n1472, A4 => n1471
                           , ZN => n1491);
   U1921 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n1612, B1 => 
                           REGISTERS_31_27_port, B2 => n1594, ZN => n1478);
   U1922 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n1648, B1 => 
                           REGISTERS_27_27_port, B2 => n1630, ZN => n1477);
   U1923 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n1684, B1 => 
                           REGISTERS_30_27_port, B2 => n1666, ZN => n1476);
   U1924 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n1711, B1 => 
                           REGISTERS_26_27_port, B2 => n1699, ZN => n1475);
   U1925 : AND4_X1 port map( A1 => n1478, A2 => n1477, A3 => n1476, A4 => n1475
                           , ZN => n1490);
   U1926 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n1611, B1 => 
                           REGISTERS_7_27_port, B2 => n1593, ZN => n1482);
   U1927 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n1647, B1 => 
                           REGISTERS_3_27_port, B2 => n1629, ZN => n1481);
   U1928 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n1683, B1 => 
                           REGISTERS_6_27_port, B2 => n1665, ZN => n1480);
   U1929 : NAND4_X1 port map( A1 => n1482, A2 => n1481, A3 => n1480, A4 => 
                           n1479, ZN => n1488);
   U1930 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n1611, B1 => 
                           REGISTERS_15_27_port, B2 => n1593, ZN => n1486);
   U1931 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n1647, B1 => 
                           REGISTERS_11_27_port, B2 => n1629, ZN => n1485);
   U1932 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n1683, B1 => 
                           REGISTERS_14_27_port, B2 => n1665, ZN => n1484);
   U1933 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n1711, B1 => 
                           REGISTERS_10_27_port, B2 => n1699, ZN => n1483);
   U1934 : NAND4_X1 port map( A1 => n1486, A2 => n1485, A3 => n1484, A4 => 
                           n1483, ZN => n1487);
   U1935 : AOI22_X1 port map( A1 => n1488, A2 => n1724, B1 => n1487, B2 => 
                           n1720, ZN => n1489);
   U1936 : OAI221_X1 port map( B1 => n1732, B2 => n1491, C1 => n1730, C2 => 
                           n1490, A => n1489, ZN => N263);
   U1937 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n1611, B1 => 
                           REGISTERS_23_28_port, B2 => n1593, ZN => n1495);
   U1938 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n1647, B1 => 
                           REGISTERS_19_28_port, B2 => n1629, ZN => n1494);
   U1939 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n1683, B1 => 
                           REGISTERS_22_28_port, B2 => n1665, ZN => n1493);
   U1940 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n1711, B1 => 
                           REGISTERS_18_28_port, B2 => n1699, ZN => n1492);
   U1941 : AND4_X1 port map( A1 => n1495, A2 => n1494, A3 => n1493, A4 => n1492
                           , ZN => n1512);
   U1942 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n1611, B1 => 
                           REGISTERS_31_28_port, B2 => n1593, ZN => n1499);
   U1943 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n1647, B1 => 
                           REGISTERS_27_28_port, B2 => n1629, ZN => n1498);
   U1944 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n1683, B1 => 
                           REGISTERS_30_28_port, B2 => n1665, ZN => n1497);
   U1945 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n1711, B1 => 
                           REGISTERS_26_28_port, B2 => n1699, ZN => n1496);
   U1946 : AND4_X1 port map( A1 => n1499, A2 => n1498, A3 => n1497, A4 => n1496
                           , ZN => n1511);
   U1947 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n1611, B1 => 
                           REGISTERS_7_28_port, B2 => n1593, ZN => n1503);
   U1948 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n1647, B1 => 
                           REGISTERS_3_28_port, B2 => n1629, ZN => n1502);
   U1949 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n1683, B1 => 
                           REGISTERS_6_28_port, B2 => n1665, ZN => n1501);
   U1950 : NAND4_X1 port map( A1 => n1503, A2 => n1502, A3 => n1501, A4 => 
                           n1500, ZN => n1509);
   U1951 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n1611, B1 => 
                           REGISTERS_15_28_port, B2 => n1593, ZN => n1507);
   U1952 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n1647, B1 => 
                           REGISTERS_11_28_port, B2 => n1629, ZN => n1506);
   U1953 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n1683, B1 => 
                           REGISTERS_14_28_port, B2 => n1665, ZN => n1505);
   U1954 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n1711, B1 => 
                           REGISTERS_10_28_port, B2 => n1698, ZN => n1504);
   U1955 : NAND4_X1 port map( A1 => n1507, A2 => n1506, A3 => n1505, A4 => 
                           n1504, ZN => n1508);
   U1956 : AOI22_X1 port map( A1 => n1509, A2 => n1724, B1 => n1508, B2 => 
                           n1720, ZN => n1510);
   U1957 : OAI221_X1 port map( B1 => n1732, B2 => n1512, C1 => n1730, C2 => 
                           n1511, A => n1510, ZN => N262);
   U1958 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n1611, B1 => 
                           REGISTERS_23_29_port, B2 => n1593, ZN => n1516);
   U1959 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n1647, B1 => 
                           REGISTERS_19_29_port, B2 => n1629, ZN => n1515);
   U1960 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n1683, B1 => 
                           REGISTERS_22_29_port, B2 => n1665, ZN => n1514);
   U1961 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n1711, B1 => 
                           REGISTERS_18_29_port, B2 => n1698, ZN => n1513);
   U1962 : AND4_X1 port map( A1 => n1516, A2 => n1515, A3 => n1514, A4 => n1513
                           , ZN => n1533);
   U1963 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n1611, B1 => 
                           REGISTERS_31_29_port, B2 => n1593, ZN => n1520);
   U1964 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n1647, B1 => 
                           REGISTERS_27_29_port, B2 => n1629, ZN => n1519);
   U1965 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n1683, B1 => 
                           REGISTERS_30_29_port, B2 => n1665, ZN => n1518);
   U1966 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n1710, B1 => 
                           REGISTERS_26_29_port, B2 => n1698, ZN => n1517);
   U1967 : AND4_X1 port map( A1 => n1520, A2 => n1519, A3 => n1518, A4 => n1517
                           , ZN => n1532);
   U1968 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n1611, B1 => 
                           REGISTERS_7_29_port, B2 => n1593, ZN => n1524);
   U1969 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n1647, B1 => 
                           REGISTERS_3_29_port, B2 => n1629, ZN => n1523);
   U1970 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n1683, B1 => 
                           REGISTERS_6_29_port, B2 => n1665, ZN => n1522);
   U1971 : NAND4_X1 port map( A1 => n1524, A2 => n1523, A3 => n1522, A4 => 
                           n1521, ZN => n1530);
   U1972 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n1611, B1 => 
                           REGISTERS_15_29_port, B2 => n1593, ZN => n1528);
   U1973 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n1647, B1 => 
                           REGISTERS_11_29_port, B2 => n1629, ZN => n1527);
   U1974 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n1683, B1 => 
                           REGISTERS_14_29_port, B2 => n1665, ZN => n1526);
   U1975 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n1710, B1 => 
                           REGISTERS_10_29_port, B2 => n1698, ZN => n1525);
   U1976 : NAND4_X1 port map( A1 => n1528, A2 => n1527, A3 => n1526, A4 => 
                           n1525, ZN => n1529);
   U1977 : AOI22_X1 port map( A1 => n1530, A2 => n1724, B1 => n1529, B2 => 
                           n1720, ZN => n1531);
   U1978 : OAI221_X1 port map( B1 => n1732, B2 => n1533, C1 => n1730, C2 => 
                           n1532, A => n1531, ZN => N261);
   U1979 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n1611, B1 => 
                           REGISTERS_23_30_port, B2 => n1593, ZN => n1537);
   U1980 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n1647, B1 => 
                           REGISTERS_19_30_port, B2 => n1629, ZN => n1536);
   U1981 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n1683, B1 => 
                           REGISTERS_22_30_port, B2 => n1665, ZN => n1535);
   U1982 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n1710, B1 => 
                           REGISTERS_18_30_port, B2 => n1698, ZN => n1534);
   U1983 : AND4_X1 port map( A1 => n1537, A2 => n1536, A3 => n1535, A4 => n1534
                           , ZN => n1554);
   U1984 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n1610, B1 => 
                           REGISTERS_31_30_port, B2 => n1592, ZN => n1541);
   U1985 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n1646, B1 => 
                           REGISTERS_27_30_port, B2 => n1628, ZN => n1540);
   U1986 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n1682, B1 => 
                           REGISTERS_30_30_port, B2 => n1664, ZN => n1539);
   U1987 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n1710, B1 => 
                           REGISTERS_26_30_port, B2 => n1698, ZN => n1538);
   U1988 : AND4_X1 port map( A1 => n1541, A2 => n1540, A3 => n1539, A4 => n1538
                           , ZN => n1553);
   U1989 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n1610, B1 => 
                           REGISTERS_7_30_port, B2 => n1592, ZN => n1545);
   U1990 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n1646, B1 => 
                           REGISTERS_3_30_port, B2 => n1628, ZN => n1544);
   U1991 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n1682, B1 => 
                           REGISTERS_6_30_port, B2 => n1664, ZN => n1543);
   U1992 : NAND4_X1 port map( A1 => n1545, A2 => n1544, A3 => n1543, A4 => 
                           n1542, ZN => n1551);
   U1993 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n1610, B1 => 
                           REGISTERS_15_30_port, B2 => n1592, ZN => n1549);
   U1994 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n1646, B1 => 
                           REGISTERS_11_30_port, B2 => n1628, ZN => n1548);
   U1995 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n1682, B1 => 
                           REGISTERS_14_30_port, B2 => n1664, ZN => n1547);
   U1996 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n1710, B1 => 
                           REGISTERS_10_30_port, B2 => n1698, ZN => n1546);
   U1997 : NAND4_X1 port map( A1 => n1549, A2 => n1548, A3 => n1547, A4 => 
                           n1546, ZN => n1550);
   U1998 : AOI22_X1 port map( A1 => n1551, A2 => n1724, B1 => n1550, B2 => 
                           n1720, ZN => n1552);
   U1999 : OAI221_X1 port map( B1 => n1732, B2 => n1554, C1 => n1730, C2 => 
                           n1553, A => n1552, ZN => N260);
   U2000 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n1610, B1 => 
                           REGISTERS_23_31_port, B2 => n1592, ZN => n1558);
   U2001 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n1646, B1 => 
                           REGISTERS_19_31_port, B2 => n1628, ZN => n1557);
   U2002 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n1682, B1 => 
                           REGISTERS_22_31_port, B2 => n1664, ZN => n1556);
   U2003 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n1710, B1 => 
                           REGISTERS_18_31_port, B2 => n1698, ZN => n1555);
   U2004 : AND4_X1 port map( A1 => n1558, A2 => n1557, A3 => n1556, A4 => n1555
                           , ZN => n1581);
   U2005 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n1610, B1 => 
                           REGISTERS_31_31_port, B2 => n1592, ZN => n1562);
   U2006 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n1646, B1 => 
                           REGISTERS_27_31_port, B2 => n1628, ZN => n1561);
   U2007 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n1682, B1 => 
                           REGISTERS_30_31_port, B2 => n1664, ZN => n1560);
   U2008 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n1710, B1 => 
                           REGISTERS_26_31_port, B2 => n1698, ZN => n1559);
   U2009 : AND4_X1 port map( A1 => n1562, A2 => n1561, A3 => n1560, A4 => n1559
                           , ZN => n1579);
   U2010 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n1610, B1 => 
                           REGISTERS_7_31_port, B2 => n1592, ZN => n1566);
   U2011 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n1646, B1 => 
                           REGISTERS_3_31_port, B2 => n1628, ZN => n1565);
   U2012 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n1682, B1 => 
                           REGISTERS_6_31_port, B2 => n1664, ZN => n1564);
   U2013 : NAND4_X1 port map( A1 => n1566, A2 => n1565, A3 => n1564, A4 => 
                           n1563, ZN => n1575);
   U2014 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n1610, B1 => 
                           REGISTERS_15_31_port, B2 => n1592, ZN => n1572);
   U2015 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n1646, B1 => 
                           REGISTERS_11_31_port, B2 => n1628, ZN => n1571);
   U2016 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n1682, B1 => 
                           REGISTERS_14_31_port, B2 => n1664, ZN => n1570);
   U2017 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n1710, B1 => 
                           REGISTERS_10_31_port, B2 => n1698, ZN => n1569);
   U2018 : NAND4_X1 port map( A1 => n1572, A2 => n1571, A3 => n1570, A4 => 
                           n1569, ZN => n1573);
   U2019 : AOI22_X1 port map( A1 => n1724, A2 => n1575, B1 => n1720, B2 => 
                           n1573, ZN => n1577);
   U2020 : OAI221_X1 port map( B1 => n1581, B2 => n1732, C1 => n1579, C2 => 
                           n1730, A => n1577, ZN => N259);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CWBU is

   port( CLOCK : in std_logic;  ALU_OP : in std_logic_vector (0 to 4);  PSW : 
         in std_logic_vector (6 downto 0);  COND_SEL : out std_logic_vector (1 
         downto 0);  CWB_SEL : in std_logic_vector (1 downto 0);  CWB_MUW_SEL :
         out std_logic_vector (1 downto 0));

end CWBU;

architecture SYN_BEHAVIORAL of CWBU is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal ALUPIPE_4_port, ALUPIPE_2_port, ALUPIPE_1_port, ALUPIPE_0_port, n1, 
      n3, n4, n5, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n2, n6, n7, n8, n9, n10, n_1562, n_1563 : std_logic;

begin
   
   ALUPIPE_reg_0_inst : DFF_X1 port map( D => ALU_OP(4), CK => CLOCK, Q => 
                           ALUPIPE_0_port, QN => n5);
   U24 : NAND3_X1 port map( A1 => n10, A2 => n2, A3 => n11, ZN => 
                           CWB_MUW_SEL(1));
   U25 : NAND3_X1 port map( A1 => n5, A2 => n4, A3 => PSW(0), ZN => n23);
   ALUPIPE_reg_3_inst : DFF_X1 port map( D => ALU_OP(1), CK => CLOCK, Q => 
                           n_1562, QN => n3);
   ALUPIPE_reg_1_inst : DFF_X1 port map( D => ALU_OP(3), CK => CLOCK, Q => 
                           ALUPIPE_1_port, QN => n4);
   ALUPIPE_reg_4_inst : DFF_X1 port map( D => ALU_OP(0), CK => CLOCK, Q => 
                           ALUPIPE_4_port, QN => n1);
   ALUPIPE_reg_2_inst : DFF_X1 port map( D => ALU_OP(2), CK => CLOCK, Q => 
                           ALUPIPE_2_port, QN => n_1563);
   U3 : INV_X1 port map( A => n14, ZN => n2);
   U4 : INV_X1 port map( A => CWB_SEL(1), ZN => n10);
   U5 : AOI221_X1 port map( B1 => PSW(1), B2 => n17, C1 => PSW(3), C2 => n13, A
                           => n22, ZN => n21);
   U6 : OAI21_X1 port map( B1 => n19, B2 => n8, A => n23, ZN => n22);
   U7 : INV_X1 port map( A => PSW(2), ZN => n8);
   U8 : AOI221_X1 port map( B1 => n17, B2 => n9, C1 => n13, C2 => n7, A => n18,
                           ZN => n16);
   U9 : INV_X1 port map( A => PSW(1), ZN => n9);
   U10 : INV_X1 port map( A => PSW(3), ZN => n7);
   U11 : OAI21_X1 port map( B1 => PSW(2), B2 => n19, A => n20, ZN => n18);
   U12 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n13);
   U13 : NOR3_X1 port map( A1 => ALUPIPE_2_port, A2 => ALUPIPE_4_port, A3 => n3
                           , ZN => n14);
   U14 : NAND4_X1 port map( A1 => ALUPIPE_2_port, A2 => n13, A3 => n3, A4 => n1
                           , ZN => n11);
   U15 : NOR2_X1 port map( A1 => n4, A2 => ALUPIPE_0_port, ZN => n17);
   U16 : AND2_X1 port map( A1 => CWB_SEL(0), A2 => n12, ZN => CWB_MUW_SEL(0));
   U17 : OAI211_X1 port map( C1 => n13, C2 => n14, A => n1, B => n15, ZN => n12
                           );
   U18 : XNOR2_X1 port map( A => n3, B => ALUPIPE_2_port, ZN => n15);
   U19 : OAI22_X1 port map( A1 => n21, A2 => n2, B1 => n11, B2 => n6, ZN => 
                           COND_SEL(0));
   U20 : OAI22_X1 port map( A1 => n16, A2 => n2, B1 => PSW(5), B2 => n11, ZN =>
                           COND_SEL(1));
   U21 : NAND2_X1 port map( A1 => ALUPIPE_0_port, A2 => n4, ZN => n19);
   U22 : OR3_X1 port map( A1 => ALUPIPE_1_port, A2 => PSW(0), A3 => 
                           ALUPIPE_0_port, ZN => n20);
   U23 : INV_X1 port map( A => PSW(5), ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 is

   port( clock, rst : in std_logic;  address : in std_logic_vector (31 downto 
         0);  d_in, w_en : in std_logic;  d_out : out std_logic);

end BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0;

architecture SYN_Behavioral of BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal BHT_0_1_port, BHT_0_0_port, BHT_1_1_port, BHT_1_0_port, BHT_2_1_port,
      BHT_2_0_port, BHT_3_1_port, BHT_3_0_port, BHT_4_1_port, BHT_4_0_port, 
      BHT_5_1_port, BHT_5_0_port, BHT_6_1_port, BHT_6_0_port, BHT_7_1_port, 
      BHT_7_0_port, n24, n31, n32, n33, n34, n37, n38, n39, n40, n42, n43, n45,
      n46, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, n62, n63, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      net36148, net36149, net36152, net46252, net46412, net60801, net60817, 
      net60838, net60842, net60854, n7, net36143, net60865, net60864, net60816,
      net36151, net36145, n66, n12, net60822, net36144, n4, n3, n2, n11, 
      N56_port, N55_port, net36154, n47, n41, n36, n1, n5, n6, n8, n9, n10, n13
      , n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, 
      n29, n30, n35, n44, n48, n58, n61, n64, n65, n67, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570,
      n_1571, n_1572 : std_logic;

begin
   d_out <= net60842;
   
   BHT_reg_7_0_inst : DFFR_X1 port map( D => n68, CK => n128, RN => n127, Q => 
                           BHT_7_0_port, QN => n24);
   U80 : NAND3_X1 port map( A1 => d_in, A2 => BHT_7_0_port, A3 => net60842, ZN 
                           => n32);
   U81 : NAND3_X1 port map( A1 => net36149, A2 => n13, A3 => d_in, ZN => n39);
   BHT_reg_5_0_inst : DFFR_X1 port map( D => n71, CK => n128, RN => n127, Q => 
                           BHT_5_0_port, QN => n122);
   BHT_reg_1_0_inst : DFFR_X1 port map( D => n79, CK => n128, RN => n127, Q => 
                           BHT_1_0_port, QN => n125);
   BHT_reg_0_0_inst : DFFR_X1 port map( D => n81, CK => n128, RN => n127, Q => 
                           BHT_0_0_port, QN => n123);
   BHT_reg_3_0_inst : DFFR_X1 port map( D => n75, CK => n128, RN => n127, Q => 
                           BHT_3_0_port, QN => n58);
   BHT_reg_3_1_inst : DFFR_X1 port map( D => n76, CK => n128, RN => n127, Q => 
                           BHT_3_1_port, QN => n_1564);
   BHT_reg_2_0_inst : DFFR_X1 port map( D => n77, CK => n128, RN => n127, Q => 
                           BHT_2_0_port, QN => n_1565);
   BHT_reg_2_1_inst : DFFR_X1 port map( D => n78, CK => n128, RN => n127, Q => 
                           BHT_2_1_port, QN => n_1566);
   BHT_reg_6_0_inst : DFFR_X1 port map( D => n69, CK => n128, RN => n127, Q => 
                           BHT_6_0_port, QN => n_1567);
   BHT_reg_5_1_inst : DFFR_X1 port map( D => n72, CK => n128, RN => n127, Q => 
                           BHT_5_1_port, QN => n_1568);
   BHT_reg_1_1_inst : DFFR_X1 port map( D => n80, CK => n128, RN => n127, Q => 
                           BHT_1_1_port, QN => n_1569);
   BHT_reg_4_1_inst : DFFR_X1 port map( D => n74, CK => n128, RN => n127, Q => 
                           BHT_4_1_port, QN => n_1570);
   BHT_reg_7_1_inst : DFFR_X1 port map( D => n85, CK => n128, RN => n127, Q => 
                           BHT_7_1_port, QN => n113);
   BHT_reg_6_1_inst : DFFR_X1 port map( D => n70, CK => n128, RN => n127, Q => 
                           BHT_6_1_port, QN => n_1571);
   BHT_reg_4_0_inst : DFFR_X1 port map( D => n73, CK => n128, RN => n127, Q => 
                           BHT_4_0_port, QN => n121);
   BHT_reg_0_1_inst : DFFR_X2 port map( D => n82, CK => n128, RN => n127, Q => 
                           BHT_0_1_port, QN => n_1572);
   U3 : AND3_X1 port map( A1 => n23, A2 => address(2), A3 => net36148, ZN => n1
                           );
   U4 : AND2_X1 port map( A1 => n84, A2 => address(2), ZN => n5);
   U5 : OR2_X1 port map( A1 => n106, A2 => n107, ZN => n6);
   U6 : OR2_X1 port map( A1 => n106, A2 => n107, ZN => n35);
   U7 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n8);
   U8 : OR2_X1 port map( A1 => n36, A2 => n117, ZN => n9);
   U9 : OR2_X1 port map( A1 => n36, A2 => n117, ZN => n116);
   U10 : OR2_X1 port map( A1 => n14, A2 => net36143, ZN => n108);
   U11 : INV_X1 port map( A => net60816, ZN => n10);
   U12 : CLKBUF_X1 port map( A => n94, Z => net60864);
   U13 : XNOR2_X1 port map( A => net60801, B => net36151, ZN => n13);
   U14 : BUF_X1 port map( A => address(1), Z => n14);
   U15 : AND2_X1 port map( A1 => n14, A2 => net60817, ZN => net60854);
   U16 : CLKBUF_X1 port map( A => n41, Z => n15);
   U17 : AND2_X1 port map( A1 => BHT_6_0_port, A2 => n84, ZN => n16);
   U18 : AND2_X1 port map( A1 => BHT_7_0_port, A2 => net60854, ZN => n17);
   U19 : NOR3_X1 port map( A1 => n16, A2 => n17, A3 => n44, ZN => n100);
   U20 : AND2_X1 port map( A1 => net36143, A2 => BHT_4_1_port, ZN => n18);
   U21 : OR2_X1 port map( A1 => n37, A2 => n19, ZN => n85);
   U22 : NAND2_X1 port map( A1 => n20, A2 => n114, ZN => n19);
   U23 : OR2_X1 port map( A1 => n112, A2 => n113, ZN => n20);
   U24 : AND2_X1 port map( A1 => BHT_6_0_port, A2 => n46, ZN => n21);
   U25 : AND2_X1 port map( A1 => BHT_7_0_port, A2 => net60854, ZN => n22);
   U26 : NOR3_X1 port map( A1 => n21, A2 => n22, A3 => net36145, ZN => n12);
   U27 : XNOR2_X1 port map( A => net36154, B => n40, ZN => n27);
   U28 : INV_X1 port map( A => n10, ZN => n23);
   U29 : NAND2_X1 port map( A1 => n30, A2 => n35, ZN => n25);
   U30 : XNOR2_X1 port map( A => net36154, B => n13, ZN => n26);
   U31 : AND3_X1 port map( A1 => n28, A2 => n29, A3 => n2, ZN => n3);
   U32 : NAND2_X1 port map( A1 => BHT_2_1_port, A2 => n46, ZN => n28);
   U33 : NAND2_X1 port map( A1 => net60822, A2 => n126, ZN => n29);
   U34 : NAND2_X1 port map( A1 => n30, A2 => n6, ZN => n99);
   U35 : OR2_X1 port map( A1 => n41, A2 => n104, ZN => n30);
   U36 : OAI22_X1 port map( A1 => n121, A2 => n124, B1 => n108, B2 => n122, ZN 
                           => n44);
   U37 : INV_X1 port map( A => address(1), ZN => n48);
   U38 : INV_X1 port map( A => n14, ZN => net36148);
   U39 : BUF_X2 port map( A => address(0), Z => net60817);
   U40 : OR2_X1 port map( A1 => n64, A2 => net60816, ZN => n61);
   U41 : OR2_X1 port map( A1 => n48, A2 => n58, ZN => n64);
   U42 : NOR2_X1 port map( A1 => net36144, A2 => n65, ZN => n11);
   U43 : NAND2_X1 port map( A1 => n67, A2 => n61, ZN => n65);
   U44 : NAND2_X1 port map( A1 => BHT_2_0_port, A2 => n83, ZN => n67);
   U45 : NOR2_X1 port map( A1 => net60817, A2 => n48, ZN => n83);
   U46 : NOR2_X1 port map( A1 => n48, A2 => net60817, ZN => n84);
   U47 : AND2_X1 port map( A1 => n120, A2 => net36143, ZN => n7);
   U48 : INV_X1 port map( A => net60838, ZN => n86);
   U49 : INV_X1 port map( A => n90, ZN => n87);
   U50 : NOR2_X1 port map( A1 => n86, A2 => n87, ZN => n88);
   U51 : NAND2_X1 port map( A1 => n25, A2 => n88, ZN => n89);
   U52 : INV_X1 port map( A => address(2), ZN => n90);
   U53 : NOR2_X1 port map( A1 => n86, A2 => n90, ZN => n91);
   U54 : NAND2_X1 port map( A1 => n99, A2 => n91, ZN => n92);
   U55 : NOR2_X1 port map( A1 => n87, A2 => net60822, ZN => n93);
   U56 : NAND2_X1 port map( A1 => n47, A2 => n95, ZN => n94);
   U57 : AND2_X1 port map( A1 => n23, A2 => n93, ZN => n95);
   U58 : INV_X1 port map( A => n84, ZN => n96);
   U59 : NAND2_X1 port map( A1 => n25, A2 => n98, ZN => n97);
   U60 : NOR2_X1 port map( A1 => n96, A2 => n87, ZN => n98);
   U61 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => n101);
   U62 : NAND2_X1 port map( A1 => n51, A2 => BHT_5_1_port, ZN => n103);
   U63 : NAND2_X1 port map( A1 => n48, A2 => n18, ZN => n102);
   U64 : OR2_X1 port map( A1 => d_in, A2 => n105, ZN => n104);
   U65 : INV_X1 port map( A => w_en, ZN => n105);
   U66 : AND2_X1 port map( A1 => N55_port, A2 => n118, ZN => n106);
   U67 : OR2_X1 port map( A1 => n105, A2 => net36154, ZN => n107);
   U68 : CLKBUF_X1 port map( A => n36, Z => net46252);
   U69 : AND2_X1 port map( A1 => n10, A2 => n90, ZN => n109);
   U70 : NAND2_X1 port map( A1 => n115, A2 => n9, ZN => n110);
   U71 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n55);
   U72 : AND2_X1 port map( A1 => n109, A2 => net60822, ZN => n111);
   U73 : BUF_X2 port map( A => net60865, Z => net46412);
   U74 : INV_X1 port map( A => net46252, ZN => n112);
   U75 : OR2_X1 port map( A1 => n113, A2 => net36149, ZN => n114);
   U76 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => n47);
   U77 : OR2_X1 port map( A1 => n41, A2 => n104, ZN => n115);
   U78 : NAND2_X1 port map( A1 => w_en, A2 => d_in, ZN => n117);
   U79 : OAI22_X1 port map( A1 => n100, A2 => n90, B1 => n11, B2 => address(2),
                           ZN => n118);
   U82 : INV_X1 port map( A => net60865, ZN => n119);
   U83 : AND2_X1 port map( A1 => n120, A2 => address(0), ZN => n51);
   U84 : INV_X1 port map( A => address(1), ZN => n120);
   U85 : OAI22_X1 port map( A1 => n124, A2 => n123, B1 => n108, B2 => n125, ZN 
                           => net36144);
   U86 : OAI22_X1 port map( A1 => n121, A2 => n124, B1 => n108, B2 => n122, ZN 
                           => net36145);
   U87 : INV_X1 port map( A => n7, ZN => n124);
   U88 : MUX2_X1 port map( A => n119, B => BHT_0_0_port, S => n94, Z => n81);
   U89 : NAND2_X1 port map( A1 => n99, A2 => n5, ZN => n42);
   U90 : NAND2_X1 port map( A1 => n47, A2 => n1, ZN => n52);
   U91 : INV_X1 port map( A => d_in, ZN => net36154);
   U92 : AOI21_X1 port map( B1 => net36152, B2 => net36154, A => n34, ZN => n33
                           );
   U93 : NAND4_X1 port map( A1 => w_en, A2 => address(2), A3 => net60822, A4 =>
                           n10, ZN => n34);
   U94 : AND2_X1 port map( A1 => N55_port, A2 => n118, ZN => n36);
   U95 : NOR2_X1 port map( A1 => N55_port, A2 => N56_port, ZN => n41);
   U96 : AOI22_X1 port map( A1 => net36149, A2 => net46252, B1 => n15, B2 => 
                           BHT_7_1_port, ZN => n38);
   U97 : BUF_X1 port map( A => N55_port, Z => net60801);
   U98 : INV_X1 port map( A => N56_port, ZN => net36151);
   U99 : OAI22_X1 port map( A1 => n4, A2 => n90, B1 => n3, B2 => address(2), ZN
                           => N55_port);
   U100 : AOI22_X1 port map( A1 => BHT_0_1_port, A2 => n7, B1 => BHT_1_1_port, 
                           B2 => n51, ZN => n2);
   U101 : AND2_X1 port map( A1 => BHT_3_1_port, A2 => net60817, ZN => n126);
   U102 : INV_X1 port map( A => net36148, ZN => net60822);
   U103 : AOI221_X1 port map( B1 => BHT_6_1_port, B2 => n84, C1 => BHT_7_1_port
                           , C2 => net60854, A => n101, ZN => n4);
   U104 : OAI22_X1 port map( A1 => n12, A2 => n90, B1 => n11, B2 => address(2),
                           ZN => N56_port);
   U105 : INV_X1 port map( A => net60817, ZN => net60816);
   U106 : OAI21_X1 port map( B1 => net60864, B2 => n26, A => n66, ZN => n82);
   U107 : INV_X1 port map( A => net36151, ZN => net60865);
   U108 : XNOR2_X1 port map( A => net60801, B => net36151, ZN => n40);
   U109 : OAI21_X1 port map( B1 => n33, B2 => BHT_7_0_port, A => n119, ZN => 
                           n31);
   U110 : NAND2_X1 port map( A1 => n94, A2 => BHT_0_1_port, ZN => n66);
   U111 : INV_X1 port map( A => address(0), ZN => net36143);
   U112 : NAND2_X1 port map( A1 => n89, A2 => BHT_1_0_port, ZN => n62);
   U113 : NAND2_X1 port map( A1 => n97, A2 => BHT_2_0_port, ZN => n59);
   U114 : NAND2_X1 port map( A1 => BHT_3_0_port, A2 => n55, ZN => n56);
   U115 : INV_X1 port map( A => net36152, ZN => net60842);
   U116 : CLKBUF_X1 port map( A => n51, Z => net60838);
   U117 : INV_X1 port map( A => rst, ZN => n127);
   U118 : INV_X1 port map( A => n34, ZN => net36149);
   U119 : NOR2_X1 port map( A1 => net36148, A2 => net60817, ZN => n46);
   U120 : OAI21_X1 port map( B1 => n27, B2 => n89, A => n63, ZN => n80);
   U121 : NAND2_X1 port map( A1 => n89, A2 => BHT_1_1_port, ZN => n63);
   U122 : OAI21_X1 port map( B1 => n27, B2 => n92, A => n50, ZN => n72);
   U123 : NAND2_X1 port map( A1 => n92, A2 => BHT_5_1_port, ZN => n50);
   U124 : NAND2_X1 port map( A1 => n92, A2 => BHT_5_0_port, ZN => n49);
   U125 : OAI21_X1 port map( B1 => n38, B2 => d_in, A => n39, ZN => n37);
   U126 : OAI21_X1 port map( B1 => n42, B2 => n26, A => n45, ZN => n70);
   U127 : NAND2_X1 port map( A1 => n42, A2 => BHT_6_0_port, ZN => n43);
   U128 : OAI211_X1 port map( C1 => net36149, C2 => n24, A => n31, B => n32, ZN
                           => n68);
   U129 : INV_X1 port map( A => clock, ZN => n128);
   U130 : OAI21_X1 port map( B1 => n27, B2 => n8, A => n57, ZN => n76);
   U131 : NAND2_X1 port map( A1 => BHT_3_1_port, A2 => n55, ZN => n57);
   U132 : NAND2_X1 port map( A1 => n42, A2 => BHT_6_1_port, ZN => n45);
   U133 : OAI21_X1 port map( B1 => n26, B2 => n97, A => n60, ZN => n78);
   U134 : NAND2_X1 port map( A1 => n97, A2 => BHT_2_1_port, ZN => n60);
   U135 : INV_X1 port map( A => net60801, ZN => net36152);
   U136 : NAND2_X1 port map( A1 => n52, A2 => BHT_4_0_port, ZN => n53);
   U137 : NAND2_X1 port map( A1 => n52, A2 => BHT_4_1_port, ZN => n54);
   U138 : OAI21_X1 port map( B1 => n27, B2 => n52, A => n54, ZN => n74);
   U139 : OAI21_X1 port map( B1 => net46412, B2 => n42, A => n43, ZN => n69);
   U140 : OAI21_X1 port map( B1 => net46412, B2 => n92, A => n49, ZN => n71);
   U141 : OAI21_X1 port map( B1 => net46412, B2 => n52, A => n53, ZN => n73);
   U142 : OAI21_X1 port map( B1 => net46412, B2 => n8, A => n56, ZN => n75);
   U143 : OAI21_X1 port map( B1 => net46412, B2 => n97, A => n59, ZN => n77);
   U144 : OAI21_X1 port map( B1 => net46412, B2 => n89, A => n62, ZN => n79);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HDU_IR_SIZE32 is

   port( clk, rst : in std_logic;  IR : in std_logic_vector (31 downto 0);  
         STALL_CODE : out std_logic_vector (1 downto 0);  IF_STALL, ID_STALL, 
         EX_STALL, MEM_STALL, WB_STALL : out std_logic);

end HDU_IR_SIZE32;

architecture SYN_behavioural of HDU_IR_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal STALL_CODE_1_port, IF_STALL_port, EX_STALL_port, cnt_mul_31_port, 
      cnt_mul_30_port, cnt_mul_29_port, cnt_mul_28_port, cnt_mul_27_port, 
      cnt_mul_26_port, cnt_mul_25_port, cnt_mul_24_port, cnt_mul_23_port, 
      cnt_mul_22_port, cnt_mul_21_port, cnt_mul_20_port, cnt_mul_19_port, 
      cnt_mul_18_port, cnt_mul_17_port, cnt_mul_16_port, cnt_mul_15_port, 
      cnt_mul_14_port, cnt_mul_13_port, cnt_mul_12_port, cnt_mul_11_port, 
      cnt_mul_10_port, cnt_mul_9_port, cnt_mul_8_port, cnt_mul_7_port, 
      cnt_mul_6_port, cnt_mul_5_port, cnt_mul_4_port, cnt_mul_3_port, 
      cnt_mul_2_port, cnt_mul_1_port, cnt_mul_0_port, N154, N155, N156, N157, 
      N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, 
      N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, 
      N182, N183, N184, N187, n98, n99, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n149, 
      n150, n151, n152, n153, n154_port, n155_port, n156_port, n157_port, 
      n158_port, n159_port, n169_port, n170_port, n171_port, n172_port, 
      n173_port, n174_port, n175_port, n176_port, n177_port, n178_port, 
      n179_port, n180_port, n181_port, n182_port, n183_port, n184_port, n185, 
      n186, n187_port, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n100, n130, STALL_CODE_0_port, n_1578, n_1579, n_1580, n_1581, 
      n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589 : 
      std_logic;

begin
   STALL_CODE <= ( STALL_CODE_1_port, STALL_CODE_0_port );
   IF_STALL <= IF_STALL_port;
   ID_STALL <= IF_STALL_port;
   EX_STALL <= EX_STALL_port;
   MEM_STALL <= EX_STALL_port;
   WB_STALL <= EX_STALL_port;
   
   cnt_mul_reg_0_inst : DFF_X1 port map( D => n202, CK => clk, Q => 
                           cnt_mul_0_port, QN => n98);
   IR_EX_reg_31_inst : DFFR_X1 port map( D => n159_port, CK => clk, RN => n15, 
                           Q => n130, QN => n_1578);
   IR_EX_reg_30_inst : DFFR_X1 port map( D => n158_port, CK => clk, RN => n15, 
                           Q => n95, QN => n_1579);
   IR_EX_reg_29_inst : DFFR_X1 port map( D => n157_port, CK => clk, RN => n15, 
                           Q => n96, QN => n_1580);
   IR_EX_reg_28_inst : DFFR_X1 port map( D => n156_port, CK => clk, RN => n15, 
                           Q => n100, QN => n_1581);
   IR_EX_reg_27_inst : DFFR_X1 port map( D => n155_port, CK => clk, RN => n15, 
                           Q => n97, QN => n_1582);
   IR_EX_reg_26_inst : DFFR_X1 port map( D => n154_port, CK => clk, RN => n15, 
                           Q => n94, QN => n1);
   IR_EX_reg_20_inst : DFFR_X1 port map( D => n153, CK => clk, RN => n15, Q => 
                           n93, QN => n_1583);
   IR_EX_reg_19_inst : DFFR_X1 port map( D => n152, CK => clk, RN => n15, Q => 
                           n92, QN => n_1584);
   IR_EX_reg_18_inst : DFFR_X1 port map( D => n151, CK => clk, RN => n15, Q => 
                           n91, QN => n_1585);
   IR_EX_reg_17_inst : DFFR_X1 port map( D => n150, CK => clk, RN => n15, Q => 
                           n90, QN => n_1586);
   IR_EX_reg_16_inst : DFFR_X1 port map( D => n149, CK => clk, RN => n15, Q => 
                           n89, QN => n_1587);
   cnt_mul_reg_1_inst : DFF_X1 port map( D => n200, CK => clk, Q => 
                           cnt_mul_1_port, QN => n_1588);
   r100 : HDU_IR_SIZE32_DW01_dec_0_DW01_dec_1 port map( A(31) => 
                           cnt_mul_31_port, A(30) => cnt_mul_30_port, A(29) => 
                           cnt_mul_29_port, A(28) => cnt_mul_28_port, A(27) => 
                           cnt_mul_27_port, A(26) => cnt_mul_26_port, A(25) => 
                           cnt_mul_25_port, A(24) => cnt_mul_24_port, A(23) => 
                           cnt_mul_23_port, A(22) => cnt_mul_22_port, A(21) => 
                           cnt_mul_21_port, A(20) => cnt_mul_20_port, A(19) => 
                           cnt_mul_19_port, A(18) => cnt_mul_18_port, A(17) => 
                           cnt_mul_17_port, A(16) => cnt_mul_16_port, A(15) => 
                           cnt_mul_15_port, A(14) => cnt_mul_14_port, A(13) => 
                           cnt_mul_13_port, A(12) => cnt_mul_12_port, A(11) => 
                           cnt_mul_11_port, A(10) => cnt_mul_10_port, A(9) => 
                           cnt_mul_9_port, A(8) => cnt_mul_8_port, A(7) => 
                           cnt_mul_7_port, A(6) => cnt_mul_6_port, A(5) => 
                           cnt_mul_5_port, A(4) => cnt_mul_4_port, A(3) => 
                           cnt_mul_3_port, A(2) => cnt_mul_2_port, A(1) => 
                           cnt_mul_1_port, A(0) => cnt_mul_0_port, SUM(31) => 
                           N184, SUM(30) => N183, SUM(29) => N182, SUM(28) => 
                           N181, SUM(27) => N180, SUM(26) => N179, SUM(25) => 
                           N178, SUM(24) => N177, SUM(23) => N176, SUM(22) => 
                           N175, SUM(21) => N174, SUM(20) => N173, SUM(19) => 
                           N172, SUM(18) => N171, SUM(17) => N170, SUM(16) => 
                           N169, SUM(15) => N168, SUM(14) => N167, SUM(13) => 
                           N166, SUM(12) => N165, SUM(11) => N164, SUM(10) => 
                           N163, SUM(9) => N162, SUM(8) => N161, SUM(7) => N160
                           , SUM(6) => N159, SUM(5) => N158, SUM(4) => N157, 
                           SUM(3) => N156, SUM(2) => N155, SUM(1) => N154, 
                           SUM(0) => n_1589);
   cnt_mul_reg_5_inst : DFF_X1 port map( D => n194, CK => clk, Q => 
                           cnt_mul_5_port, QN => n104);
   cnt_mul_reg_6_inst : DFF_X1 port map( D => n193, CK => clk, Q => 
                           cnt_mul_6_port, QN => n105);
   cnt_mul_reg_4_inst : DFF_X1 port map( D => n195, CK => clk, Q => 
                           cnt_mul_4_port, QN => n103);
   cnt_mul_reg_3_inst : DFF_X1 port map( D => n196, CK => clk, Q => 
                           cnt_mul_3_port, QN => n102);
   cnt_mul_reg_2_inst : DFF_X1 port map( D => n197, CK => clk, Q => 
                           cnt_mul_2_port, QN => n101);
   cnt_mul_reg_26_inst : DFF_X1 port map( D => n173_port, CK => clk, Q => 
                           cnt_mul_26_port, QN => n125);
   cnt_mul_reg_25_inst : DFF_X1 port map( D => n174_port, CK => clk, Q => 
                           cnt_mul_25_port, QN => n124);
   cnt_mul_reg_24_inst : DFF_X1 port map( D => n175_port, CK => clk, Q => 
                           cnt_mul_24_port, QN => n123);
   cnt_mul_reg_23_inst : DFF_X1 port map( D => n176_port, CK => clk, Q => 
                           cnt_mul_23_port, QN => n122);
   cnt_mul_reg_22_inst : DFF_X1 port map( D => n177_port, CK => clk, Q => 
                           cnt_mul_22_port, QN => n121);
   cnt_mul_reg_21_inst : DFF_X1 port map( D => n178_port, CK => clk, Q => 
                           cnt_mul_21_port, QN => n120);
   cnt_mul_reg_20_inst : DFF_X1 port map( D => n179_port, CK => clk, Q => 
                           cnt_mul_20_port, QN => n119);
   cnt_mul_reg_19_inst : DFF_X1 port map( D => n180_port, CK => clk, Q => 
                           cnt_mul_19_port, QN => n118);
   cnt_mul_reg_18_inst : DFF_X1 port map( D => n181_port, CK => clk, Q => 
                           cnt_mul_18_port, QN => n117);
   cnt_mul_reg_17_inst : DFF_X1 port map( D => n182_port, CK => clk, Q => 
                           cnt_mul_17_port, QN => n116);
   cnt_mul_reg_16_inst : DFF_X1 port map( D => n183_port, CK => clk, Q => 
                           cnt_mul_16_port, QN => n115);
   cnt_mul_reg_15_inst : DFF_X1 port map( D => n184_port, CK => clk, Q => 
                           cnt_mul_15_port, QN => n114);
   cnt_mul_reg_14_inst : DFF_X1 port map( D => n185, CK => clk, Q => 
                           cnt_mul_14_port, QN => n113);
   cnt_mul_reg_13_inst : DFF_X1 port map( D => n186, CK => clk, Q => 
                           cnt_mul_13_port, QN => n112);
   cnt_mul_reg_12_inst : DFF_X1 port map( D => n187_port, CK => clk, Q => 
                           cnt_mul_12_port, QN => n111);
   cnt_mul_reg_11_inst : DFF_X1 port map( D => n188, CK => clk, Q => 
                           cnt_mul_11_port, QN => n110);
   cnt_mul_reg_10_inst : DFF_X1 port map( D => n189, CK => clk, Q => 
                           cnt_mul_10_port, QN => n109);
   cnt_mul_reg_9_inst : DFF_X1 port map( D => n190, CK => clk, Q => 
                           cnt_mul_9_port, QN => n108);
   cnt_mul_reg_30_inst : DFF_X1 port map( D => n169_port, CK => clk, Q => 
                           cnt_mul_30_port, QN => n129);
   cnt_mul_reg_29_inst : DFF_X1 port map( D => n170_port, CK => clk, Q => 
                           cnt_mul_29_port, QN => n128);
   cnt_mul_reg_28_inst : DFF_X1 port map( D => n171_port, CK => clk, Q => 
                           cnt_mul_28_port, QN => n127);
   cnt_mul_reg_27_inst : DFF_X1 port map( D => n172_port, CK => clk, Q => 
                           cnt_mul_27_port, QN => n126);
   cnt_mul_reg_31_inst : DFF_X1 port map( D => n198, CK => clk, Q => 
                           cnt_mul_31_port, QN => n99);
   cnt_mul_reg_8_inst : DFF_X1 port map( D => n191, CK => clk, Q => 
                           cnt_mul_8_port, QN => n107);
   cnt_mul_reg_7_inst : DFF_X1 port map( D => n192, CK => clk, Q => 
                           cnt_mul_7_port, QN => n106);
   STALL_MUL_reg : DFF_X1 port map( D => n201, CK => clk, Q => EX_STALL_port, 
                           QN => n199);
   U3 : INV_X1 port map( A => n107, ZN => n2);
   U4 : BUF_X1 port map( A => n7, Z => n10);
   U5 : NAND3_X1 port map( A1 => n3, A2 => n4, A3 => n5, ZN => n30);
   U6 : NOR3_X1 port map( A1 => IR(10), A2 => IR(5), A3 => IR(4), ZN => n3);
   U7 : NOR4_X1 port map( A1 => IR(9), A2 => IR(8), A3 => IR(7), A4 => IR(6), 
                           ZN => n4);
   U8 : NOR4_X1 port map( A1 => n63, A2 => n64, A3 => IR(0), A4 => n65, ZN => 
                           n5);
   U9 : AND2_X1 port map( A1 => n199, A2 => n30, ZN => n7);
   U10 : INV_X1 port map( A => n106, ZN => n6);
   U11 : BUF_X1 port map( A => n32, Z => n12);
   U12 : BUF_X1 port map( A => n32, Z => n13);
   U13 : BUF_X1 port map( A => n32, Z => n14);
   U14 : INV_X1 port map( A => rst, ZN => n15);
   U15 : INV_X1 port map( A => n10, ZN => n8);
   U16 : INV_X1 port map( A => n10, ZN => n9);
   U17 : BUF_X1 port map( A => n7, Z => n11);
   U18 : NOR3_X1 port map( A1 => cnt_mul_0_port, A2 => cnt_mul_11_port, A3 => 
                           cnt_mul_10_port, ZN => n19);
   U19 : NOR4_X1 port map( A1 => cnt_mul_15_port, A2 => cnt_mul_14_port, A3 => 
                           cnt_mul_13_port, A4 => cnt_mul_12_port, ZN => n18);
   U20 : NOR4_X1 port map( A1 => cnt_mul_19_port, A2 => cnt_mul_18_port, A3 => 
                           cnt_mul_17_port, A4 => cnt_mul_16_port, ZN => n17);
   U21 : NOR4_X1 port map( A1 => cnt_mul_22_port, A2 => cnt_mul_21_port, A3 => 
                           cnt_mul_20_port, A4 => cnt_mul_1_port, ZN => n16);
   U22 : AND4_X1 port map( A1 => n19, A2 => n18, A3 => n17, A4 => n16, ZN => 
                           n25);
   U23 : NOR4_X1 port map( A1 => cnt_mul_26_port, A2 => cnt_mul_25_port, A3 => 
                           cnt_mul_24_port, A4 => cnt_mul_23_port, ZN => n23);
   U24 : NOR4_X1 port map( A1 => cnt_mul_2_port, A2 => cnt_mul_29_port, A3 => 
                           cnt_mul_28_port, A4 => cnt_mul_27_port, ZN => n22);
   U25 : NOR4_X1 port map( A1 => cnt_mul_5_port, A2 => cnt_mul_4_port, A3 => 
                           cnt_mul_3_port, A4 => cnt_mul_30_port, ZN => n21);
   U26 : NOR4_X1 port map( A1 => cnt_mul_9_port, A2 => n2, A3 => n6, A4 => 
                           cnt_mul_6_port, ZN => n20);
   U27 : AND4_X1 port map( A1 => n23, A2 => n22, A3 => n21, A4 => n20, ZN => 
                           n24);
   U28 : AOI21_X1 port map( B1 => n25, B2 => n24, A => cnt_mul_31_port, ZN => 
                           N187);
   U29 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n202);
   U30 : XOR2_X1 port map( A => n8, B => n98, Z => n26);
   U31 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => n200);
   U32 : INV_X1 port map( A => n29, ZN => n28);
   U33 : MUX2_X1 port map( A => N154, B => cnt_mul_1_port, S => n11, Z => n29);
   U34 : NAND3_X1 port map( A1 => n30, A2 => n31, A3 => n8, ZN => n27);
   U35 : OAI22_X1 port map( A1 => n14, A2 => n33, B1 => n99, B2 => n8, ZN => 
                           n198);
   U36 : INV_X1 port map( A => N184, ZN => n33);
   U37 : OAI22_X1 port map( A1 => n14, A2 => n34, B1 => n101, B2 => n8, ZN => 
                           n197);
   U38 : INV_X1 port map( A => N155, ZN => n34);
   U39 : OAI22_X1 port map( A1 => n14, A2 => n35, B1 => n102, B2 => n8, ZN => 
                           n196);
   U40 : INV_X1 port map( A => N156, ZN => n35);
   U41 : OAI22_X1 port map( A1 => n14, A2 => n36, B1 => n103, B2 => n8, ZN => 
                           n195);
   U42 : INV_X1 port map( A => N157, ZN => n36);
   U43 : OAI22_X1 port map( A1 => n14, A2 => n37, B1 => n104, B2 => n8, ZN => 
                           n194);
   U44 : INV_X1 port map( A => N158, ZN => n37);
   U45 : OAI22_X1 port map( A1 => n14, A2 => n38, B1 => n105, B2 => n8, ZN => 
                           n193);
   U46 : INV_X1 port map( A => N159, ZN => n38);
   U47 : OAI22_X1 port map( A1 => n14, A2 => n39, B1 => n106, B2 => n8, ZN => 
                           n192);
   U48 : INV_X1 port map( A => N160, ZN => n39);
   U49 : OAI22_X1 port map( A1 => n14, A2 => n40, B1 => n107, B2 => n8, ZN => 
                           n191);
   U50 : INV_X1 port map( A => N161, ZN => n40);
   U51 : OAI22_X1 port map( A1 => n13, A2 => n41, B1 => n108, B2 => n8, ZN => 
                           n190);
   U52 : INV_X1 port map( A => N162, ZN => n41);
   U53 : OAI22_X1 port map( A1 => n13, A2 => n42, B1 => n109, B2 => n8, ZN => 
                           n189);
   U54 : INV_X1 port map( A => N163, ZN => n42);
   U55 : OAI22_X1 port map( A1 => n13, A2 => n43, B1 => n110, B2 => n8, ZN => 
                           n188);
   U56 : INV_X1 port map( A => N164, ZN => n43);
   U57 : OAI22_X1 port map( A1 => n13, A2 => n44, B1 => n111, B2 => n8, ZN => 
                           n187_port);
   U58 : INV_X1 port map( A => N165, ZN => n44);
   U59 : OAI22_X1 port map( A1 => n13, A2 => n45, B1 => n112, B2 => n9, ZN => 
                           n186);
   U60 : INV_X1 port map( A => N166, ZN => n45);
   U61 : OAI22_X1 port map( A1 => n13, A2 => n46, B1 => n113, B2 => n9, ZN => 
                           n185);
   U62 : INV_X1 port map( A => N167, ZN => n46);
   U63 : OAI22_X1 port map( A1 => n13, A2 => n47, B1 => n114, B2 => n9, ZN => 
                           n184_port);
   U64 : INV_X1 port map( A => N168, ZN => n47);
   U65 : OAI22_X1 port map( A1 => n13, A2 => n48, B1 => n115, B2 => n9, ZN => 
                           n183_port);
   U66 : INV_X1 port map( A => N169, ZN => n48);
   U67 : OAI22_X1 port map( A1 => n13, A2 => n49, B1 => n116, B2 => n9, ZN => 
                           n182_port);
   U68 : INV_X1 port map( A => N170, ZN => n49);
   U69 : OAI22_X1 port map( A1 => n13, A2 => n50, B1 => n117, B2 => n9, ZN => 
                           n181_port);
   U70 : INV_X1 port map( A => N171, ZN => n50);
   U71 : OAI22_X1 port map( A1 => n13, A2 => n51, B1 => n118, B2 => n9, ZN => 
                           n180_port);
   U72 : INV_X1 port map( A => N172, ZN => n51);
   U73 : OAI22_X1 port map( A1 => n12, A2 => n52, B1 => n119, B2 => n9, ZN => 
                           n179_port);
   U74 : INV_X1 port map( A => N173, ZN => n52);
   U75 : OAI22_X1 port map( A1 => n12, A2 => n53, B1 => n120, B2 => n9, ZN => 
                           n178_port);
   U76 : INV_X1 port map( A => N174, ZN => n53);
   U77 : OAI22_X1 port map( A1 => n12, A2 => n54, B1 => n121, B2 => n9, ZN => 
                           n177_port);
   U78 : INV_X1 port map( A => N175, ZN => n54);
   U79 : OAI22_X1 port map( A1 => n12, A2 => n55, B1 => n122, B2 => n9, ZN => 
                           n176_port);
   U80 : INV_X1 port map( A => N176, ZN => n55);
   U81 : OAI22_X1 port map( A1 => n12, A2 => n56, B1 => n123, B2 => n9, ZN => 
                           n175_port);
   U82 : INV_X1 port map( A => N177, ZN => n56);
   U83 : OAI22_X1 port map( A1 => n12, A2 => n57, B1 => n124, B2 => n9, ZN => 
                           n174_port);
   U84 : INV_X1 port map( A => N178, ZN => n57);
   U85 : OAI22_X1 port map( A1 => n12, A2 => n58, B1 => n125, B2 => n9, ZN => 
                           n173_port);
   U86 : INV_X1 port map( A => N179, ZN => n58);
   U87 : OAI22_X1 port map( A1 => n12, A2 => n59, B1 => n126, B2 => n9, ZN => 
                           n172_port);
   U88 : INV_X1 port map( A => N180, ZN => n59);
   U89 : OAI22_X1 port map( A1 => n12, A2 => n60, B1 => n127, B2 => n9, ZN => 
                           n171_port);
   U90 : INV_X1 port map( A => N181, ZN => n60);
   U91 : OAI22_X1 port map( A1 => n12, A2 => n61, B1 => n128, B2 => n9, ZN => 
                           n170_port);
   U92 : INV_X1 port map( A => N182, ZN => n61);
   U93 : OAI22_X1 port map( A1 => n12, A2 => n62, B1 => n129, B2 => n9, ZN => 
                           n169_port);
   U94 : INV_X1 port map( A => N183, ZN => n62);
   U95 : INV_X1 port map( A => n201, ZN => n32);
   U96 : AOI21_X1 port map( B1 => n30, B2 => n31, A => n11, ZN => n201);
   U97 : INV_X1 port map( A => N187, ZN => n31);
   U98 : INV_X1 port map( A => IR(26), ZN => n64);
   U99 : NAND3_X1 port map( A1 => IR(2), A2 => IR(1), A3 => IR(3), ZN => n63);
   U100 : MUX2_X1 port map( A => n130, B => IR(31), S => n199, Z => n159_port);
   U101 : MUX2_X1 port map( A => n95, B => IR(30), S => n199, Z => n158_port);
   U102 : MUX2_X1 port map( A => n96, B => IR(29), S => n199, Z => n157_port);
   U103 : MUX2_X1 port map( A => n100, B => IR(28), S => n199, Z => n156_port);
   U104 : MUX2_X1 port map( A => n97, B => IR(27), S => n199, Z => n155_port);
   U105 : MUX2_X1 port map( A => n94, B => IR(26), S => n199, Z => n154_port);
   U106 : MUX2_X1 port map( A => n93, B => IR(20), S => n199, Z => n153);
   U107 : MUX2_X1 port map( A => n92, B => IR(19), S => n199, Z => n152);
   U108 : MUX2_X1 port map( A => n91, B => IR(18), S => n199, Z => n151);
   U109 : MUX2_X1 port map( A => n90, B => IR(17), S => n199, Z => n150);
   U110 : MUX2_X1 port map( A => n89, B => IR(16), S => n199, Z => n149);
   U111 : NOR2_X1 port map( A1 => n199, A2 => STALL_CODE_0_port, ZN => 
                           STALL_CODE_1_port);
   U112 : INV_X1 port map( A => n66, ZN => STALL_CODE_0_port);
   U113 : NAND2_X1 port map( A1 => n199, A2 => n66, ZN => IF_STALL_port);
   U114 : NAND3_X1 port map( A1 => n130, A2 => n67, A3 => n68, ZN => n66);
   U115 : AOI211_X1 port map( C1 => n69, C2 => n70, A => n95, B => n96, ZN => 
                           n68);
   U116 : NAND4_X1 port map( A1 => n71, A2 => n72, A3 => n73, A4 => n74, ZN => 
                           n70);
   U117 : NOR3_X1 port map( A1 => n75, A2 => n76, A3 => n77, ZN => n74);
   U118 : XOR2_X1 port map( A => n89, B => IR(21), Z => n77);
   U119 : XOR2_X1 port map( A => n90, B => IR(22), Z => n76);
   U120 : XOR2_X1 port map( A => n93, B => IR(25), Z => n75);
   U121 : XNOR2_X1 port map( A => n91, B => IR(23), ZN => n73);
   U122 : OR4_X1 port map( A1 => n78, A2 => n79, A3 => IR(29), A4 => IR(31), ZN
                           => n72);
   U123 : MUX2_X1 port map( A => n80, B => IR(28), S => IR(27), Z => n78);
   U124 : AOI21_X1 port map( B1 => IR(28), B2 => IR(26), A => n81, ZN => n80);
   U125 : INV_X1 port map( A => IR(30), ZN => n81);
   U126 : XNOR2_X1 port map( A => n92, B => IR(24), ZN => n71);
   U127 : NAND4_X1 port map( A1 => n82, A2 => n79, A3 => n83, A4 => n84, ZN => 
                           n69);
   U128 : NOR3_X1 port map( A1 => n85, A2 => n86, A3 => n87, ZN => n84);
   U129 : XOR2_X1 port map( A => n89, B => IR(16), Z => n87);
   U130 : XOR2_X1 port map( A => n90, B => IR(17), Z => n86);
   U131 : XOR2_X1 port map( A => n93, B => IR(20), Z => n85);
   U132 : XNOR2_X1 port map( A => IR(18), B => n91, ZN => n83);
   U133 : NOR2_X1 port map( A1 => n65, A2 => IR(26), ZN => n79);
   U134 : OR4_X1 port map( A1 => IR(30), A2 => IR(31), A3 => IR(29), A4 => n88,
                           ZN => n65);
   U135 : OR2_X1 port map( A1 => IR(28), A2 => IR(27), ZN => n88);
   U136 : XNOR2_X1 port map( A => IR(19), B => n92, ZN => n82);
   U137 : OAI21_X1 port map( B1 => n100, B2 => n1, A => n97, ZN => n67);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWDU_IR_SIZE32 is

   port( CLOCK, RESET, EN : in std_logic;  IR : in std_logic_vector (31 downto 
         0);  FWD_A, FWD_B : out std_logic_vector (1 downto 0);  FWD_B2 : out 
         std_logic;  ZDU_SEL : out std_logic_vector (1 downto 0));

end FWDU_IR_SIZE32;

architecture SYN_BEHAVIORAL of FWDU_IR_SIZE32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal FWD_B2_port, ZDU_SEL_1_port, ZDU_SEL_0_port, n106, n107, n108, n109, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n175, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n174, n176, n177, n_1590, 
      n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, 
      n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, 
      n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, 
      n_1618, n_1619, n_1620, n_1621, n_1622 : std_logic;

begin
   FWD_B2 <= FWD_B2_port;
   ZDU_SEL <= ( ZDU_SEL_1_port, ZDU_SEL_0_port );
   
   IR_EX_reg_31_inst : DFFR_X1 port map( D => n175, CK => CLOCK, RN => n7, Q =>
                           n121, QN => n2);
   IR_EX_reg_30_inst : DFFR_X1 port map( D => n173, CK => CLOCK, RN => n7, Q =>
                           n123, QN => n_1590);
   IR_EX_reg_29_inst : DFFR_X1 port map( D => n172, CK => CLOCK, RN => n7, Q =>
                           n122, QN => n_1591);
   IR_EX_reg_28_inst : DFFR_X1 port map( D => n171, CK => CLOCK, RN => n7, Q =>
                           n110, QN => n_1592);
   IR_EX_reg_27_inst : DFFR_X1 port map( D => n170, CK => CLOCK, RN => n7, Q =>
                           n105, QN => n_1593);
   IR_EX_reg_26_inst : DFFR_X1 port map( D => n169, CK => CLOCK, RN => n7, Q =>
                           n104, QN => n_1594);
   IR_EX_reg_20_inst : DFFR_X1 port map( D => n168, CK => CLOCK, RN => n7, Q =>
                           n120, QN => n_1595);
   IR_EX_reg_19_inst : DFFR_X1 port map( D => n167, CK => CLOCK, RN => n7, Q =>
                           n118, QN => n_1596);
   IR_EX_reg_18_inst : DFFR_X1 port map( D => n166, CK => CLOCK, RN => n7, Q =>
                           n116, QN => n_1597);
   IR_EX_reg_17_inst : DFFR_X1 port map( D => n165, CK => CLOCK, RN => n7, Q =>
                           n114, QN => n_1598);
   IR_EX_reg_16_inst : DFFR_X1 port map( D => n164, CK => CLOCK, RN => n7, Q =>
                           n112, QN => n_1599);
   IR_EX_reg_15_inst : DFFR_X1 port map( D => n163, CK => CLOCK, RN => n8, Q =>
                           n119, QN => n_1600);
   IR_EX_reg_14_inst : DFFR_X1 port map( D => n162, CK => CLOCK, RN => n8, Q =>
                           n117, QN => n_1601);
   IR_EX_reg_13_inst : DFFR_X1 port map( D => n161, CK => CLOCK, RN => n8, Q =>
                           n115, QN => n_1602);
   IR_EX_reg_12_inst : DFFR_X1 port map( D => n160, CK => CLOCK, RN => n8, Q =>
                           n113, QN => n_1603);
   IR_EX_reg_11_inst : DFFR_X1 port map( D => n159, CK => CLOCK, RN => n8, Q =>
                           n111, QN => n_1604);
   IR_MEM_reg_31_inst : DFFR_X1 port map( D => n158, CK => CLOCK, RN => n8, Q 
                           => n134, QN => n_1605);
   IR_MEM_reg_30_inst : DFFR_X1 port map( D => n157, CK => CLOCK, RN => n8, Q 
                           => n176, QN => n1);
   IR_MEM_reg_29_inst : DFFR_X1 port map( D => n156, CK => CLOCK, RN => n8, Q 
                           => n177, QN => n_1606);
   IR_MEM_reg_28_inst : DFFR_X1 port map( D => n155, CK => CLOCK, RN => n8, Q 
                           => n135, QN => n_1607);
   IR_MEM_reg_27_inst : DFFR_X1 port map( D => n154, CK => CLOCK, RN => n8, Q 
                           => n174, QN => n_1608);
   IR_MEM_reg_20_inst : DFFR_X1 port map( D => n153, CK => CLOCK, RN => n8, Q 
                           => n133, QN => n_1609);
   IR_MEM_reg_19_inst : DFFR_X1 port map( D => n152, CK => CLOCK, RN => n9, Q 
                           => n131, QN => n_1610);
   IR_MEM_reg_18_inst : DFFR_X1 port map( D => n151, CK => CLOCK, RN => n9, Q 
                           => n129, QN => n_1611);
   IR_MEM_reg_17_inst : DFFR_X1 port map( D => n150, CK => CLOCK, RN => n9, Q 
                           => n127, QN => n_1612);
   IR_MEM_reg_16_inst : DFFR_X1 port map( D => n149, CK => CLOCK, RN => n9, Q 
                           => n125, QN => n_1613);
   IR_MEM_reg_15_inst : DFFR_X1 port map( D => n148, CK => CLOCK, RN => n9, Q 
                           => n132, QN => n_1614);
   IR_MEM_reg_14_inst : DFFR_X1 port map( D => n147, CK => CLOCK, RN => n9, Q 
                           => n130, QN => n_1615);
   IR_MEM_reg_13_inst : DFFR_X1 port map( D => n146, CK => CLOCK, RN => n9, Q 
                           => n128, QN => n_1616);
   IR_MEM_reg_12_inst : DFFR_X1 port map( D => n145, CK => CLOCK, RN => n9, Q 
                           => n126, QN => n_1617);
   IR_MEM_reg_11_inst : DFFR_X1 port map( D => n144, CK => CLOCK, RN => n9, Q 
                           => n124, QN => n_1618);
   FWD_B2_tmp2_reg : DFF_X1 port map( D => n143, CK => CLOCK, Q => n103, QN => 
                           n_1619);
   FWD_B2_reg : DFF_X1 port map( D => n142, CK => CLOCK, Q => FWD_B2_port, QN 
                           => n_1620);
   FWD_A_reg_1_inst : DFF_X1 port map( D => n141, CK => CLOCK, Q => FWD_A(1), 
                           QN => n109);
   FWD_A_reg_0_inst : DFF_X1 port map( D => n140, CK => CLOCK, Q => FWD_A(0), 
                           QN => n108);
   FWD_B_reg_1_inst : DFF_X1 port map( D => n139, CK => CLOCK, Q => FWD_B(1), 
                           QN => n107);
   FWD_B_reg_0_inst : DFF_X1 port map( D => n138, CK => CLOCK, Q => FWD_B(0), 
                           QN => n106);
   ZDU_SEL_reg_1_inst : DFF_X1 port map( D => n137, CK => CLOCK, Q => 
                           ZDU_SEL_1_port, QN => n_1621);
   ZDU_SEL_reg_0_inst : DFF_X1 port map( D => n136, CK => CLOCK, Q => 
                           ZDU_SEL_0_port, QN => n_1622);
   U2 : NOR4_X2 port map( A1 => n135, A2 => n134, A3 => n174, A4 => n102, ZN =>
                           n83);
   U3 : NOR4_X2 port map( A1 => n110, A2 => n105, A3 => n121, A4 => n97, ZN => 
                           n92);
   U4 : BUF_X1 port map( A => EN, Z => n6);
   U5 : BUF_X1 port map( A => n10, Z => n8);
   U6 : BUF_X1 port map( A => n10, Z => n7);
   U7 : BUF_X1 port map( A => n10, Z => n9);
   U8 : BUF_X1 port map( A => n6, Z => n5);
   U9 : BUF_X1 port map( A => n6, Z => n4);
   U10 : BUF_X1 port map( A => n6, Z => n3);
   U11 : INV_X1 port map( A => RESET, ZN => n10);
   U12 : MUX2_X1 port map( A => n121, B => IR(31), S => n3, Z => n175);
   U13 : MUX2_X1 port map( A => n123, B => IR(30), S => n3, Z => n173);
   U14 : MUX2_X1 port map( A => n122, B => IR(29), S => n3, Z => n172);
   U15 : MUX2_X1 port map( A => n110, B => IR(28), S => n3, Z => n171);
   U16 : MUX2_X1 port map( A => n105, B => IR(27), S => n3, Z => n170);
   U17 : MUX2_X1 port map( A => n104, B => IR(26), S => n3, Z => n169);
   U18 : MUX2_X1 port map( A => n120, B => IR(20), S => n3, Z => n168);
   U19 : MUX2_X1 port map( A => n118, B => IR(19), S => n3, Z => n167);
   U20 : MUX2_X1 port map( A => n116, B => IR(18), S => n3, Z => n166);
   U21 : MUX2_X1 port map( A => n114, B => IR(17), S => n3, Z => n165);
   U22 : MUX2_X1 port map( A => n112, B => IR(16), S => n3, Z => n164);
   U23 : MUX2_X1 port map( A => n119, B => IR(15), S => n4, Z => n163);
   U24 : MUX2_X1 port map( A => n117, B => IR(14), S => n4, Z => n162);
   U25 : MUX2_X1 port map( A => n115, B => IR(13), S => n4, Z => n161);
   U26 : MUX2_X1 port map( A => n113, B => IR(12), S => n4, Z => n160);
   U27 : MUX2_X1 port map( A => n111, B => IR(11), S => n4, Z => n159);
   U28 : MUX2_X1 port map( A => n134, B => n121, S => n4, Z => n158);
   U29 : MUX2_X1 port map( A => n176, B => n123, S => n4, Z => n157);
   U30 : MUX2_X1 port map( A => n177, B => n122, S => n4, Z => n156);
   U31 : MUX2_X1 port map( A => n135, B => n110, S => n4, Z => n155);
   U32 : MUX2_X1 port map( A => n174, B => n105, S => n4, Z => n154);
   U33 : MUX2_X1 port map( A => n133, B => n120, S => n4, Z => n153);
   U34 : MUX2_X1 port map( A => n131, B => n118, S => n5, Z => n152);
   U35 : MUX2_X1 port map( A => n129, B => n116, S => n5, Z => n151);
   U36 : MUX2_X1 port map( A => n127, B => n114, S => n5, Z => n150);
   U37 : MUX2_X1 port map( A => n125, B => n112, S => n5, Z => n149);
   U38 : MUX2_X1 port map( A => n132, B => n119, S => n5, Z => n148);
   U39 : MUX2_X1 port map( A => n130, B => n117, S => n5, Z => n147);
   U40 : MUX2_X1 port map( A => n128, B => n115, S => n5, Z => n146);
   U41 : MUX2_X1 port map( A => n126, B => n113, S => n5, Z => n145);
   U42 : MUX2_X1 port map( A => n124, B => n111, S => n5, Z => n144);
   U43 : MUX2_X1 port map( A => n103, B => n11, S => n12, Z => n143);
   U44 : AND4_X1 port map( A1 => n13, A2 => n14, A3 => IR(31), A4 => IR(29), ZN
                           => n11);
   U45 : AND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n13);
   U46 : INV_X1 port map( A => IR(30), ZN => n18);
   U47 : OR4_X1 port map( A1 => IR(19), A2 => IR(20), A3 => IR(18), A4 => n19, 
                           ZN => n16);
   U48 : OR2_X1 port map( A1 => IR(17), A2 => IR(16), ZN => n19);
   U49 : NAND2_X1 port map( A1 => IR(27), A2 => n20, ZN => n15);
   U50 : MUX2_X1 port map( A => FWD_B2_port, B => n103, S => n12, Z => n142);
   U51 : OAI21_X1 port map( B1 => n109, B2 => n12, A => n21, ZN => n141);
   U52 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n21);
   U53 : NOR2_X1 port map( A1 => n26, A2 => n27, ZN => n25);
   U54 : OAI22_X1 port map( A1 => n108, A2 => n12, B1 => n27, B2 => n28, ZN => 
                           n140);
   U55 : OR2_X1 port map( A1 => n23, A2 => n22, ZN => n28);
   U56 : OAI21_X1 port map( B1 => n107, B2 => n12, A => n29, ZN => n139);
   U57 : NAND4_X1 port map( A1 => n24, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           n29);
   U58 : NOR2_X1 port map( A1 => n27, A2 => n33, ZN => n32);
   U59 : INV_X1 port map( A => n34, ZN => n33);
   U60 : OAI21_X1 port map( B1 => n35, B2 => n36, A => n37, ZN => n31);
   U61 : NAND4_X1 port map( A1 => n38, A2 => n39, A3 => n40, A4 => n41, ZN => 
                           n37);
   U62 : NOR2_X1 port map( A1 => n42, A2 => n43, ZN => n41);
   U63 : XOR2_X1 port map( A => IR(18), B => n44, Z => n43);
   U64 : XOR2_X1 port map( A => IR(20), B => n45, Z => n42);
   U65 : XNOR2_X1 port map( A => n46, B => IR(16), ZN => n40);
   U66 : XNOR2_X1 port map( A => n47, B => IR(17), ZN => n39);
   U67 : XNOR2_X1 port map( A => n48, B => IR(19), ZN => n38);
   U68 : INV_X1 port map( A => n49, ZN => n36);
   U69 : INV_X1 port map( A => n50, ZN => n24);
   U70 : OAI22_X1 port map( A1 => n106, A2 => n12, B1 => n27, B2 => n30, ZN => 
                           n138);
   U71 : NAND3_X1 port map( A1 => n34, A2 => n14, A3 => n51, ZN => n30);
   U72 : AOI21_X1 port map( B1 => n49, B2 => n20, A => n22, ZN => n51);
   U73 : INV_X1 port map( A => IR(26), ZN => n20);
   U74 : NOR4_X1 port map( A1 => n52, A2 => n2, A3 => n123, A4 => n122, ZN => 
                           n49);
   U75 : MUX2_X1 port map( A => n105, B => n110, S => n104, Z => n52);
   U76 : INV_X1 port map( A => n35, ZN => n14);
   U77 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           n35);
   U78 : NOR2_X1 port map( A1 => n57, A2 => n58, ZN => n56);
   U79 : XOR2_X1 port map( A => IR(17), B => n59, Z => n58);
   U80 : XOR2_X1 port map( A => IR(20), B => n60, Z => n57);
   U81 : XNOR2_X1 port map( A => n61, B => IR(19), ZN => n55);
   U82 : XNOR2_X1 port map( A => n62, B => IR(16), ZN => n54);
   U83 : XNOR2_X1 port map( A => n63, B => IR(18), ZN => n53);
   U84 : NOR2_X1 port map( A1 => n64, A2 => IR(28), ZN => n34);
   U85 : OAI221_X1 port map( B1 => n22, B2 => n65, C1 => n50, C2 => n66, A => 
                           n12, ZN => n27);
   U86 : NOR3_X1 port map( A1 => n177, A2 => n134, A3 => n67, ZN => n50);
   U87 : MUX2_X1 port map( A => n68, B => n135, S => n174, Z => n67);
   U88 : NAND2_X1 port map( A1 => n1, A2 => n135, ZN => n68);
   U89 : NOR3_X1 port map( A1 => n122, A2 => n121, A3 => n69, ZN => n22);
   U90 : INV_X1 port map( A => n70, ZN => n69);
   U91 : MUX2_X1 port map( A => n105, B => n71, S => n110, Z => n70);
   U92 : NOR2_X1 port map( A1 => n105, A2 => n123, ZN => n71);
   U93 : MUX2_X1 port map( A => ZDU_SEL_1_port, B => n72, S => n12, Z => n137);
   U94 : NOR4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           n72);
   U95 : INV_X1 port map( A => n23, ZN => n75);
   U96 : OR3_X1 port map( A1 => n26, A2 => n17, A3 => n64, ZN => n73);
   U97 : INV_X1 port map( A => IR(28), ZN => n17);
   U98 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           n26);
   U99 : NOR2_X1 port map( A1 => n81, A2 => n82, ZN => n80);
   U100 : XOR2_X1 port map( A => IR(24), B => n48, Z => n82);
   U101 : XOR2_X1 port map( A => IR(25), B => n45, Z => n81);
   U102 : XNOR2_X1 port map( A => n46, B => IR(21), ZN => n79);
   U103 : MUX2_X1 port map( A => n125, B => n124, S => n83, Z => n46);
   U104 : XNOR2_X1 port map( A => n47, B => IR(22), ZN => n78);
   U105 : MUX2_X1 port map( A => n127, B => n126, S => n83, Z => n47);
   U106 : XNOR2_X1 port map( A => n44, B => IR(23), ZN => n77);
   U107 : MUX2_X1 port map( A => n129, B => n128, S => n83, Z => n44);
   U108 : MUX2_X1 port map( A => ZDU_SEL_0_port, B => n84, S => n12, Z => n136)
                           ;
   U109 : AND2_X1 port map( A1 => n5, A2 => n9, ZN => n12);
   U110 : NOR3_X1 port map( A1 => n85, A2 => n23, A3 => n64, ZN => n84);
   U111 : OR4_X1 port map( A1 => IR(27), A2 => IR(29), A3 => IR(30), A4 => 
                           IR(31), ZN => n64);
   U112 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           n23);
   U113 : NOR2_X1 port map( A1 => n90, A2 => n91, ZN => n89);
   U114 : XOR2_X1 port map( A => IR(23), B => n63, Z => n91);
   U115 : MUX2_X1 port map( A => n116, B => n115, S => n92, Z => n63);
   U116 : XOR2_X1 port map( A => IR(22), B => n59, Z => n90);
   U117 : MUX2_X1 port map( A => n114, B => n113, S => n92, Z => n59);
   U118 : XNOR2_X1 port map( A => n62, B => IR(21), ZN => n88);
   U119 : MUX2_X1 port map( A => n112, B => n111, S => n92, Z => n62);
   U120 : XNOR2_X1 port map( A => n60, B => IR(25), ZN => n87);
   U121 : XNOR2_X1 port map( A => n61, B => IR(24), ZN => n86);
   U122 : NAND3_X1 port map( A1 => n66, A2 => n65, A3 => IR(28), ZN => n85);
   U123 : INV_X1 port map( A => n76, ZN => n65);
   U124 : NOR3_X1 port map( A1 => n60, A2 => n61, A3 => n93, ZN => n76);
   U125 : INV_X1 port map( A => n94, ZN => n93);
   U126 : MUX2_X1 port map( A => n95, B => n96, S => n92, Z => n94);
   U127 : NOR3_X1 port map( A1 => n115, A2 => n111, A3 => n113, ZN => n96);
   U128 : NOR3_X1 port map( A1 => n116, A2 => n112, A3 => n114, ZN => n95);
   U129 : MUX2_X1 port map( A => n118, B => n117, S => n92, Z => n61);
   U130 : MUX2_X1 port map( A => n120, B => n119, S => n92, Z => n60);
   U131 : OR2_X1 port map( A1 => n122, A2 => n123, ZN => n97);
   U132 : INV_X1 port map( A => n74, ZN => n66);
   U133 : NOR3_X1 port map( A1 => n48, A2 => n45, A3 => n98, ZN => n74);
   U134 : INV_X1 port map( A => n99, ZN => n98);
   U135 : MUX2_X1 port map( A => n100, B => n101, S => n83, Z => n99);
   U136 : NOR3_X1 port map( A1 => n128, A2 => n124, A3 => n126, ZN => n101);
   U137 : NOR3_X1 port map( A1 => n129, A2 => n125, A3 => n127, ZN => n100);
   U138 : MUX2_X1 port map( A => n133, B => n132, S => n83, Z => n45);
   U139 : MUX2_X1 port map( A => n131, B => n130, S => n83, Z => n48);
   U140 : OR2_X1 port map( A1 => n176, A2 => n177, ZN => n102);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( CLOCK : in std_logic;  AluOpcode : in std_logic_vector (0 to 4);  A, B
         : in std_logic_vector (31 downto 0);  Cin : in std_logic;  ALU_out : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic;  COND : out
         std_logic_vector (5 downto 0));

end ALU_NBIT32;

architecture SYN_BEHAVIORAL of ALU_NBIT32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX4to1_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUL
      port( CLOCK : in std_logic;  A, B : in std_logic_vector (15 downto 0);  Y
            : out std_logic_vector (31 downto 0));
   end component;
   
   component CMP_NBIT32
      port( SUM : in std_logic_vector (31 downto 0);  Cout : in std_logic;  
            A_L_B, A_LE_B, A_G_B, A_GE_B, A_E_B, A_NE_B : out std_logic);
   end component;
   
   component LOGIC_NBIT32_N_SELECTOR4
      port( S : in std_logic_vector (3 downto 0);  A, B : in std_logic_vector 
            (31 downto 0);  O : out std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER
      port( data_in : in std_logic_vector (31 downto 0);  R : in 
            std_logic_vector (4 downto 0);  conf : in std_logic_vector (1 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  ADD_SUB, Cin : in 
            std_logic;  S : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   component AND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal Cout_port, cin_internal, en_adder, A_adder_31_port, A_adder_30_port, 
      A_adder_29_port, A_adder_28_port, A_adder_27_port, A_adder_26_port, 
      A_adder_25_port, A_adder_24_port, A_adder_23_port, A_adder_22_port, 
      A_adder_21_port, A_adder_20_port, A_adder_19_port, A_adder_18_port, 
      A_adder_17_port, A_adder_16_port, A_adder_15_port, A_adder_14_port, 
      A_adder_13_port, A_adder_12_port, A_adder_11_port, A_adder_10_port, 
      A_adder_9_port, A_adder_8_port, A_adder_7_port, A_adder_6_port, 
      A_adder_5_port, A_adder_4_port, A_adder_3_port, A_adder_2_port, 
      A_adder_1_port, A_adder_0_port, B_adder_31_port, B_adder_30_port, 
      B_adder_29_port, B_adder_28_port, B_adder_27_port, B_adder_26_port, 
      B_adder_25_port, B_adder_24_port, B_adder_23_port, B_adder_22_port, 
      B_adder_21_port, B_adder_20_port, B_adder_19_port, B_adder_18_port, 
      B_adder_17_port, B_adder_16_port, B_adder_15_port, B_adder_14_port, 
      B_adder_13_port, B_adder_12_port, B_adder_11_port, B_adder_10_port, 
      B_adder_9_port, B_adder_8_port, B_adder_7_port, B_adder_6_port, 
      B_adder_5_port, B_adder_4_port, B_adder_3_port, B_adder_2_port, 
      B_adder_1_port, B_adder_0_port, en_logic, A_logic_31_port, 
      A_logic_30_port, A_logic_29_port, A_logic_28_port, A_logic_27_port, 
      A_logic_26_port, A_logic_25_port, A_logic_24_port, A_logic_23_port, 
      A_logic_22_port, A_logic_21_port, A_logic_20_port, A_logic_19_port, 
      A_logic_18_port, A_logic_17_port, A_logic_16_port, A_logic_15_port, 
      A_logic_14_port, A_logic_13_port, A_logic_12_port, A_logic_11_port, 
      A_logic_10_port, A_logic_9_port, A_logic_8_port, A_logic_7_port, 
      A_logic_6_port, A_logic_5_port, A_logic_4_port, A_logic_3_port, 
      A_logic_2_port, A_logic_1_port, A_logic_0_port, B_logic_31_port, 
      B_logic_30_port, B_logic_29_port, B_logic_28_port, B_logic_27_port, 
      B_logic_26_port, B_logic_25_port, B_logic_24_port, B_logic_23_port, 
      B_logic_22_port, B_logic_21_port, B_logic_20_port, B_logic_19_port, 
      B_logic_18_port, B_logic_17_port, B_logic_16_port, B_logic_15_port, 
      B_logic_14_port, B_logic_13_port, B_logic_12_port, B_logic_11_port, 
      B_logic_10_port, B_logic_9_port, B_logic_8_port, B_logic_7_port, 
      B_logic_6_port, B_logic_5_port, B_logic_4_port, B_logic_3_port, 
      B_logic_2_port, B_logic_1_port, B_logic_0_port, en_shifter, 
      A_shifter_31_port, A_shifter_30_port, A_shifter_29_port, 
      A_shifter_28_port, A_shifter_27_port, A_shifter_26_port, 
      A_shifter_25_port, A_shifter_24_port, A_shifter_23_port, 
      A_shifter_22_port, A_shifter_21_port, A_shifter_20_port, 
      A_shifter_19_port, A_shifter_18_port, A_shifter_17_port, 
      A_shifter_16_port, A_shifter_15_port, A_shifter_14_port, 
      A_shifter_13_port, A_shifter_12_port, A_shifter_11_port, 
      A_shifter_10_port, A_shifter_9_port, A_shifter_8_port, A_shifter_7_port, 
      A_shifter_6_port, A_shifter_5_port, A_shifter_4_port, A_shifter_3_port, 
      A_shifter_2_port, A_shifter_1_port, A_shifter_0_port, B_shifter_4_port, 
      B_shifter_3_port, B_shifter_2_port, B_shifter_1_port, B_shifter_0_port, 
      en_cmp, in_cmp_31_port, in_cmp_30_port, in_cmp_29_port, in_cmp_28_port, 
      in_cmp_27_port, in_cmp_26_port, in_cmp_25_port, in_cmp_24_port, 
      in_cmp_23_port, in_cmp_22_port, in_cmp_21_port, in_cmp_20_port, 
      in_cmp_19_port, in_cmp_18_port, in_cmp_17_port, in_cmp_16_port, 
      in_cmp_15_port, in_cmp_14_port, in_cmp_13_port, in_cmp_12_port, 
      in_cmp_11_port, in_cmp_10_port, in_cmp_9_port, in_cmp_8_port, 
      in_cmp_7_port, in_cmp_6_port, in_cmp_5_port, in_cmp_4_port, in_cmp_3_port
      , in_cmp_2_port, in_cmp_1_port, in_cmp_0_port, out_adder_31_port, 
      out_adder_30_port, out_adder_29_port, out_adder_28_port, 
      out_adder_27_port, out_adder_26_port, out_adder_25_port, 
      out_adder_24_port, out_adder_23_port, out_adder_22_port, 
      out_adder_21_port, out_adder_20_port, out_adder_19_port, 
      out_adder_18_port, out_adder_17_port, out_adder_16_port, 
      out_adder_15_port, out_adder_14_port, out_adder_13_port, 
      out_adder_12_port, out_adder_11_port, out_adder_10_port, out_adder_9_port
      , out_adder_8_port, out_adder_7_port, out_adder_6_port, out_adder_5_port,
      out_adder_4_port, out_adder_3_port, out_adder_2_port, out_adder_1_port, 
      out_adder_0_port, A_mul_15_port, A_mul_14_port, A_mul_13_port, 
      A_mul_12_port, A_mul_11_port, A_mul_10_port, A_mul_9_port, A_mul_8_port, 
      A_mul_7_port, A_mul_6_port, A_mul_5_port, A_mul_4_port, A_mul_3_port, 
      A_mul_2_port, A_mul_1_port, A_mul_0_port, B_mul_15_port, B_mul_14_port, 
      B_mul_13_port, B_mul_12_port, B_mul_11_port, B_mul_10_port, B_mul_9_port,
      B_mul_8_port, B_mul_7_port, B_mul_6_port, B_mul_5_port, B_mul_4_port, 
      B_mul_3_port, B_mul_2_port, B_mul_1_port, B_mul_0_port, conf_1_port, 
      conf_0_port, out_shifter_31_port, out_shifter_30_port, 
      out_shifter_29_port, out_shifter_28_port, out_shifter_27_port, 
      out_shifter_26_port, out_shifter_25_port, out_shifter_24_port, 
      out_shifter_23_port, out_shifter_22_port, out_shifter_21_port, 
      out_shifter_20_port, out_shifter_19_port, out_shifter_18_port, 
      out_shifter_17_port, out_shifter_16_port, out_shifter_15_port, 
      out_shifter_14_port, out_shifter_13_port, out_shifter_12_port, 
      out_shifter_11_port, out_shifter_10_port, out_shifter_9_port, 
      out_shifter_8_port, out_shifter_7_port, out_shifter_6_port, 
      out_shifter_5_port, out_shifter_4_port, out_shifter_3_port, 
      out_shifter_2_port, out_shifter_1_port, out_shifter_0_port, 
      logic_sel_3_port, logic_sel_2_port, logic_sel_1_port, logic_sel_0_port, 
      out_logic_31_port, out_logic_30_port, out_logic_29_port, 
      out_logic_28_port, out_logic_27_port, out_logic_26_port, 
      out_logic_25_port, out_logic_24_port, out_logic_23_port, 
      out_logic_22_port, out_logic_21_port, out_logic_20_port, 
      out_logic_19_port, out_logic_18_port, out_logic_17_port, 
      out_logic_16_port, out_logic_15_port, out_logic_14_port, 
      out_logic_13_port, out_logic_12_port, out_logic_11_port, 
      out_logic_10_port, out_logic_9_port, out_logic_8_port, out_logic_7_port, 
      out_logic_6_port, out_logic_5_port, out_logic_4_port, out_logic_3_port, 
      out_logic_2_port, out_logic_1_port, out_logic_0_port, out_mul_31_port, 
      out_mul_30_port, out_mul_29_port, out_mul_28_port, out_mul_27_port, 
      out_mul_26_port, out_mul_25_port, out_mul_24_port, out_mul_23_port, 
      out_mul_22_port, out_mul_21_port, out_mul_20_port, out_mul_19_port, 
      out_mul_18_port, out_mul_17_port, out_mul_16_port, out_mul_15_port, 
      out_mul_14_port, out_mul_13_port, out_mul_12_port, out_mul_11_port, 
      out_mul_10_port, out_mul_9_port, out_mul_8_port, out_mul_7_port, 
      out_mul_6_port, out_mul_5_port, out_mul_4_port, out_mul_3_port, 
      out_mul_2_port, out_mul_1_port, out_mul_0_port, mux_out_1_port, 
      mux_out_0_port, N88, N89, N90, N91, N92, N93, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n1, n2, n3, n4, n5, n6, n7, n8, n9, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62 : std_logic;

begin
   Cout <= Cout_port;
   
   conf_reg_1_inst : DLH_X1 port map( G => N91, D => N93, Q => conf_1_port);
   conf_reg_0_inst : DLH_X1 port map( G => N91, D => N92, Q => conf_0_port);
   logic_sel_reg_3_inst : DLH_X1 port map( G => n50, D => N90, Q => 
                           logic_sel_3_port);
   logic_sel_reg_2_inst : DLH_X1 port map( G => n49, D => N89, Q => 
                           logic_sel_2_port);
   logic_sel_reg_1_inst : DLH_X1 port map( G => n50, D => N89, Q => 
                           logic_sel_1_port);
   logic_sel_reg_0_inst : DLH_X1 port map( G => n49, D => N88, Q => 
                           logic_sel_0_port);
   U37 : NAND3_X1 port map( A1 => n14, A2 => n57, A3 => n15, ZN => n12);
   U38 : XOR2_X1 port map( A => AluOpcode(3), B => AluOpcode(4), Z => n14);
   U39 : NAND3_X1 port map( A1 => n60, A2 => n57, A3 => AluOpcode(1), ZN => n18
                           );
   U40 : XOR2_X1 port map( A => AluOpcode(2), B => n19, Z => n23);
   U41 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n29, ZN => N89);
   U42 : NAND3_X1 port map( A1 => n56, A2 => AluOpcode(4), A3 => AluOpcode(1), 
                           ZN => n29);
   U43 : NAND3_X1 port map( A1 => AluOpcode(2), A2 => n57, A3 => AluOpcode(3), 
                           ZN => n17);
   U44 : NAND3_X1 port map( A1 => n11, A2 => n62, A3 => n15, ZN => n28);
   U45 : NAND3_X1 port map( A1 => AluOpcode(0), A2 => n62, A3 => n15, ZN => n25
                           );
   ADDER_A_i_0 : AND2_0 port map( A => A(0), B => n6, Y => A_adder_0_port);
   ADDER_B_i_0 : AND2_228 port map( A => B(0), B => en_adder, Y => 
                           B_adder_0_port);
   ADDER_A_i_1 : AND2_227 port map( A => A(1), B => n3, Y => A_adder_1_port);
   ADDER_B_i_1 : AND2_226 port map( A => B(1), B => n6, Y => B_adder_1_port);
   ADDER_A_i_2 : AND2_225 port map( A => A(2), B => n4, Y => A_adder_2_port);
   ADDER_B_i_2 : AND2_224 port map( A => B(2), B => n5, Y => B_adder_2_port);
   ADDER_A_i_3 : AND2_223 port map( A => A(3), B => n7, Y => A_adder_3_port);
   ADDER_B_i_3 : AND2_222 port map( A => B(3), B => n6, Y => B_adder_3_port);
   ADDER_A_i_4 : AND2_221 port map( A => A(4), B => n7, Y => A_adder_4_port);
   ADDER_B_i_4 : AND2_220 port map( A => B(4), B => n2, Y => B_adder_4_port);
   ADDER_A_i_5 : AND2_219 port map( A => A(5), B => n3, Y => A_adder_5_port);
   ADDER_B_i_5 : AND2_218 port map( A => B(5), B => n6, Y => B_adder_5_port);
   ADDER_A_i_6 : AND2_217 port map( A => A(6), B => n7, Y => A_adder_6_port);
   ADDER_B_i_6 : AND2_216 port map( A => B(6), B => n4, Y => B_adder_6_port);
   ADDER_A_i_7 : AND2_215 port map( A => A(7), B => n7, Y => A_adder_7_port);
   ADDER_B_i_7 : AND2_214 port map( A => B(7), B => n6, Y => B_adder_7_port);
   ADDER_A_i_8 : AND2_213 port map( A => A(8), B => n4, Y => A_adder_8_port);
   ADDER_B_i_8 : AND2_212 port map( A => B(8), B => n2, Y => B_adder_8_port);
   ADDER_A_i_9 : AND2_211 port map( A => A(9), B => n7, Y => A_adder_9_port);
   ADDER_B_i_9 : AND2_210 port map( A => B(9), B => n3, Y => B_adder_9_port);
   ADDER_A_i_10 : AND2_209 port map( A => A(10), B => n7, Y => A_adder_10_port)
                           ;
   ADDER_B_i_10 : AND2_208 port map( A => B(10), B => n4, Y => B_adder_10_port)
                           ;
   ADDER_A_i_11 : AND2_207 port map( A => A(11), B => n3, Y => A_adder_11_port)
                           ;
   ADDER_B_i_11 : AND2_206 port map( A => B(11), B => n7, Y => B_adder_11_port)
                           ;
   ADDER_A_i_12 : AND2_205 port map( A => A(12), B => n2, Y => A_adder_12_port)
                           ;
   ADDER_B_i_12 : AND2_204 port map( A => B(12), B => n4, Y => B_adder_12_port)
                           ;
   ADDER_A_i_13 : AND2_203 port map( A => A(13), B => n7, Y => A_adder_13_port)
                           ;
   ADDER_B_i_13 : AND2_202 port map( A => B(13), B => n6, Y => B_adder_13_port)
                           ;
   ADDER_A_i_14 : AND2_201 port map( A => A(14), B => n4, Y => A_adder_14_port)
                           ;
   ADDER_B_i_14 : AND2_200 port map( A => B(14), B => n2, Y => B_adder_14_port)
                           ;
   ADDER_A_i_15 : AND2_199 port map( A => A(15), B => n3, Y => A_adder_15_port)
                           ;
   ADDER_B_i_15 : AND2_198 port map( A => B(15), B => n6, Y => B_adder_15_port)
                           ;
   ADDER_A_i_16 : AND2_197 port map( A => A(16), B => n3, Y => A_adder_16_port)
                           ;
   ADDER_B_i_16 : AND2_196 port map( A => B(16), B => n2, Y => B_adder_16_port)
                           ;
   ADDER_A_i_17 : AND2_195 port map( A => A(17), B => n3, Y => A_adder_17_port)
                           ;
   ADDER_B_i_17 : AND2_194 port map( A => B(17), B => n7, Y => B_adder_17_port)
                           ;
   ADDER_A_i_18 : AND2_193 port map( A => A(18), B => n7, Y => A_adder_18_port)
                           ;
   ADDER_B_i_18 : AND2_192 port map( A => B(18), B => n4, Y => B_adder_18_port)
                           ;
   ADDER_A_i_19 : AND2_191 port map( A => A(19), B => n3, Y => A_adder_19_port)
                           ;
   ADDER_B_i_19 : AND2_190 port map( A => B(19), B => n4, Y => B_adder_19_port)
                           ;
   ADDER_A_i_20 : AND2_189 port map( A => A(20), B => n2, Y => A_adder_20_port)
                           ;
   ADDER_B_i_20 : AND2_188 port map( A => B(20), B => n2, Y => B_adder_20_port)
                           ;
   ADDER_A_i_21 : AND2_187 port map( A => A(21), B => n2, Y => A_adder_21_port)
                           ;
   ADDER_B_i_21 : AND2_186 port map( A => B(21), B => n3, Y => B_adder_21_port)
                           ;
   ADDER_A_i_22 : AND2_185 port map( A => A(22), B => n2, Y => A_adder_22_port)
                           ;
   ADDER_B_i_22 : AND2_184 port map( A => B(22), B => n4, Y => B_adder_22_port)
                           ;
   ADDER_A_i_23 : AND2_183 port map( A => A(23), B => n2, Y => A_adder_23_port)
                           ;
   ADDER_B_i_23 : AND2_182 port map( A => B(23), B => n3, Y => B_adder_23_port)
                           ;
   ADDER_A_i_24 : AND2_181 port map( A => A(24), B => n4, Y => A_adder_24_port)
                           ;
   ADDER_B_i_24 : AND2_180 port map( A => B(24), B => n4, Y => B_adder_24_port)
                           ;
   ADDER_A_i_25 : AND2_179 port map( A => A(25), B => n7, Y => A_adder_25_port)
                           ;
   ADDER_B_i_25 : AND2_178 port map( A => B(25), B => n4, Y => B_adder_25_port)
                           ;
   ADDER_A_i_26 : AND2_177 port map( A => A(26), B => n3, Y => A_adder_26_port)
                           ;
   ADDER_B_i_26 : AND2_176 port map( A => B(26), B => n3, Y => B_adder_26_port)
                           ;
   ADDER_A_i_27 : AND2_175 port map( A => A(27), B => n4, Y => A_adder_27_port)
                           ;
   ADDER_B_i_27 : AND2_174 port map( A => B(27), B => n4, Y => B_adder_27_port)
                           ;
   ADDER_A_i_28 : AND2_173 port map( A => A(28), B => n3, Y => A_adder_28_port)
                           ;
   ADDER_B_i_28 : AND2_172 port map( A => B(28), B => n2, Y => B_adder_28_port)
                           ;
   ADDER_A_i_29 : AND2_171 port map( A => A(29), B => n3, Y => A_adder_29_port)
                           ;
   ADDER_B_i_29 : AND2_170 port map( A => B(29), B => n7, Y => B_adder_29_port)
                           ;
   ADDER_A_i_30 : AND2_169 port map( A => A(30), B => n2, Y => A_adder_30_port)
                           ;
   ADDER_B_i_30 : AND2_168 port map( A => B(30), B => n2, Y => B_adder_30_port)
                           ;
   ADDER_A_i_31 : AND2_167 port map( A => A(31), B => n7, Y => A_adder_31_port)
                           ;
   ADDER_B_i_31 : AND2_166 port map( A => B(31), B => n4, Y => B_adder_31_port)
                           ;
   LOGIC_A_i_0 : AND2_165 port map( A => A(0), B => n44, Y => A_logic_0_port);
   LOGIC_B_i_0 : AND2_164 port map( A => B(0), B => n48, Y => B_logic_0_port);
   LOGIC_A_i_1 : AND2_163 port map( A => A(1), B => n49, Y => A_logic_1_port);
   LOGIC_B_i_1 : AND2_162 port map( A => B(1), B => n49, Y => B_logic_1_port);
   LOGIC_A_i_2 : AND2_161 port map( A => A(2), B => n49, Y => A_logic_2_port);
   LOGIC_B_i_2 : AND2_160 port map( A => B(2), B => n49, Y => B_logic_2_port);
   LOGIC_A_i_3 : AND2_159 port map( A => A(3), B => n49, Y => A_logic_3_port);
   LOGIC_B_i_3 : AND2_158 port map( A => B(3), B => n49, Y => B_logic_3_port);
   LOGIC_A_i_4 : AND2_157 port map( A => A(4), B => n49, Y => A_logic_4_port);
   LOGIC_B_i_4 : AND2_156 port map( A => B(4), B => n49, Y => B_logic_4_port);
   LOGIC_A_i_5 : AND2_155 port map( A => A(5), B => n49, Y => A_logic_5_port);
   LOGIC_B_i_5 : AND2_154 port map( A => B(5), B => n48, Y => B_logic_5_port);
   LOGIC_A_i_6 : AND2_153 port map( A => A(6), B => n48, Y => A_logic_6_port);
   LOGIC_B_i_6 : AND2_152 port map( A => B(6), B => n48, Y => B_logic_6_port);
   LOGIC_A_i_7 : AND2_151 port map( A => A(7), B => n48, Y => A_logic_7_port);
   LOGIC_B_i_7 : AND2_150 port map( A => B(7), B => n48, Y => B_logic_7_port);
   LOGIC_A_i_8 : AND2_149 port map( A => A(8), B => n48, Y => A_logic_8_port);
   LOGIC_B_i_8 : AND2_148 port map( A => B(8), B => n48, Y => B_logic_8_port);
   LOGIC_A_i_9 : AND2_147 port map( A => A(9), B => n48, Y => A_logic_9_port);
   LOGIC_B_i_9 : AND2_146 port map( A => B(9), B => n48, Y => B_logic_9_port);
   LOGIC_A_i_10 : AND2_145 port map( A => A(10), B => n48, Y => A_logic_10_port
                           );
   LOGIC_B_i_10 : AND2_144 port map( A => B(10), B => n47, Y => B_logic_10_port
                           );
   LOGIC_A_i_11 : AND2_143 port map( A => A(11), B => n47, Y => A_logic_11_port
                           );
   LOGIC_B_i_11 : AND2_142 port map( A => B(11), B => n47, Y => B_logic_11_port
                           );
   LOGIC_A_i_12 : AND2_141 port map( A => A(12), B => n47, Y => A_logic_12_port
                           );
   LOGIC_B_i_12 : AND2_140 port map( A => B(12), B => n47, Y => B_logic_12_port
                           );
   LOGIC_A_i_13 : AND2_139 port map( A => A(13), B => n47, Y => A_logic_13_port
                           );
   LOGIC_B_i_13 : AND2_138 port map( A => B(13), B => n47, Y => B_logic_13_port
                           );
   LOGIC_A_i_14 : AND2_137 port map( A => A(14), B => n47, Y => A_logic_14_port
                           );
   LOGIC_B_i_14 : AND2_136 port map( A => B(14), B => n47, Y => B_logic_14_port
                           );
   LOGIC_A_i_15 : AND2_135 port map( A => A(15), B => n47, Y => A_logic_15_port
                           );
   LOGIC_B_i_15 : AND2_134 port map( A => B(15), B => n47, Y => B_logic_15_port
                           );
   LOGIC_A_i_16 : AND2_133 port map( A => A(16), B => n46, Y => A_logic_16_port
                           );
   LOGIC_B_i_16 : AND2_132 port map( A => B(16), B => n46, Y => B_logic_16_port
                           );
   LOGIC_A_i_17 : AND2_131 port map( A => A(17), B => n46, Y => A_logic_17_port
                           );
   LOGIC_B_i_17 : AND2_130 port map( A => B(17), B => n46, Y => B_logic_17_port
                           );
   LOGIC_A_i_18 : AND2_129 port map( A => A(18), B => n46, Y => A_logic_18_port
                           );
   LOGIC_B_i_18 : AND2_128 port map( A => B(18), B => n46, Y => B_logic_18_port
                           );
   LOGIC_A_i_19 : AND2_127 port map( A => A(19), B => n46, Y => A_logic_19_port
                           );
   LOGIC_B_i_19 : AND2_126 port map( A => B(19), B => n46, Y => B_logic_19_port
                           );
   LOGIC_A_i_20 : AND2_125 port map( A => A(20), B => n46, Y => A_logic_20_port
                           );
   LOGIC_B_i_20 : AND2_124 port map( A => B(20), B => n46, Y => B_logic_20_port
                           );
   LOGIC_A_i_21 : AND2_123 port map( A => A(21), B => n45, Y => A_logic_21_port
                           );
   LOGIC_B_i_21 : AND2_122 port map( A => B(21), B => n45, Y => B_logic_21_port
                           );
   LOGIC_A_i_22 : AND2_121 port map( A => A(22), B => n45, Y => A_logic_22_port
                           );
   LOGIC_B_i_22 : AND2_120 port map( A => B(22), B => n45, Y => B_logic_22_port
                           );
   LOGIC_A_i_23 : AND2_119 port map( A => A(23), B => n45, Y => A_logic_23_port
                           );
   LOGIC_B_i_23 : AND2_118 port map( A => B(23), B => n45, Y => B_logic_23_port
                           );
   LOGIC_A_i_24 : AND2_117 port map( A => A(24), B => n45, Y => A_logic_24_port
                           );
   LOGIC_B_i_24 : AND2_116 port map( A => B(24), B => n45, Y => B_logic_24_port
                           );
   LOGIC_A_i_25 : AND2_115 port map( A => A(25), B => n45, Y => A_logic_25_port
                           );
   LOGIC_B_i_25 : AND2_114 port map( A => B(25), B => n45, Y => B_logic_25_port
                           );
   LOGIC_A_i_26 : AND2_113 port map( A => A(26), B => n46, Y => A_logic_26_port
                           );
   LOGIC_B_i_26 : AND2_112 port map( A => B(26), B => n45, Y => B_logic_26_port
                           );
   LOGIC_A_i_27 : AND2_111 port map( A => A(27), B => n44, Y => A_logic_27_port
                           );
   LOGIC_B_i_27 : AND2_110 port map( A => B(27), B => n44, Y => B_logic_27_port
                           );
   LOGIC_A_i_28 : AND2_109 port map( A => A(28), B => n44, Y => A_logic_28_port
                           );
   LOGIC_B_i_28 : AND2_108 port map( A => B(28), B => n44, Y => B_logic_28_port
                           );
   LOGIC_A_i_29 : AND2_107 port map( A => A(29), B => n44, Y => A_logic_29_port
                           );
   LOGIC_B_i_29 : AND2_106 port map( A => B(29), B => n44, Y => B_logic_29_port
                           );
   LOGIC_A_i_30 : AND2_105 port map( A => A(30), B => n44, Y => A_logic_30_port
                           );
   LOGIC_B_i_30 : AND2_104 port map( A => B(30), B => n44, Y => B_logic_30_port
                           );
   LOGIC_A_i_31 : AND2_103 port map( A => A(31), B => n44, Y => A_logic_31_port
                           );
   LOGIC_B_i_31 : AND2_102 port map( A => B(31), B => n44, Y => B_logic_31_port
                           );
   SHIFTER_A_i_0 : AND2_101 port map( A => A(0), B => n36, Y => 
                           A_shifter_0_port);
   SHIFTER_A_i_1 : AND2_100 port map( A => A(1), B => n36, Y => 
                           A_shifter_1_port);
   SHIFTER_A_i_2 : AND2_99 port map( A => A(2), B => n36, Y => A_shifter_2_port
                           );
   SHIFTER_A_i_3 : AND2_98 port map( A => A(3), B => n36, Y => A_shifter_3_port
                           );
   SHIFTER_A_i_4 : AND2_97 port map( A => A(4), B => n36, Y => A_shifter_4_port
                           );
   SHIFTER_A_i_5 : AND2_96 port map( A => A(5), B => n36, Y => A_shifter_5_port
                           );
   SHIFTER_A_i_6 : AND2_95 port map( A => A(6), B => n36, Y => A_shifter_6_port
                           );
   SHIFTER_A_i_7 : AND2_94 port map( A => A(7), B => n36, Y => A_shifter_7_port
                           );
   SHIFTER_A_i_8 : AND2_93 port map( A => A(8), B => n36, Y => A_shifter_8_port
                           );
   SHIFTER_A_i_9 : AND2_92 port map( A => A(9), B => n36, Y => A_shifter_9_port
                           );
   SHIFTER_A_i_10 : AND2_91 port map( A => A(10), B => n36, Y => 
                           A_shifter_10_port);
   SHIFTER_A_i_11 : AND2_90 port map( A => A(11), B => n37, Y => 
                           A_shifter_11_port);
   SHIFTER_A_i_12 : AND2_89 port map( A => A(12), B => n37, Y => 
                           A_shifter_12_port);
   SHIFTER_A_i_13 : AND2_88 port map( A => A(13), B => n37, Y => 
                           A_shifter_13_port);
   SHIFTER_A_i_14 : AND2_87 port map( A => A(14), B => n37, Y => 
                           A_shifter_14_port);
   SHIFTER_A_i_15 : AND2_86 port map( A => A(15), B => n37, Y => 
                           A_shifter_15_port);
   SHIFTER_A_i_16 : AND2_85 port map( A => A(16), B => n37, Y => 
                           A_shifter_16_port);
   SHIFTER_A_i_17 : AND2_84 port map( A => A(17), B => n37, Y => 
                           A_shifter_17_port);
   SHIFTER_A_i_18 : AND2_83 port map( A => A(18), B => n37, Y => 
                           A_shifter_18_port);
   SHIFTER_A_i_19 : AND2_82 port map( A => A(19), B => n37, Y => 
                           A_shifter_19_port);
   SHIFTER_A_i_20 : AND2_81 port map( A => A(20), B => n37, Y => 
                           A_shifter_20_port);
   SHIFTER_A_i_21 : AND2_80 port map( A => A(21), B => n37, Y => 
                           A_shifter_21_port);
   SHIFTER_A_i_22 : AND2_79 port map( A => A(22), B => n38, Y => 
                           A_shifter_22_port);
   SHIFTER_A_i_23 : AND2_78 port map( A => A(23), B => n38, Y => 
                           A_shifter_23_port);
   SHIFTER_A_i_24 : AND2_77 port map( A => A(24), B => n38, Y => 
                           A_shifter_24_port);
   SHIFTER_A_i_25 : AND2_76 port map( A => A(25), B => n38, Y => 
                           A_shifter_25_port);
   SHIFTER_A_i_26 : AND2_75 port map( A => A(26), B => n38, Y => 
                           A_shifter_26_port);
   SHIFTER_A_i_27 : AND2_74 port map( A => A(27), B => n38, Y => 
                           A_shifter_27_port);
   SHIFTER_A_i_28 : AND2_73 port map( A => A(28), B => n38, Y => 
                           A_shifter_28_port);
   SHIFTER_A_i_29 : AND2_72 port map( A => A(29), B => n38, Y => 
                           A_shifter_29_port);
   SHIFTER_A_i_30 : AND2_71 port map( A => A(30), B => n38, Y => 
                           A_shifter_30_port);
   SHIFTER_A_i_31 : AND2_70 port map( A => A(31), B => n38, Y => 
                           A_shifter_31_port);
   SHIFTER_B_i_0 : AND2_69 port map( A => B(0), B => n38, Y => B_shifter_0_port
                           );
   SHIFTER_B_i_1 : AND2_68 port map( A => B(1), B => n39, Y => B_shifter_1_port
                           );
   SHIFTER_B_i_2 : AND2_67 port map( A => B(2), B => n39, Y => B_shifter_2_port
                           );
   SHIFTER_B_i_3 : AND2_66 port map( A => B(3), B => n39, Y => B_shifter_3_port
                           );
   SHIFTER_B_i_4 : AND2_65 port map( A => B(4), B => n39, Y => B_shifter_4_port
                           );
   SUM_i_0 : AND2_64 port map( A => out_adder_0_port, B => n35, Y => 
                           in_cmp_0_port);
   SUM_i_1 : AND2_63 port map( A => out_adder_1_port, B => n35, Y => 
                           in_cmp_1_port);
   SUM_i_2 : AND2_62 port map( A => out_adder_2_port, B => n34, Y => 
                           in_cmp_2_port);
   SUM_i_3 : AND2_61 port map( A => out_adder_3_port, B => n34, Y => 
                           in_cmp_3_port);
   SUM_i_4 : AND2_60 port map( A => out_adder_4_port, B => n34, Y => 
                           in_cmp_4_port);
   SUM_i_5 : AND2_59 port map( A => out_adder_5_port, B => n34, Y => 
                           in_cmp_5_port);
   SUM_i_6 : AND2_58 port map( A => out_adder_6_port, B => n34, Y => 
                           in_cmp_6_port);
   SUM_i_7 : AND2_57 port map( A => out_adder_7_port, B => n34, Y => 
                           in_cmp_7_port);
   SUM_i_8 : AND2_56 port map( A => out_adder_8_port, B => n34, Y => 
                           in_cmp_8_port);
   SUM_i_9 : AND2_55 port map( A => out_adder_9_port, B => n34, Y => 
                           in_cmp_9_port);
   SUM_i_10 : AND2_54 port map( A => out_adder_10_port, B => n34, Y => 
                           in_cmp_10_port);
   SUM_i_11 : AND2_53 port map( A => out_adder_11_port, B => n34, Y => 
                           in_cmp_11_port);
   SUM_i_12 : AND2_52 port map( A => out_adder_12_port, B => n34, Y => 
                           in_cmp_12_port);
   SUM_i_13 : AND2_51 port map( A => out_adder_13_port, B => n34, Y => 
                           in_cmp_13_port);
   SUM_i_14 : AND2_50 port map( A => out_adder_14_port, B => n34, Y => 
                           in_cmp_14_port);
   SUM_i_15 : AND2_49 port map( A => out_adder_15_port, B => n34, Y => 
                           in_cmp_15_port);
   SUM_i_16 : AND2_48 port map( A => out_adder_16_port, B => n34, Y => 
                           in_cmp_16_port);
   SUM_i_17 : AND2_47 port map( A => out_adder_17_port, B => n34, Y => 
                           in_cmp_17_port);
   SUM_i_18 : AND2_46 port map( A => out_adder_18_port, B => n33, Y => 
                           in_cmp_18_port);
   SUM_i_19 : AND2_45 port map( A => out_adder_19_port, B => n33, Y => 
                           in_cmp_19_port);
   SUM_i_20 : AND2_44 port map( A => out_adder_20_port, B => n33, Y => 
                           in_cmp_20_port);
   SUM_i_21 : AND2_43 port map( A => out_adder_21_port, B => n33, Y => 
                           in_cmp_21_port);
   SUM_i_22 : AND2_42 port map( A => out_adder_22_port, B => n33, Y => 
                           in_cmp_22_port);
   SUM_i_23 : AND2_41 port map( A => out_adder_23_port, B => n33, Y => 
                           in_cmp_23_port);
   SUM_i_24 : AND2_40 port map( A => out_adder_24_port, B => n33, Y => 
                           in_cmp_24_port);
   SUM_i_25 : AND2_39 port map( A => out_adder_25_port, B => n33, Y => 
                           in_cmp_25_port);
   SUM_i_26 : AND2_38 port map( A => out_adder_26_port, B => n33, Y => 
                           in_cmp_26_port);
   SUM_i_27 : AND2_37 port map( A => out_adder_27_port, B => n33, Y => 
                           in_cmp_27_port);
   SUM_i_28 : AND2_36 port map( A => out_adder_28_port, B => n33, Y => 
                           in_cmp_28_port);
   SUM_i_29 : AND2_35 port map( A => out_adder_29_port, B => n33, Y => 
                           in_cmp_29_port);
   SUM_i_30 : AND2_34 port map( A => out_adder_30_port, B => n33, Y => 
                           in_cmp_30_port);
   SUM_i_31 : AND2_33 port map( A => out_adder_31_port, B => n33, Y => 
                           in_cmp_31_port);
   MUL_A_i_0 : AND2_32 port map( A => A(0), B => n8, Y => A_mul_0_port);
   MUL_B_i_0 : AND2_31 port map( A => B(0), B => n8, Y => B_mul_0_port);
   MUL_A_i_1 : AND2_30 port map( A => A(1), B => n8, Y => A_mul_1_port);
   MUL_B_i_1 : AND2_29 port map( A => B(1), B => n8, Y => B_mul_1_port);
   MUL_A_i_2 : AND2_28 port map( A => A(2), B => n8, Y => A_mul_2_port);
   MUL_B_i_2 : AND2_27 port map( A => B(2), B => n8, Y => B_mul_2_port);
   MUL_A_i_3 : AND2_26 port map( A => A(3), B => n8, Y => A_mul_3_port);
   MUL_B_i_3 : AND2_25 port map( A => B(3), B => n8, Y => B_mul_3_port);
   MUL_A_i_4 : AND2_24 port map( A => A(4), B => n8, Y => A_mul_4_port);
   MUL_B_i_4 : AND2_23 port map( A => B(4), B => n8, Y => B_mul_4_port);
   MUL_A_i_5 : AND2_22 port map( A => A(5), B => n8, Y => A_mul_5_port);
   MUL_B_i_5 : AND2_21 port map( A => B(5), B => n9, Y => B_mul_5_port);
   MUL_A_i_6 : AND2_20 port map( A => A(6), B => n9, Y => A_mul_6_port);
   MUL_B_i_6 : AND2_19 port map( A => B(6), B => n9, Y => B_mul_6_port);
   MUL_A_i_7 : AND2_18 port map( A => A(7), B => n9, Y => A_mul_7_port);
   MUL_B_i_7 : AND2_17 port map( A => B(7), B => n9, Y => B_mul_7_port);
   MUL_A_i_8 : AND2_16 port map( A => A(8), B => n9, Y => A_mul_8_port);
   MUL_B_i_8 : AND2_15 port map( A => B(8), B => n9, Y => B_mul_8_port);
   MUL_A_i_9 : AND2_14 port map( A => A(9), B => n9, Y => A_mul_9_port);
   MUL_B_i_9 : AND2_13 port map( A => B(9), B => n9, Y => B_mul_9_port);
   MUL_A_i_10 : AND2_12 port map( A => A(10), B => n9, Y => A_mul_10_port);
   MUL_B_i_10 : AND2_11 port map( A => B(10), B => n9, Y => B_mul_10_port);
   MUL_A_i_11 : AND2_10 port map( A => A(11), B => n30, Y => A_mul_11_port);
   MUL_B_i_11 : AND2_9 port map( A => B(11), B => n30, Y => B_mul_11_port);
   MUL_A_i_12 : AND2_8 port map( A => A(12), B => n30, Y => A_mul_12_port);
   MUL_B_i_12 : AND2_7 port map( A => B(12), B => n30, Y => B_mul_12_port);
   MUL_A_i_13 : AND2_6 port map( A => A(13), B => n30, Y => A_mul_13_port);
   MUL_B_i_13 : AND2_5 port map( A => B(13), B => n30, Y => B_mul_13_port);
   MUL_A_i_14 : AND2_4 port map( A => A(14), B => n30, Y => A_mul_14_port);
   MUL_B_i_14 : AND2_3 port map( A => B(14), B => n30, Y => B_mul_14_port);
   MUL_A_i_15 : AND2_2 port map( A => A(15), B => n30, Y => A_mul_15_port);
   MUL_B_i_15 : AND2_1 port map( A => B(15), B => n30, Y => B_mul_15_port);
   ADD : ADDER_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A_adder_31_port, 
                           A(30) => A_adder_30_port, A(29) => A_adder_29_port, 
                           A(28) => A_adder_28_port, A(27) => A_adder_27_port, 
                           A(26) => A_adder_26_port, A(25) => A_adder_25_port, 
                           A(24) => A_adder_24_port, A(23) => A_adder_23_port, 
                           A(22) => A_adder_22_port, A(21) => A_adder_21_port, 
                           A(20) => A_adder_20_port, A(19) => A_adder_19_port, 
                           A(18) => A_adder_18_port, A(17) => A_adder_17_port, 
                           A(16) => A_adder_16_port, A(15) => A_adder_15_port, 
                           A(14) => A_adder_14_port, A(13) => A_adder_13_port, 
                           A(12) => A_adder_12_port, A(11) => A_adder_11_port, 
                           A(10) => A_adder_10_port, A(9) => A_adder_9_port, 
                           A(8) => A_adder_8_port, A(7) => A_adder_7_port, A(6)
                           => A_adder_6_port, A(5) => A_adder_5_port, A(4) => 
                           A_adder_4_port, A(3) => A_adder_3_port, A(2) => 
                           A_adder_2_port, A(1) => A_adder_1_port, A(0) => 
                           A_adder_0_port, B(31) => B_adder_31_port, B(30) => 
                           B_adder_30_port, B(29) => B_adder_29_port, B(28) => 
                           B_adder_28_port, B(27) => B_adder_27_port, B(26) => 
                           B_adder_26_port, B(25) => B_adder_25_port, B(24) => 
                           B_adder_24_port, B(23) => B_adder_23_port, B(22) => 
                           B_adder_22_port, B(21) => B_adder_21_port, B(20) => 
                           B_adder_20_port, B(19) => B_adder_19_port, B(18) => 
                           B_adder_18_port, B(17) => B_adder_17_port, B(16) => 
                           B_adder_16_port, B(15) => B_adder_15_port, B(14) => 
                           B_adder_14_port, B(13) => B_adder_13_port, B(12) => 
                           B_adder_12_port, B(11) => B_adder_11_port, B(10) => 
                           B_adder_10_port, B(9) => B_adder_9_port, B(8) => 
                           B_adder_8_port, B(7) => B_adder_7_port, B(6) => 
                           B_adder_6_port, B(5) => B_adder_5_port, B(4) => 
                           B_adder_4_port, B(3) => B_adder_3_port, B(2) => 
                           B_adder_2_port, B(1) => B_adder_1_port, B(0) => 
                           B_adder_0_port, ADD_SUB => n55, Cin => cin_internal,
                           S(31) => out_adder_31_port, S(30) => 
                           out_adder_30_port, S(29) => out_adder_29_port, S(28)
                           => out_adder_28_port, S(27) => out_adder_27_port, 
                           S(26) => out_adder_26_port, S(25) => 
                           out_adder_25_port, S(24) => out_adder_24_port, S(23)
                           => out_adder_23_port, S(22) => out_adder_22_port, 
                           S(21) => out_adder_21_port, S(20) => 
                           out_adder_20_port, S(19) => out_adder_19_port, S(18)
                           => out_adder_18_port, S(17) => out_adder_17_port, 
                           S(16) => out_adder_16_port, S(15) => 
                           out_adder_15_port, S(14) => out_adder_14_port, S(13)
                           => out_adder_13_port, S(12) => out_adder_12_port, 
                           S(11) => out_adder_11_port, S(10) => 
                           out_adder_10_port, S(9) => out_adder_9_port, S(8) =>
                           out_adder_8_port, S(7) => out_adder_7_port, S(6) => 
                           out_adder_6_port, S(5) => out_adder_5_port, S(4) => 
                           out_adder_4_port, S(3) => out_adder_3_port, S(2) => 
                           out_adder_2_port, S(1) => out_adder_1_port, S(0) => 
                           out_adder_0_port, Cout => Cout_port);
   SHIFT : SHIFTER port map( data_in(31) => A_shifter_31_port, data_in(30) => 
                           A_shifter_30_port, data_in(29) => A_shifter_29_port,
                           data_in(28) => A_shifter_28_port, data_in(27) => 
                           A_shifter_27_port, data_in(26) => A_shifter_26_port,
                           data_in(25) => A_shifter_25_port, data_in(24) => 
                           A_shifter_24_port, data_in(23) => A_shifter_23_port,
                           data_in(22) => A_shifter_22_port, data_in(21) => 
                           A_shifter_21_port, data_in(20) => A_shifter_20_port,
                           data_in(19) => A_shifter_19_port, data_in(18) => 
                           A_shifter_18_port, data_in(17) => A_shifter_17_port,
                           data_in(16) => A_shifter_16_port, data_in(15) => 
                           A_shifter_15_port, data_in(14) => A_shifter_14_port,
                           data_in(13) => A_shifter_13_port, data_in(12) => 
                           A_shifter_12_port, data_in(11) => A_shifter_11_port,
                           data_in(10) => A_shifter_10_port, data_in(9) => 
                           A_shifter_9_port, data_in(8) => A_shifter_8_port, 
                           data_in(7) => A_shifter_7_port, data_in(6) => 
                           A_shifter_6_port, data_in(5) => A_shifter_5_port, 
                           data_in(4) => A_shifter_4_port, data_in(3) => 
                           A_shifter_3_port, data_in(2) => A_shifter_2_port, 
                           data_in(1) => A_shifter_1_port, data_in(0) => 
                           A_shifter_0_port, R(4) => B_shifter_4_port, R(3) => 
                           B_shifter_3_port, R(2) => B_shifter_2_port, R(1) => 
                           B_shifter_1_port, R(0) => B_shifter_0_port, conf(1) 
                           => conf_1_port, conf(0) => conf_0_port, data_out(31)
                           => out_shifter_31_port, data_out(30) => 
                           out_shifter_30_port, data_out(29) => 
                           out_shifter_29_port, data_out(28) => 
                           out_shifter_28_port, data_out(27) => 
                           out_shifter_27_port, data_out(26) => 
                           out_shifter_26_port, data_out(25) => 
                           out_shifter_25_port, data_out(24) => 
                           out_shifter_24_port, data_out(23) => 
                           out_shifter_23_port, data_out(22) => 
                           out_shifter_22_port, data_out(21) => 
                           out_shifter_21_port, data_out(20) => 
                           out_shifter_20_port, data_out(19) => 
                           out_shifter_19_port, data_out(18) => 
                           out_shifter_18_port, data_out(17) => 
                           out_shifter_17_port, data_out(16) => 
                           out_shifter_16_port, data_out(15) => 
                           out_shifter_15_port, data_out(14) => 
                           out_shifter_14_port, data_out(13) => 
                           out_shifter_13_port, data_out(12) => 
                           out_shifter_12_port, data_out(11) => 
                           out_shifter_11_port, data_out(10) => 
                           out_shifter_10_port, data_out(9) => 
                           out_shifter_9_port, data_out(8) => 
                           out_shifter_8_port, data_out(7) => 
                           out_shifter_7_port, data_out(6) => 
                           out_shifter_6_port, data_out(5) => 
                           out_shifter_5_port, data_out(4) => 
                           out_shifter_4_port, data_out(3) => 
                           out_shifter_3_port, data_out(2) => 
                           out_shifter_2_port, data_out(1) => 
                           out_shifter_1_port, data_out(0) => 
                           out_shifter_0_port);
   LOGICALS : LOGIC_NBIT32_N_SELECTOR4 port map( S(3) => logic_sel_3_port, S(2)
                           => logic_sel_2_port, S(1) => logic_sel_1_port, S(0) 
                           => logic_sel_0_port, A(31) => A_logic_31_port, A(30)
                           => A_logic_30_port, A(29) => A_logic_29_port, A(28) 
                           => A_logic_28_port, A(27) => A_logic_27_port, A(26) 
                           => A_logic_26_port, A(25) => A_logic_25_port, A(24) 
                           => A_logic_24_port, A(23) => A_logic_23_port, A(22) 
                           => A_logic_22_port, A(21) => A_logic_21_port, A(20) 
                           => A_logic_20_port, A(19) => A_logic_19_port, A(18) 
                           => A_logic_18_port, A(17) => A_logic_17_port, A(16) 
                           => A_logic_16_port, A(15) => A_logic_15_port, A(14) 
                           => A_logic_14_port, A(13) => A_logic_13_port, A(12) 
                           => A_logic_12_port, A(11) => A_logic_11_port, A(10) 
                           => A_logic_10_port, A(9) => A_logic_9_port, A(8) => 
                           A_logic_8_port, A(7) => A_logic_7_port, A(6) => 
                           A_logic_6_port, A(5) => A_logic_5_port, A(4) => 
                           A_logic_4_port, A(3) => A_logic_3_port, A(2) => 
                           A_logic_2_port, A(1) => A_logic_1_port, A(0) => 
                           A_logic_0_port, B(31) => B_logic_31_port, B(30) => 
                           B_logic_30_port, B(29) => B_logic_29_port, B(28) => 
                           B_logic_28_port, B(27) => B_logic_27_port, B(26) => 
                           B_logic_26_port, B(25) => B_logic_25_port, B(24) => 
                           B_logic_24_port, B(23) => B_logic_23_port, B(22) => 
                           B_logic_22_port, B(21) => B_logic_21_port, B(20) => 
                           B_logic_20_port, B(19) => B_logic_19_port, B(18) => 
                           B_logic_18_port, B(17) => B_logic_17_port, B(16) => 
                           B_logic_16_port, B(15) => B_logic_15_port, B(14) => 
                           B_logic_14_port, B(13) => B_logic_13_port, B(12) => 
                           B_logic_12_port, B(11) => B_logic_11_port, B(10) => 
                           B_logic_10_port, B(9) => B_logic_9_port, B(8) => 
                           B_logic_8_port, B(7) => B_logic_7_port, B(6) => 
                           B_logic_6_port, B(5) => B_logic_5_port, B(4) => 
                           B_logic_4_port, B(3) => B_logic_3_port, B(2) => 
                           B_logic_2_port, B(1) => B_logic_1_port, B(0) => 
                           B_logic_0_port, O(31) => out_logic_31_port, O(30) =>
                           out_logic_30_port, O(29) => out_logic_29_port, O(28)
                           => out_logic_28_port, O(27) => out_logic_27_port, 
                           O(26) => out_logic_26_port, O(25) => 
                           out_logic_25_port, O(24) => out_logic_24_port, O(23)
                           => out_logic_23_port, O(22) => out_logic_22_port, 
                           O(21) => out_logic_21_port, O(20) => 
                           out_logic_20_port, O(19) => out_logic_19_port, O(18)
                           => out_logic_18_port, O(17) => out_logic_17_port, 
                           O(16) => out_logic_16_port, O(15) => 
                           out_logic_15_port, O(14) => out_logic_14_port, O(13)
                           => out_logic_13_port, O(12) => out_logic_12_port, 
                           O(11) => out_logic_11_port, O(10) => 
                           out_logic_10_port, O(9) => out_logic_9_port, O(8) =>
                           out_logic_8_port, O(7) => out_logic_7_port, O(6) => 
                           out_logic_6_port, O(5) => out_logic_5_port, O(4) => 
                           out_logic_4_port, O(3) => out_logic_3_port, O(2) => 
                           out_logic_2_port, O(1) => out_logic_1_port, O(0) => 
                           out_logic_0_port);
   COMPARATOR : CMP_NBIT32 port map( SUM(31) => in_cmp_31_port, SUM(30) => 
                           in_cmp_30_port, SUM(29) => in_cmp_29_port, SUM(28) 
                           => in_cmp_28_port, SUM(27) => in_cmp_27_port, 
                           SUM(26) => in_cmp_26_port, SUM(25) => in_cmp_25_port
                           , SUM(24) => in_cmp_24_port, SUM(23) => 
                           in_cmp_23_port, SUM(22) => in_cmp_22_port, SUM(21) 
                           => in_cmp_21_port, SUM(20) => in_cmp_20_port, 
                           SUM(19) => in_cmp_19_port, SUM(18) => in_cmp_18_port
                           , SUM(17) => in_cmp_17_port, SUM(16) => 
                           in_cmp_16_port, SUM(15) => in_cmp_15_port, SUM(14) 
                           => in_cmp_14_port, SUM(13) => in_cmp_13_port, 
                           SUM(12) => in_cmp_12_port, SUM(11) => in_cmp_11_port
                           , SUM(10) => in_cmp_10_port, SUM(9) => in_cmp_9_port
                           , SUM(8) => in_cmp_8_port, SUM(7) => in_cmp_7_port, 
                           SUM(6) => in_cmp_6_port, SUM(5) => in_cmp_5_port, 
                           SUM(4) => in_cmp_4_port, SUM(3) => in_cmp_3_port, 
                           SUM(2) => in_cmp_2_port, SUM(1) => in_cmp_1_port, 
                           SUM(0) => in_cmp_0_port, Cout => Cout_port, A_L_B =>
                           COND(0), A_LE_B => COND(1), A_G_B => COND(2), A_GE_B
                           => COND(3), A_E_B => COND(4), A_NE_B => COND(5));
   MULTIPLIER : MUL port map( CLOCK => CLOCK, A(15) => A_mul_15_port, A(14) => 
                           A_mul_14_port, A(13) => A_mul_13_port, A(12) => 
                           A_mul_12_port, A(11) => A_mul_11_port, A(10) => 
                           A_mul_10_port, A(9) => A_mul_9_port, A(8) => 
                           A_mul_8_port, A(7) => A_mul_7_port, A(6) => 
                           A_mul_6_port, A(5) => A_mul_5_port, A(4) => 
                           A_mul_4_port, A(3) => A_mul_3_port, A(2) => 
                           A_mul_2_port, A(1) => A_mul_1_port, A(0) => 
                           A_mul_0_port, B(15) => B_mul_15_port, B(14) => 
                           B_mul_14_port, B(13) => B_mul_13_port, B(12) => 
                           B_mul_12_port, B(11) => B_mul_11_port, B(10) => 
                           B_mul_10_port, B(9) => B_mul_9_port, B(8) => 
                           B_mul_8_port, B(7) => B_mul_7_port, B(6) => 
                           B_mul_6_port, B(5) => B_mul_5_port, B(4) => 
                           B_mul_4_port, B(3) => B_mul_3_port, B(2) => 
                           B_mul_2_port, B(1) => B_mul_1_port, B(0) => 
                           B_mul_0_port, Y(31) => out_mul_31_port, Y(30) => 
                           out_mul_30_port, Y(29) => out_mul_29_port, Y(28) => 
                           out_mul_28_port, Y(27) => out_mul_27_port, Y(26) => 
                           out_mul_26_port, Y(25) => out_mul_25_port, Y(24) => 
                           out_mul_24_port, Y(23) => out_mul_23_port, Y(22) => 
                           out_mul_22_port, Y(21) => out_mul_21_port, Y(20) => 
                           out_mul_20_port, Y(19) => out_mul_19_port, Y(18) => 
                           out_mul_18_port, Y(17) => out_mul_17_port, Y(16) => 
                           out_mul_16_port, Y(15) => out_mul_15_port, Y(14) => 
                           out_mul_14_port, Y(13) => out_mul_13_port, Y(12) => 
                           out_mul_12_port, Y(11) => out_mul_11_port, Y(10) => 
                           out_mul_10_port, Y(9) => out_mul_9_port, Y(8) => 
                           out_mul_8_port, Y(7) => out_mul_7_port, Y(6) => 
                           out_mul_6_port, Y(5) => out_mul_5_port, Y(4) => 
                           out_mul_4_port, Y(3) => out_mul_3_port, Y(2) => 
                           out_mul_2_port, Y(1) => out_mul_1_port, Y(0) => 
                           out_mul_0_port);
   OUTPUT_SEL : MUX4to1_NBIT32_1 port map( A(31) => out_adder_31_port, A(30) =>
                           out_adder_30_port, A(29) => out_adder_29_port, A(28)
                           => out_adder_28_port, A(27) => out_adder_27_port, 
                           A(26) => out_adder_26_port, A(25) => 
                           out_adder_25_port, A(24) => out_adder_24_port, A(23)
                           => out_adder_23_port, A(22) => out_adder_22_port, 
                           A(21) => out_adder_21_port, A(20) => 
                           out_adder_20_port, A(19) => out_adder_19_port, A(18)
                           => out_adder_18_port, A(17) => out_adder_17_port, 
                           A(16) => out_adder_16_port, A(15) => 
                           out_adder_15_port, A(14) => out_adder_14_port, A(13)
                           => out_adder_13_port, A(12) => out_adder_12_port, 
                           A(11) => out_adder_11_port, A(10) => 
                           out_adder_10_port, A(9) => out_adder_9_port, A(8) =>
                           out_adder_8_port, A(7) => out_adder_7_port, A(6) => 
                           out_adder_6_port, A(5) => out_adder_5_port, A(4) => 
                           out_adder_4_port, A(3) => out_adder_3_port, A(2) => 
                           out_adder_2_port, A(1) => out_adder_1_port, A(0) => 
                           out_adder_0_port, B(31) => out_logic_31_port, B(30) 
                           => out_logic_30_port, B(29) => out_logic_29_port, 
                           B(28) => out_logic_28_port, B(27) => 
                           out_logic_27_port, B(26) => out_logic_26_port, B(25)
                           => out_logic_25_port, B(24) => out_logic_24_port, 
                           B(23) => out_logic_23_port, B(22) => 
                           out_logic_22_port, B(21) => out_logic_21_port, B(20)
                           => out_logic_20_port, B(19) => out_logic_19_port, 
                           B(18) => out_logic_18_port, B(17) => 
                           out_logic_17_port, B(16) => out_logic_16_port, B(15)
                           => out_logic_15_port, B(14) => out_logic_14_port, 
                           B(13) => out_logic_13_port, B(12) => 
                           out_logic_12_port, B(11) => out_logic_11_port, B(10)
                           => out_logic_10_port, B(9) => out_logic_9_port, B(8)
                           => out_logic_8_port, B(7) => out_logic_7_port, B(6) 
                           => out_logic_6_port, B(5) => out_logic_5_port, B(4) 
                           => out_logic_4_port, B(3) => out_logic_3_port, B(2) 
                           => out_logic_2_port, B(1) => out_logic_1_port, B(0) 
                           => out_logic_0_port, C(31) => out_shifter_31_port, 
                           C(30) => out_shifter_30_port, C(29) => 
                           out_shifter_29_port, C(28) => out_shifter_28_port, 
                           C(27) => out_shifter_27_port, C(26) => 
                           out_shifter_26_port, C(25) => out_shifter_25_port, 
                           C(24) => out_shifter_24_port, C(23) => 
                           out_shifter_23_port, C(22) => out_shifter_22_port, 
                           C(21) => out_shifter_21_port, C(20) => 
                           out_shifter_20_port, C(19) => out_shifter_19_port, 
                           C(18) => out_shifter_18_port, C(17) => 
                           out_shifter_17_port, C(16) => out_shifter_16_port, 
                           C(15) => out_shifter_15_port, C(14) => 
                           out_shifter_14_port, C(13) => out_shifter_13_port, 
                           C(12) => out_shifter_12_port, C(11) => 
                           out_shifter_11_port, C(10) => out_shifter_10_port, 
                           C(9) => out_shifter_9_port, C(8) => 
                           out_shifter_8_port, C(7) => out_shifter_7_port, C(6)
                           => out_shifter_6_port, C(5) => out_shifter_5_port, 
                           C(4) => out_shifter_4_port, C(3) => 
                           out_shifter_3_port, C(2) => out_shifter_2_port, C(1)
                           => out_shifter_1_port, C(0) => out_shifter_0_port, 
                           D(31) => out_mul_31_port, D(30) => out_mul_30_port, 
                           D(29) => out_mul_29_port, D(28) => out_mul_28_port, 
                           D(27) => out_mul_27_port, D(26) => out_mul_26_port, 
                           D(25) => out_mul_25_port, D(24) => out_mul_24_port, 
                           D(23) => out_mul_23_port, D(22) => out_mul_22_port, 
                           D(21) => out_mul_21_port, D(20) => out_mul_20_port, 
                           D(19) => out_mul_19_port, D(18) => out_mul_18_port, 
                           D(17) => out_mul_17_port, D(16) => out_mul_16_port, 
                           D(15) => out_mul_15_port, D(14) => out_mul_14_port, 
                           D(13) => out_mul_13_port, D(12) => out_mul_12_port, 
                           D(11) => out_mul_11_port, D(10) => out_mul_10_port, 
                           D(9) => out_mul_9_port, D(8) => out_mul_8_port, D(7)
                           => out_mul_7_port, D(6) => out_mul_6_port, D(5) => 
                           out_mul_5_port, D(4) => out_mul_4_port, D(3) => 
                           out_mul_3_port, D(2) => out_mul_2_port, D(1) => 
                           out_mul_1_port, D(0) => out_mul_0_port, SEL(1) => 
                           mux_out_1_port, SEL(0) => mux_out_0_port, Y(31) => 
                           ALU_out(31), Y(30) => ALU_out(30), Y(29) => 
                           ALU_out(29), Y(28) => ALU_out(28), Y(27) => 
                           ALU_out(27), Y(26) => ALU_out(26), Y(25) => 
                           ALU_out(25), Y(24) => ALU_out(24), Y(23) => 
                           ALU_out(23), Y(22) => ALU_out(22), Y(21) => 
                           ALU_out(21), Y(20) => ALU_out(20), Y(19) => 
                           ALU_out(19), Y(18) => ALU_out(18), Y(17) => 
                           ALU_out(17), Y(16) => ALU_out(16), Y(15) => 
                           ALU_out(15), Y(14) => ALU_out(14), Y(13) => 
                           ALU_out(13), Y(12) => ALU_out(12), Y(11) => 
                           ALU_out(11), Y(10) => ALU_out(10), Y(9) => 
                           ALU_out(9), Y(8) => ALU_out(8), Y(7) => ALU_out(7), 
                           Y(6) => ALU_out(6), Y(5) => ALU_out(5), Y(4) => 
                           ALU_out(4), Y(3) => ALU_out(3), Y(2) => ALU_out(2), 
                           Y(1) => ALU_out(1), Y(0) => ALU_out(0));
   U3 : BUF_X1 port map( A => en_adder, Z => n7);
   U4 : BUF_X1 port map( A => en_cmp, Z => n33);
   U5 : BUF_X1 port map( A => n5, Z => n2);
   U6 : BUF_X1 port map( A => n1, Z => n31);
   U7 : BUF_X1 port map( A => en_adder, Z => n4);
   U8 : BUF_X1 port map( A => en_adder, Z => n3);
   U9 : AND3_X1 port map( A1 => n58, A2 => n60, A3 => n11, ZN => n1);
   U10 : BUF_X1 port map( A => n43, Z => n52);
   U11 : BUF_X1 port map( A => n43, Z => n51);
   U12 : OR2_X1 port map( A1 => n30, A2 => n49, ZN => mux_out_0_port);
   U13 : BUF_X1 port map( A => n31, Z => n30);
   U14 : BUF_X1 port map( A => n40, Z => n39);
   U15 : OR2_X1 port map( A1 => n32, A2 => n39, ZN => mux_out_1_port);
   U16 : BUF_X1 port map( A => n40, Z => n38);
   U17 : BUF_X1 port map( A => n40, Z => n37);
   U18 : BUF_X1 port map( A => n31, Z => n9);
   U19 : BUF_X1 port map( A => n42, Z => n40);
   U20 : BUF_X1 port map( A => n51, Z => n49);
   U21 : BUF_X1 port map( A => n51, Z => n48);
   U22 : BUF_X1 port map( A => n52, Z => n46);
   U23 : BUF_X1 port map( A => n52, Z => n45);
   U24 : BUF_X1 port map( A => n52, Z => n47);
   U25 : BUF_X1 port map( A => n41, Z => n36);
   U26 : BUF_X1 port map( A => n42, Z => n41);
   U27 : BUF_X1 port map( A => n51, Z => n50);
   U28 : BUF_X1 port map( A => n32, Z => n8);
   U29 : BUF_X1 port map( A => n1, Z => n32);
   U30 : BUF_X1 port map( A => en_adder, Z => n6);
   U31 : INV_X1 port map( A => n22, ZN => n58);
   U32 : BUF_X1 port map( A => en_shifter, Z => n42);
   U33 : BUF_X1 port map( A => n53, Z => n44);
   U34 : BUF_X1 port map( A => n43, Z => n53);
   U35 : NOR3_X1 port map( A1 => n59, A2 => n62, A3 => n10, ZN => N92);
   U36 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => N88);
   U46 : NAND2_X1 port map( A1 => Cin, A2 => n15, ZN => n16);
   U47 : INV_X1 port map( A => AluOpcode(4), ZN => n62);
   U48 : BUF_X1 port map( A => en_logic, Z => n43);
   U49 : INV_X1 port map( A => N89, ZN => n54);
   U50 : NOR3_X1 port map( A1 => n22, A2 => n11, A3 => n23, ZN => N90);
   U51 : BUF_X1 port map( A => en_adder, Z => n5);
   U52 : INV_X1 port map( A => AluOpcode(3), ZN => n61);
   U53 : NAND2_X1 port map( A1 => AluOpcode(4), A2 => n59, ZN => n22);
   U54 : NOR3_X1 port map( A1 => n10, A2 => AluOpcode(1), A3 => AluOpcode(4), 
                           ZN => N93);
   U55 : INV_X1 port map( A => AluOpcode(1), ZN => n59);
   U56 : CLKBUF_X1 port map( A => en_cmp, Z => n34);
   U57 : CLKBUF_X1 port map( A => en_cmp, Z => n35);
   U58 : INV_X1 port map( A => AluOpcode(0), ZN => n57);
   U59 : NAND4_X1 port map( A1 => n26, A2 => n24, A3 => n25, A4 => n54, ZN => 
                           en_logic);
   U60 : AOI22_X1 port map( A1 => n21, A2 => n62, B1 => AluOpcode(1), B2 => 
                           AluOpcode(2), ZN => n20);
   U61 : NAND2_X1 port map( A1 => AluOpcode(2), A2 => n19, ZN => n10);
   U62 : NOR2_X1 port map( A1 => AluOpcode(1), A2 => AluOpcode(2), ZN => n15);
   U63 : INV_X1 port map( A => AluOpcode(2), ZN => n60);
   U64 : OAI22_X1 port map( A1 => n15, A2 => n57, B1 => AluOpcode(3), B2 => n20
                           , ZN => N91);
   U65 : NAND4_X1 port map( A1 => n58, A2 => AluOpcode(3), A3 => n60, A4 => n57
                           , ZN => n26);
   U66 : NAND4_X1 port map( A1 => n58, A2 => AluOpcode(2), A3 => n61, A4 => n57
                           , ZN => n27);
   U67 : NOR2_X1 port map( A1 => n57, A2 => n61, ZN => n11);
   U68 : INV_X1 port map( A => n17, ZN => n56);
   U69 : NOR2_X1 port map( A1 => AluOpcode(0), A2 => AluOpcode(1), ZN => n21);
   U70 : NOR4_X1 port map( A1 => n16, A2 => n61, A3 => AluOpcode(0), A4 => 
                           AluOpcode(4), ZN => cin_internal);
   U71 : NAND4_X1 port map( A1 => n58, A2 => AluOpcode(0), A3 => n61, A4 => n60
                           , ZN => n24);
   U72 : NOR2_X1 port map( A1 => AluOpcode(3), A2 => AluOpcode(0), ZN => n19);
   U73 : NOR2_X1 port map( A1 => n10, A2 => n58, ZN => en_shifter);
   U74 : INV_X1 port map( A => n13, ZN => n55);
   U75 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => en_adder);
   U76 : AOI21_X1 port map( B1 => n62, B2 => n56, A => n33, ZN => n13);
   U77 : OAI21_X1 port map( B1 => AluOpcode(1), B2 => n17, A => n18, ZN => 
                           en_cmp);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT5 is

   port( A, B, C : in std_logic_vector (4 downto 0);  SEL : in std_logic_vector
         (1 downto 0);  Y : out std_logic_vector (4 downto 0));

end MUX3to1_NBIT5;

architecture SYN_Behavioral of MUX3to1_NBIT5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n7, n8, n9, n10, n11, n12_port, n13, n14, n1, n2, n3, n4, n5, n6
      : std_logic;

begin
   
   Y_reg_4_inst : DLH_X1 port map( G => N12, D => n1, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => N12, D => n2, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => N12, D => n3, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => n4, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => n5, Q => Y(0));
   U3 : NOR2_X1 port map( A1 => n6, A2 => SEL(0), ZN => n9);
   U4 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n8);
   U5 : AND2_X1 port map( A1 => SEL(0), A2 => n6, ZN => n10);
   U6 : NAND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => N12);
   U7 : INV_X1 port map( A => SEL(1), ZN => n6);
   U8 : INV_X1 port map( A => n14, ZN => n5);
   U9 : AOI222_X1 port map( A1 => A(0), A2 => n8, B1 => C(0), B2 => n9, C1 => 
                           B(0), C2 => n10, ZN => n14);
   U10 : INV_X1 port map( A => n13, ZN => n4);
   U11 : AOI222_X1 port map( A1 => A(1), A2 => n8, B1 => C(1), B2 => n9, C1 => 
                           B(1), C2 => n10, ZN => n13);
   U12 : INV_X1 port map( A => n12_port, ZN => n3);
   U13 : AOI222_X1 port map( A1 => A(2), A2 => n8, B1 => C(2), B2 => n9, C1 => 
                           B(2), C2 => n10, ZN => n12_port);
   U14 : INV_X1 port map( A => n11, ZN => n2);
   U15 : AOI222_X1 port map( A1 => A(3), A2 => n8, B1 => C(3), B2 => n9, C1 => 
                           B(3), C2 => n10, ZN => n11);
   U16 : INV_X1 port map( A => n7, ZN => n1);
   U17 : AOI222_X1 port map( A1 => A(4), A2 => n8, B1 => C(4), B2 => n9, C1 => 
                           B(4), C2 => n10, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX4to1_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX4to1_NBIT32_0;

architecture SYN_Behavioral of MUX4to1_NBIT32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n76);
   U2 : BUF_X1 port map( A => n7, Z => n72);
   U3 : BUF_X1 port map( A => n4, Z => n81);
   U4 : BUF_X1 port map( A => n5, Z => n77);
   U5 : BUF_X1 port map( A => n76, Z => n73);
   U6 : BUF_X1 port map( A => n76, Z => n74);
   U7 : BUF_X1 port map( A => n81, Z => n82);
   U8 : BUF_X1 port map( A => n81, Z => n83);
   U9 : BUF_X1 port map( A => n72, Z => n1);
   U10 : BUF_X1 port map( A => n72, Z => n70);
   U11 : BUF_X1 port map( A => n77, Z => n78);
   U12 : BUF_X1 port map( A => n77, Z => n79);
   U13 : BUF_X1 port map( A => n76, Z => n75);
   U14 : BUF_X1 port map( A => n81, Z => n84);
   U15 : BUF_X1 port map( A => n72, Z => n71);
   U16 : BUF_X1 port map( A => n77, Z => n80);
   U17 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(0));
   U18 : AOI22_X1 port map( A1 => D(0), A2 => n82, B1 => C(0), B2 => n78, ZN =>
                           n69);
   U19 : AOI22_X1 port map( A1 => B(0), A2 => n73, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U20 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(1));
   U21 : AOI22_X1 port map( A1 => D(1), A2 => n82, B1 => C(1), B2 => n78, ZN =>
                           n47);
   U22 : AOI22_X1 port map( A1 => B(1), A2 => n73, B1 => A(1), B2 => n1, ZN => 
                           n46);
   U23 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(2));
   U24 : AOI22_X1 port map( A1 => D(2), A2 => n83, B1 => C(2), B2 => n79, ZN =>
                           n25);
   U25 : AOI22_X1 port map( A1 => B(2), A2 => n74, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U26 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(3));
   U27 : AOI22_X1 port map( A1 => D(3), A2 => n84, B1 => C(3), B2 => n80, ZN =>
                           n19);
   U28 : AOI22_X1 port map( A1 => B(3), A2 => n75, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U29 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(4));
   U30 : AOI22_X1 port map( A1 => D(4), A2 => n84, B1 => C(4), B2 => n80, ZN =>
                           n17);
   U31 : AOI22_X1 port map( A1 => B(4), A2 => n75, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U32 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(5));
   U33 : AOI22_X1 port map( A1 => D(5), A2 => n84, B1 => C(5), B2 => n80, ZN =>
                           n15);
   U34 : AOI22_X1 port map( A1 => B(5), A2 => n75, B1 => A(5), B2 => n71, ZN =>
                           n14);
   U35 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(6));
   U36 : AOI22_X1 port map( A1 => D(6), A2 => n84, B1 => C(6), B2 => n80, ZN =>
                           n13);
   U37 : AOI22_X1 port map( A1 => B(6), A2 => n75, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U38 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(7));
   U39 : AOI22_X1 port map( A1 => D(7), A2 => n84, B1 => C(7), B2 => n80, ZN =>
                           n11);
   U40 : AOI22_X1 port map( A1 => B(7), A2 => n75, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U41 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(8));
   U42 : AOI22_X1 port map( A1 => D(8), A2 => n84, B1 => C(8), B2 => n80, ZN =>
                           n9);
   U43 : AOI22_X1 port map( A1 => B(8), A2 => n75, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U44 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(9));
   U45 : AOI22_X1 port map( A1 => D(9), A2 => n84, B1 => C(9), B2 => n80, ZN =>
                           n3);
   U46 : AOI22_X1 port map( A1 => B(9), A2 => n75, B1 => A(9), B2 => n71, ZN =>
                           n2);
   U47 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(10));
   U48 : AOI22_X1 port map( A1 => D(10), A2 => n82, B1 => C(10), B2 => n78, ZN 
                           => n67);
   U49 : AOI22_X1 port map( A1 => B(10), A2 => n73, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U50 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(11));
   U51 : AOI22_X1 port map( A1 => D(11), A2 => n82, B1 => C(11), B2 => n78, ZN 
                           => n65);
   U52 : AOI22_X1 port map( A1 => B(11), A2 => n73, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U53 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(12));
   U54 : AOI22_X1 port map( A1 => D(12), A2 => n82, B1 => C(12), B2 => n78, ZN 
                           => n63);
   U55 : AOI22_X1 port map( A1 => B(12), A2 => n73, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U56 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(13));
   U57 : AOI22_X1 port map( A1 => D(13), A2 => n82, B1 => C(13), B2 => n78, ZN 
                           => n61);
   U58 : AOI22_X1 port map( A1 => B(13), A2 => n73, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U59 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(14));
   U60 : AOI22_X1 port map( A1 => D(14), A2 => n82, B1 => C(14), B2 => n78, ZN 
                           => n59);
   U61 : AOI22_X1 port map( A1 => B(14), A2 => n73, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U62 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(15));
   U63 : AOI22_X1 port map( A1 => D(15), A2 => n82, B1 => C(15), B2 => n78, ZN 
                           => n57);
   U64 : AOI22_X1 port map( A1 => B(15), A2 => n73, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U65 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(27));
   U66 : AOI22_X1 port map( A1 => D(27), A2 => n83, B1 => C(27), B2 => n79, ZN 
                           => n31);
   U67 : AOI22_X1 port map( A1 => B(27), A2 => n74, B1 => A(27), B2 => n70, ZN 
                           => n30);
   U68 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(16));
   U69 : AOI22_X1 port map( A1 => B(16), A2 => n73, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U70 : AOI22_X1 port map( A1 => D(16), A2 => n82, B1 => C(16), B2 => n78, ZN 
                           => n55);
   U71 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(17));
   U72 : AOI22_X1 port map( A1 => B(17), A2 => n73, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U73 : AOI22_X1 port map( A1 => D(17), A2 => n82, B1 => C(17), B2 => n78, ZN 
                           => n53);
   U74 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(18));
   U75 : AOI22_X1 port map( A1 => B(18), A2 => n73, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U76 : AOI22_X1 port map( A1 => D(18), A2 => n82, B1 => C(18), B2 => n78, ZN 
                           => n51);
   U77 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(19));
   U78 : AOI22_X1 port map( A1 => B(19), A2 => n73, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U79 : AOI22_X1 port map( A1 => D(19), A2 => n82, B1 => C(19), B2 => n78, ZN 
                           => n49);
   U80 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(20));
   U81 : AOI22_X1 port map( A1 => B(20), A2 => n74, B1 => A(20), B2 => n70, ZN 
                           => n44);
   U82 : AOI22_X1 port map( A1 => D(20), A2 => n83, B1 => C(20), B2 => n79, ZN 
                           => n45);
   U83 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(21));
   U84 : AOI22_X1 port map( A1 => B(21), A2 => n74, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U85 : AOI22_X1 port map( A1 => D(21), A2 => n83, B1 => C(21), B2 => n79, ZN 
                           => n43);
   U86 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(22));
   U87 : AOI22_X1 port map( A1 => B(22), A2 => n74, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U88 : AOI22_X1 port map( A1 => D(22), A2 => n83, B1 => C(22), B2 => n79, ZN 
                           => n41);
   U89 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(23));
   U90 : AOI22_X1 port map( A1 => B(23), A2 => n74, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U91 : AOI22_X1 port map( A1 => D(23), A2 => n83, B1 => C(23), B2 => n79, ZN 
                           => n39);
   U92 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(24));
   U93 : AOI22_X1 port map( A1 => B(24), A2 => n74, B1 => A(24), B2 => n70, ZN 
                           => n36);
   U94 : AOI22_X1 port map( A1 => D(24), A2 => n83, B1 => C(24), B2 => n79, ZN 
                           => n37);
   U95 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(25));
   U96 : AOI22_X1 port map( A1 => B(25), A2 => n74, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U97 : AOI22_X1 port map( A1 => D(25), A2 => n83, B1 => C(25), B2 => n79, ZN 
                           => n35);
   U98 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(26));
   U99 : AOI22_X1 port map( A1 => B(26), A2 => n74, B1 => A(26), B2 => n70, ZN 
                           => n32);
   U100 : AOI22_X1 port map( A1 => D(26), A2 => n83, B1 => C(26), B2 => n79, ZN
                           => n33);
   U101 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(28));
   U102 : AOI22_X1 port map( A1 => B(28), A2 => n74, B1 => A(28), B2 => n70, ZN
                           => n28);
   U103 : AOI22_X1 port map( A1 => D(28), A2 => n83, B1 => C(28), B2 => n79, ZN
                           => n29);
   U104 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(29));
   U105 : AOI22_X1 port map( A1 => B(29), A2 => n74, B1 => A(29), B2 => n70, ZN
                           => n26);
   U106 : AOI22_X1 port map( A1 => D(29), A2 => n83, B1 => C(29), B2 => n79, ZN
                           => n27);
   U107 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(30));
   U108 : AOI22_X1 port map( A1 => B(30), A2 => n74, B1 => A(30), B2 => n70, ZN
                           => n22);
   U109 : AOI22_X1 port map( A1 => D(30), A2 => n83, B1 => C(30), B2 => n79, ZN
                           => n23);
   U110 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(31));
   U111 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n71, ZN
                           => n20);
   U112 : AOI22_X1 port map( A1 => D(31), A2 => n84, B1 => C(31), B2 => n80, ZN
                           => n21);
   U113 : NOR2_X1 port map( A1 => n85, A2 => SEL(1), ZN => n6);
   U114 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => n7);
   U115 : INV_X1 port map( A => SEL(0), ZN => n85);
   U116 : AND2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n4);
   U117 : AND2_X1 port map( A1 => SEL(1), A2 => n85, ZN => n5);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT2 is

   port( A, B, C, SEL : in std_logic_vector (1 downto 0);  Y : out 
         std_logic_vector (1 downto 0));

end MUX3to1_NBIT2;

architecture SYN_Behavioral of MUX3to1_NBIT2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, N13, N14, n2, n3, n4, n5, n1 : std_logic;

begin
   
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => N14, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => N13, Q => Y(0));
   U9 : NAND3_X1 port map( A1 => C(1), A2 => n1, A3 => SEL(1), ZN => n3);
   U10 : NAND3_X1 port map( A1 => SEL(1), A2 => n1, A3 => C(0), ZN => n5);
   U3 : INV_X1 port map( A => SEL(0), ZN => n1);
   U4 : NAND2_X1 port map( A1 => SEL(0), A2 => SEL(1), ZN => N12);
   U5 : OAI21_X1 port map( B1 => SEL(1), B2 => n4, A => n5, ZN => N13);
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => SEL(0), ZN 
                           => n4);
   U7 : OAI21_X1 port map( B1 => SEL(1), B2 => n2, A => n3, ZN => N14);
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => SEL(0), B2 => B(1), ZN 
                           => n2);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX5to1_NBIT32_0 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX5to1_NBIT32_0;

architecture SYN_Behavioral of MUX5to1_NBIT32_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n1, n2, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
      n94, n95, n96, n97, n98 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n91, D => N57, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n91, D => N56, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n91, D => N55, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n91, D => N54, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n91, D => N53, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n91, D => N52, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n91, D => N51, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n91, D => N50, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n91, D => N49, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n91, D => N48, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n92, D => N47, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n92, D => N46, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n92, D => N45, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n92, D => N44, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n92, D => N43, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n92, D => N42, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n92, D => N41, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n92, D => N40, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n92, D => N39, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n92, D => N38, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n93, D => N37, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n93, D => N36, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n93, D => N35, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n93, D => N34, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n93, D => N33, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n93, D => N32, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n93, D => N31, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n93, D => N30, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n93, D => N29, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n93, D => N28, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n94, D => N27, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n94, D => N26, Q => Y(0));
   U3 : BUF_X1 port map( A => N25, Z => n95);
   U4 : BUF_X1 port map( A => n7, Z => n82);
   U5 : BUF_X1 port map( A => n5, Z => n90);
   U6 : BUF_X1 port map( A => n8, Z => n78);
   U7 : BUF_X1 port map( A => n9, Z => n74);
   U8 : BUF_X1 port map( A => n6, Z => n83);
   U9 : BUF_X1 port map( A => n95, Z => n93);
   U10 : BUF_X1 port map( A => n95, Z => n92);
   U11 : BUF_X1 port map( A => n95, Z => n94);
   U12 : BUF_X1 port map( A => n96, Z => n91);
   U13 : BUF_X1 port map( A => N25, Z => n96);
   U14 : OR4_X1 port map( A1 => n86, A2 => n79, A3 => n72, A4 => n87, ZN => N25
                           );
   U15 : OR2_X1 port map( A1 => n73, A2 => n77, ZN => n72);
   U16 : BUF_X1 port map( A => n90, Z => n87);
   U17 : BUF_X1 port map( A => n90, Z => n88);
   U18 : BUF_X1 port map( A => n78, Z => n76);
   U19 : BUF_X1 port map( A => n78, Z => n75);
   U20 : BUF_X1 port map( A => n74, Z => n2);
   U21 : BUF_X1 port map( A => n74, Z => n1);
   U22 : BUF_X1 port map( A => n83, Z => n85);
   U23 : BUF_X1 port map( A => n83, Z => n84);
   U24 : BUF_X1 port map( A => n82, Z => n79);
   U25 : BUF_X1 port map( A => n82, Z => n80);
   U26 : BUF_X1 port map( A => n83, Z => n86);
   U27 : BUF_X1 port map( A => n82, Z => n81);
   U28 : BUF_X1 port map( A => n78, Z => n77);
   U29 : BUF_X1 port map( A => n74, Z => n73);
   U30 : BUF_X1 port map( A => n90, Z => n89);
   U31 : INV_X1 port map( A => SEL(0), ZN => n97);
   U32 : INV_X1 port map( A => SEL(1), ZN => n98);
   U33 : NOR3_X1 port map( A1 => n97, A2 => SEL(2), A3 => n98, ZN => n7);
   U34 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n98, ZN => n5);
   U35 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n97, ZN => n8);
   U36 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n9);
   U37 : AND3_X1 port map( A1 => n97, A2 => n98, A3 => SEL(2), ZN => n6);
   U38 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N26);
   U39 : AOI22_X1 port map( A1 => B(0), A2 => n77, B1 => A(0), B2 => n73, ZN =>
                           n70);
   U40 : AOI222_X1 port map( A1 => C(0), A2 => n87, B1 => E(0), B2 => n86, C1 
                           => D(0), C2 => n79, ZN => n71);
   U41 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N27);
   U42 : AOI22_X1 port map( A1 => B(1), A2 => n77, B1 => A(1), B2 => n73, ZN =>
                           n68);
   U43 : AOI222_X1 port map( A1 => C(1), A2 => n87, B1 => E(1), B2 => n86, C1 
                           => D(1), C2 => n79, ZN => n69);
   U44 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N28);
   U45 : AOI22_X1 port map( A1 => B(2), A2 => n77, B1 => A(2), B2 => n73, ZN =>
                           n66);
   U46 : AOI222_X1 port map( A1 => C(2), A2 => n87, B1 => E(2), B2 => n86, C1 
                           => D(2), C2 => n79, ZN => n67);
   U47 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N29);
   U48 : AOI22_X1 port map( A1 => B(3), A2 => n77, B1 => A(3), B2 => n73, ZN =>
                           n64);
   U49 : AOI222_X1 port map( A1 => C(3), A2 => n87, B1 => E(3), B2 => n86, C1 
                           => D(3), C2 => n79, ZN => n65);
   U50 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N30);
   U51 : AOI22_X1 port map( A1 => B(4), A2 => n77, B1 => A(4), B2 => n73, ZN =>
                           n62);
   U52 : AOI222_X1 port map( A1 => C(4), A2 => n87, B1 => E(4), B2 => n86, C1 
                           => D(4), C2 => n79, ZN => n63);
   U53 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N31);
   U54 : AOI22_X1 port map( A1 => B(5), A2 => n77, B1 => A(5), B2 => n73, ZN =>
                           n60);
   U55 : AOI222_X1 port map( A1 => C(5), A2 => n87, B1 => E(5), B2 => n86, C1 
                           => D(5), C2 => n79, ZN => n61);
   U56 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N32);
   U57 : AOI22_X1 port map( A1 => B(6), A2 => n77, B1 => A(6), B2 => n73, ZN =>
                           n58);
   U58 : AOI222_X1 port map( A1 => C(6), A2 => n87, B1 => E(6), B2 => n86, C1 
                           => D(6), C2 => n79, ZN => n59);
   U59 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => N33);
   U60 : AOI22_X1 port map( A1 => B(7), A2 => n77, B1 => A(7), B2 => n73, ZN =>
                           n56_port);
   U61 : AOI222_X1 port map( A1 => C(7), A2 => n87, B1 => E(7), B2 => n86, C1 
                           => D(7), C2 => n79, ZN => n57_port);
   U62 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => N34);
   U63 : AOI22_X1 port map( A1 => B(8), A2 => n76, B1 => A(8), B2 => n2, ZN => 
                           n54_port);
   U64 : AOI222_X1 port map( A1 => C(8), A2 => n87, B1 => E(8), B2 => n85, C1 
                           => D(8), C2 => n79, ZN => n55_port);
   U65 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => N35);
   U66 : AOI22_X1 port map( A1 => B(9), A2 => n76, B1 => A(9), B2 => n2, ZN => 
                           n52_port);
   U67 : AOI222_X1 port map( A1 => C(9), A2 => n87, B1 => E(9), B2 => n85, C1 
                           => D(9), C2 => n79, ZN => n53_port);
   U68 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => N36);
   U69 : AOI22_X1 port map( A1 => B(10), A2 => n76, B1 => A(10), B2 => n2, ZN 
                           => n50_port);
   U70 : AOI222_X1 port map( A1 => C(10), A2 => n87, B1 => E(10), B2 => n85, C1
                           => D(10), C2 => n79, ZN => n51_port);
   U71 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => N37);
   U72 : AOI22_X1 port map( A1 => B(11), A2 => n76, B1 => A(11), B2 => n2, ZN 
                           => n48_port);
   U73 : AOI222_X1 port map( A1 => C(11), A2 => n87, B1 => E(11), B2 => n85, C1
                           => D(11), C2 => n80, ZN => n49_port);
   U74 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => N38);
   U75 : AOI22_X1 port map( A1 => B(12), A2 => n76, B1 => A(12), B2 => n2, ZN 
                           => n46_port);
   U76 : AOI222_X1 port map( A1 => C(12), A2 => n88, B1 => E(12), B2 => n85, C1
                           => D(12), C2 => n80, ZN => n47_port);
   U77 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => N39);
   U78 : AOI22_X1 port map( A1 => B(13), A2 => n76, B1 => A(13), B2 => n2, ZN 
                           => n44_port);
   U79 : AOI222_X1 port map( A1 => C(13), A2 => n88, B1 => E(13), B2 => n85, C1
                           => D(13), C2 => n80, ZN => n45_port);
   U80 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => N40);
   U81 : AOI22_X1 port map( A1 => B(14), A2 => n76, B1 => A(14), B2 => n2, ZN 
                           => n42_port);
   U82 : AOI222_X1 port map( A1 => C(14), A2 => n88, B1 => E(14), B2 => n85, C1
                           => D(14), C2 => n80, ZN => n43_port);
   U83 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => N41);
   U84 : AOI22_X1 port map( A1 => B(15), A2 => n76, B1 => A(15), B2 => n2, ZN 
                           => n40_port);
   U85 : AOI222_X1 port map( A1 => C(15), A2 => n88, B1 => E(15), B2 => n85, C1
                           => D(15), C2 => n80, ZN => n41_port);
   U86 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => N42);
   U87 : AOI22_X1 port map( A1 => B(16), A2 => n76, B1 => A(16), B2 => n2, ZN 
                           => n38_port);
   U88 : AOI222_X1 port map( A1 => C(16), A2 => n88, B1 => E(16), B2 => n85, C1
                           => D(16), C2 => n80, ZN => n39_port);
   U89 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => N43);
   U90 : AOI22_X1 port map( A1 => B(17), A2 => n76, B1 => A(17), B2 => n2, ZN 
                           => n36_port);
   U91 : AOI222_X1 port map( A1 => C(17), A2 => n88, B1 => E(17), B2 => n85, C1
                           => D(17), C2 => n80, ZN => n37_port);
   U92 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => N44);
   U93 : AOI22_X1 port map( A1 => B(18), A2 => n76, B1 => A(18), B2 => n2, ZN 
                           => n34_port);
   U94 : AOI222_X1 port map( A1 => C(18), A2 => n88, B1 => E(18), B2 => n85, C1
                           => D(18), C2 => n80, ZN => n35_port);
   U95 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => N45);
   U96 : AOI22_X1 port map( A1 => B(19), A2 => n76, B1 => A(19), B2 => n2, ZN 
                           => n32_port);
   U97 : AOI222_X1 port map( A1 => C(19), A2 => n88, B1 => E(19), B2 => n85, C1
                           => D(19), C2 => n80, ZN => n33_port);
   U98 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => N46);
   U99 : AOI22_X1 port map( A1 => B(20), A2 => n75, B1 => A(20), B2 => n1, ZN 
                           => n30_port);
   U100 : AOI222_X1 port map( A1 => C(20), A2 => n88, B1 => E(20), B2 => n84, 
                           C1 => D(20), C2 => n80, ZN => n31_port);
   U101 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => N47);
   U102 : AOI22_X1 port map( A1 => B(21), A2 => n75, B1 => A(21), B2 => n1, ZN 
                           => n28_port);
   U103 : AOI222_X1 port map( A1 => C(21), A2 => n88, B1 => E(21), B2 => n84, 
                           C1 => D(21), C2 => n80, ZN => n29_port);
   U104 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => N48);
   U105 : AOI22_X1 port map( A1 => B(22), A2 => n75, B1 => A(22), B2 => n1, ZN 
                           => n26_port);
   U106 : AOI222_X1 port map( A1 => C(22), A2 => n88, B1 => E(22), B2 => n84, 
                           C1 => D(22), C2 => n80, ZN => n27_port);
   U107 : NAND2_X1 port map( A1 => n24, A2 => n25_port, ZN => N49);
   U108 : AOI22_X1 port map( A1 => B(23), A2 => n75, B1 => A(23), B2 => n1, ZN 
                           => n24);
   U109 : AOI222_X1 port map( A1 => C(23), A2 => n88, B1 => E(23), B2 => n84, 
                           C1 => D(23), C2 => n81, ZN => n25_port);
   U110 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => N50);
   U111 : AOI22_X1 port map( A1 => B(24), A2 => n75, B1 => A(24), B2 => n1, ZN 
                           => n22);
   U112 : AOI222_X1 port map( A1 => C(24), A2 => n88, B1 => E(24), B2 => n84, 
                           C1 => D(24), C2 => n81, ZN => n23);
   U113 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => N51);
   U114 : AOI22_X1 port map( A1 => B(25), A2 => n75, B1 => A(25), B2 => n1, ZN 
                           => n20);
   U115 : AOI222_X1 port map( A1 => C(25), A2 => n89, B1 => E(25), B2 => n84, 
                           C1 => D(25), C2 => n81, ZN => n21);
   U116 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => N52);
   U117 : AOI22_X1 port map( A1 => B(26), A2 => n75, B1 => A(26), B2 => n1, ZN 
                           => n18);
   U118 : AOI222_X1 port map( A1 => C(26), A2 => n89, B1 => E(26), B2 => n84, 
                           C1 => D(26), C2 => n81, ZN => n19);
   U119 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => N53);
   U120 : AOI22_X1 port map( A1 => B(27), A2 => n75, B1 => A(27), B2 => n1, ZN 
                           => n16);
   U121 : AOI222_X1 port map( A1 => C(27), A2 => n89, B1 => E(27), B2 => n84, 
                           C1 => D(27), C2 => n81, ZN => n17);
   U122 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => N54);
   U123 : AOI22_X1 port map( A1 => B(28), A2 => n75, B1 => A(28), B2 => n1, ZN 
                           => n14);
   U124 : AOI222_X1 port map( A1 => C(28), A2 => n89, B1 => E(28), B2 => n84, 
                           C1 => D(28), C2 => n81, ZN => n15);
   U125 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => N55);
   U126 : AOI22_X1 port map( A1 => B(29), A2 => n75, B1 => A(29), B2 => n1, ZN 
                           => n12);
   U127 : AOI222_X1 port map( A1 => C(29), A2 => n89, B1 => E(29), B2 => n84, 
                           C1 => D(29), C2 => n81, ZN => n13);
   U128 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => N56);
   U129 : AOI22_X1 port map( A1 => B(30), A2 => n75, B1 => A(30), B2 => n1, ZN 
                           => n10);
   U130 : AOI222_X1 port map( A1 => C(30), A2 => n89, B1 => E(30), B2 => n84, 
                           C1 => D(30), C2 => n81, ZN => n11);
   U131 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N57);
   U132 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n1, ZN 
                           => n3);
   U133 : AOI222_X1 port map( A1 => C(31), A2 => n89, B1 => E(31), B2 => n84, 
                           C1 => D(31), C2 => n81, ZN => n4);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX2to1_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX2to1_NBIT32_0;

architecture SYN_BEHAVIORAL of MUX2to1_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : BUF_X2 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U5 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U6 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U8 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U9 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U11 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U12 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U13 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U14 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U15 : MUX2_X1 port map( A => A(11), B => B(11), S => n2, Z => Y(11));
   U16 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U17 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U20 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U21 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U22 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U23 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U24 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U26 : MUX2_X1 port map( A => A(22), B => B(22), S => n3, Z => Y(22));
   U27 : MUX2_X1 port map( A => A(23), B => B(23), S => n3, Z => Y(23));
   U28 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U29 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U30 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U31 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U32 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U33 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U34 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U35 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX3to1_NBIT32_0 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX3to1_NBIT32_0;

architecture SYN_Behavioral of MUX3to1_NBIT32_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N12, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12_port, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
      , n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n69, n70, n71 : 
      std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => N12, D => n4, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => N12, D => n5, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => N12, D => n6, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => N12, D => n7, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => N12, D => n8, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => N12, D => n9, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => N12, D => n10, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => N12, D => n11, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => N12, D => n12_port, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => N12, D => n13, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => N12, D => n14, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => N12, D => n15, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => N12, D => n16, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => N12, D => n17, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => N12, D => n18, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => N12, D => n19, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => N12, D => n20, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => N12, D => n21, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => N12, D => n22, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => N12, D => n23, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => N12, D => n24, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => N12, D => n25, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => N12, D => n26, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => N12, D => n27, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => N12, D => n28, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => N12, D => n29, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => N12, D => n30, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => N12, D => n31, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => N12, D => n32, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => N12, D => n33, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => N12, D => n69, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => N12, D => n70, Q => Y(0));
   U3 : NOR2_X2 port map( A1 => SEL(0), A2 => SEL(1), ZN => n35);
   U4 : AND2_X2 port map( A1 => SEL(0), A2 => n71, ZN => n37);
   U5 : NOR2_X2 port map( A1 => n71, A2 => SEL(0), ZN => n36);
   U6 : OR3_X1 port map( A1 => n37, A2 => n2, A3 => n1, ZN => N12);
   U7 : BUF_X1 port map( A => n36, Z => n1);
   U8 : BUF_X1 port map( A => n35, Z => n2);
   U9 : BUF_X1 port map( A => n35, Z => n3);
   U10 : INV_X1 port map( A => SEL(1), ZN => n71);
   U11 : INV_X1 port map( A => n68, ZN => n70);
   U12 : AOI222_X1 port map( A1 => A(0), A2 => n2, B1 => C(0), B2 => n1, C1 => 
                           B(0), C2 => n37, ZN => n68);
   U13 : INV_X1 port map( A => n67, ZN => n69);
   U14 : AOI222_X1 port map( A1 => A(1), A2 => n2, B1 => C(1), B2 => n1, C1 => 
                           B(1), C2 => n37, ZN => n67);
   U15 : INV_X1 port map( A => n66, ZN => n33);
   U16 : AOI222_X1 port map( A1 => A(2), A2 => n2, B1 => C(2), B2 => n1, C1 => 
                           B(2), C2 => n37, ZN => n66);
   U17 : INV_X1 port map( A => n65, ZN => n32);
   U18 : AOI222_X1 port map( A1 => A(3), A2 => n2, B1 => C(3), B2 => n1, C1 => 
                           B(3), C2 => n37, ZN => n65);
   U19 : INV_X1 port map( A => n64, ZN => n31);
   U20 : AOI222_X1 port map( A1 => A(4), A2 => n2, B1 => C(4), B2 => n1, C1 => 
                           B(4), C2 => n37, ZN => n64);
   U21 : INV_X1 port map( A => n63, ZN => n30);
   U22 : AOI222_X1 port map( A1 => A(5), A2 => n2, B1 => C(5), B2 => n1, C1 => 
                           B(5), C2 => n37, ZN => n63);
   U23 : INV_X1 port map( A => n62, ZN => n29);
   U24 : AOI222_X1 port map( A1 => A(6), A2 => n2, B1 => C(6), B2 => n1, C1 => 
                           B(6), C2 => n37, ZN => n62);
   U25 : INV_X1 port map( A => n61, ZN => n28);
   U26 : AOI222_X1 port map( A1 => A(7), A2 => n2, B1 => C(7), B2 => n1, C1 => 
                           B(7), C2 => n37, ZN => n61);
   U27 : INV_X1 port map( A => n60, ZN => n27);
   U28 : AOI222_X1 port map( A1 => A(8), A2 => n2, B1 => C(8), B2 => n36, C1 =>
                           B(8), C2 => n37, ZN => n60);
   U29 : INV_X1 port map( A => n59, ZN => n26);
   U30 : AOI222_X1 port map( A1 => A(9), A2 => n2, B1 => C(9), B2 => n36, C1 =>
                           B(9), C2 => n37, ZN => n59);
   U31 : INV_X1 port map( A => n58, ZN => n25);
   U32 : AOI222_X1 port map( A1 => A(10), A2 => n2, B1 => C(10), B2 => n36, C1 
                           => B(10), C2 => n37, ZN => n58);
   U33 : INV_X1 port map( A => n57, ZN => n24);
   U34 : AOI222_X1 port map( A1 => A(11), A2 => n35, B1 => C(11), B2 => n36, C1
                           => B(11), C2 => n37, ZN => n57);
   U35 : INV_X1 port map( A => n56, ZN => n23);
   U36 : AOI222_X1 port map( A1 => A(12), A2 => n35, B1 => C(12), B2 => n36, C1
                           => B(12), C2 => n37, ZN => n56);
   U37 : INV_X1 port map( A => n55, ZN => n22);
   U38 : AOI222_X1 port map( A1 => A(13), A2 => n35, B1 => C(13), B2 => n36, C1
                           => B(13), C2 => n37, ZN => n55);
   U39 : INV_X1 port map( A => n54, ZN => n21);
   U40 : AOI222_X1 port map( A1 => A(14), A2 => n35, B1 => C(14), B2 => n36, C1
                           => B(14), C2 => n37, ZN => n54);
   U41 : INV_X1 port map( A => n53, ZN => n20);
   U42 : AOI222_X1 port map( A1 => A(15), A2 => n35, B1 => C(15), B2 => n36, C1
                           => B(15), C2 => n37, ZN => n53);
   U43 : INV_X1 port map( A => n52, ZN => n19);
   U44 : AOI222_X1 port map( A1 => A(16), A2 => n35, B1 => C(16), B2 => n36, C1
                           => B(16), C2 => n37, ZN => n52);
   U45 : INV_X1 port map( A => n51, ZN => n18);
   U46 : AOI222_X1 port map( A1 => A(17), A2 => n35, B1 => C(17), B2 => n36, C1
                           => B(17), C2 => n37, ZN => n51);
   U47 : INV_X1 port map( A => n50, ZN => n17);
   U48 : AOI222_X1 port map( A1 => A(18), A2 => n35, B1 => C(18), B2 => n36, C1
                           => B(18), C2 => n37, ZN => n50);
   U49 : INV_X1 port map( A => n49, ZN => n16);
   U50 : AOI222_X1 port map( A1 => A(19), A2 => n35, B1 => C(19), B2 => n36, C1
                           => B(19), C2 => n37, ZN => n49);
   U51 : INV_X1 port map( A => n48, ZN => n15);
   U52 : AOI222_X1 port map( A1 => A(20), A2 => n35, B1 => C(20), B2 => n1, C1 
                           => B(20), C2 => n37, ZN => n48);
   U53 : INV_X1 port map( A => n47, ZN => n14);
   U54 : AOI222_X1 port map( A1 => A(21), A2 => n35, B1 => C(21), B2 => n1, C1 
                           => B(21), C2 => n37, ZN => n47);
   U55 : INV_X1 port map( A => n46, ZN => n13);
   U56 : AOI222_X1 port map( A1 => A(22), A2 => n35, B1 => C(22), B2 => n1, C1 
                           => B(22), C2 => n37, ZN => n46);
   U57 : INV_X1 port map( A => n45, ZN => n12_port);
   U58 : AOI222_X1 port map( A1 => A(23), A2 => n3, B1 => C(23), B2 => n1, C1 
                           => B(23), C2 => n37, ZN => n45);
   U59 : INV_X1 port map( A => n44, ZN => n11);
   U60 : AOI222_X1 port map( A1 => A(24), A2 => n3, B1 => C(24), B2 => n1, C1 
                           => B(24), C2 => n37, ZN => n44);
   U61 : INV_X1 port map( A => n43, ZN => n10);
   U62 : AOI222_X1 port map( A1 => A(25), A2 => n3, B1 => C(25), B2 => n1, C1 
                           => B(25), C2 => n37, ZN => n43);
   U63 : INV_X1 port map( A => n42, ZN => n9);
   U64 : AOI222_X1 port map( A1 => A(26), A2 => n3, B1 => C(26), B2 => n1, C1 
                           => B(26), C2 => n37, ZN => n42);
   U65 : INV_X1 port map( A => n41, ZN => n8);
   U66 : AOI222_X1 port map( A1 => A(27), A2 => n3, B1 => C(27), B2 => n1, C1 
                           => B(27), C2 => n37, ZN => n41);
   U67 : INV_X1 port map( A => n40, ZN => n7);
   U68 : AOI222_X1 port map( A1 => A(28), A2 => n3, B1 => C(28), B2 => n1, C1 
                           => B(28), C2 => n37, ZN => n40);
   U69 : INV_X1 port map( A => n39, ZN => n6);
   U70 : AOI222_X1 port map( A1 => A(29), A2 => n3, B1 => C(29), B2 => n1, C1 
                           => B(29), C2 => n37, ZN => n39);
   U71 : INV_X1 port map( A => n38, ZN => n5);
   U72 : AOI222_X1 port map( A1 => A(30), A2 => n3, B1 => C(30), B2 => n1, C1 
                           => B(30), C2 => n37, ZN => n38);
   U73 : INV_X1 port map( A => n34, ZN => n4);
   U74 : AOI222_X1 port map( A1 => A(31), A2 => n3, B1 => C(31), B2 => n1, C1 
                           => B(31), C2 => n37, ZN => n34);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PC_adder_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Sum : out std_logic_vector 
         (31 downto 0));

end PC_adder_0;

architecture SYN_Behavioral of PC_adder_0 is

   component PC_adder_0_DW01_add_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1623 : std_logic;

begin
   
   n1 <= '0';
   add_16 : PC_adder_0_DW01_add_2 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(31) => Sum(31), 
                           SUM(30) => Sum(30), SUM(29) => Sum(29), SUM(28) => 
                           Sum(28), SUM(27) => Sum(27), SUM(26) => Sum(26), 
                           SUM(25) => Sum(25), SUM(24) => Sum(24), SUM(23) => 
                           Sum(23), SUM(22) => Sum(22), SUM(21) => Sum(21), 
                           SUM(20) => Sum(20), SUM(19) => Sum(19), SUM(18) => 
                           Sum(18), SUM(17) => Sum(17), SUM(16) => Sum(16), 
                           SUM(15) => Sum(15), SUM(14) => Sum(14), SUM(13) => 
                           Sum(13), SUM(12) => Sum(12), SUM(11) => Sum(11), 
                           SUM(10) => Sum(10), SUM(9) => Sum(9), SUM(8) => 
                           Sum(8), SUM(7) => Sum(7), SUM(6) => Sum(6), SUM(5) 
                           => Sum(5), SUM(4) => Sum(4), SUM(3) => Sum(3), 
                           SUM(2) => Sum(2), SUM(1) => Sum(1), SUM(0) => Sum(0)
                           , CO => n_1623);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT7 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (6 
         downto 0);  data_out : out std_logic_vector (6 downto 0));

end REG_NBIT7;

architecture SYN_Behavioral of REG_NBIT7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n22, n21, n23, n24, n25 : std_logic;

begin
   
   reg_reg_6_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n25, Q => 
                           data_out(6), QN => n14);
   reg_reg_5_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n25, Q => 
                           data_out(5), QN => n13);
   reg_reg_4_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n25, Q => 
                           data_out(4), QN => n12);
   reg_reg_3_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n25, Q => 
                           data_out(3), QN => n11);
   reg_reg_2_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n25, Q => 
                           data_out(2), QN => n10);
   reg_reg_1_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n25, Q => 
                           data_out(1), QN => n9);
   reg_reg_0_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n25, Q => 
                           data_out(0), QN => n8);
   U2 : INV_X1 port map( A => reset, ZN => n25);
   U3 : BUF_X1 port map( A => n24, Z => n21);
   U4 : BUF_X1 port map( A => n24, Z => n23);
   U5 : BUF_X1 port map( A => enable, Z => n24);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n21, A => n3, ZN => n17);
   U7 : NAND2_X1 port map( A1 => data_in(2), A2 => n21, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n8, B2 => n21, A => n1, ZN => n15);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n21, A => n2, ZN => n16);
   U10 : OAI21_X1 port map( B1 => n12, B2 => n21, A => n5, ZN => n19);
   U11 : OAI21_X1 port map( B1 => n13, B2 => n23, A => n6, ZN => n20);
   U12 : OAI21_X1 port map( B1 => n14, B2 => n21, A => n7, ZN => n22);
   U13 : NAND2_X1 port map( A1 => data_in(6), A2 => n21, ZN => n7);
   U14 : NAND2_X1 port map( A1 => data_in(3), A2 => n21, ZN => n4);
   U15 : NAND2_X1 port map( A1 => data_in(1), A2 => n21, ZN => n2);
   U16 : OAI21_X1 port map( B1 => n11, B2 => n21, A => n4, ZN => n18);
   U17 : NAND2_X1 port map( A1 => data_in(5), A2 => n21, ZN => n6);
   U18 : NAND2_X1 port map( A1 => data_in(4), A2 => n21, ZN => n5);
   U19 : NAND2_X1 port map( A1 => n23, A2 => data_in(0), ZN => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FFD_0;

architecture SYN_BEHAVIORAL of FFD_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2, n4, n1, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n1, Q => Q, QN => n2);
   U2 : INV_X1 port map( A => RESET, ZN => n1);
   U3 : INV_X1 port map( A => n2, ZN => n3);
   U4 : MUX2_X1 port map( A => n3, B => D, S => ENABLE, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_NBIT32_0 is

   port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector (31 
         downto 0);  data_out : out std_logic_vector (31 downto 0));

end REG_NBIT32_0;

architecture SYN_Behavioral of REG_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_27_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n97, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, data_out_16_port, data_out_17_port, 
      data_out_18_port, data_out_19_port, data_out_20_port, data_out_21_port, 
      data_out_22_port, data_out_23_port, data_out_24_port, data_out_25_port, 
      data_out_26_port, data_out_28_port, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639 : std_logic;

begin
   data_out <= ( data_out_31_port, data_out_30_port, data_out_29_port, 
      data_out_28_port, data_out_27_port, data_out_26_port, data_out_25_port, 
      data_out_24_port, data_out_23_port, data_out_22_port, data_out_21_port, 
      data_out_20_port, data_out_19_port, data_out_18_port, data_out_17_port, 
      data_out_16_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   reg_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n25, Q => 
                           data_out_31_port, QN => n_1624);
   reg_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n25, Q => 
                           data_out_30_port, QN => n_1625);
   reg_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n25, Q => 
                           data_out_29_port, QN => n_1626);
   reg_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n25, Q => 
                           data_out_28_port, QN => n_1627);
   reg_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n25, Q => 
                           data_out_26_port, QN => n_1628);
   reg_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n26, Q => 
                           data_out_25_port, QN => n_1629);
   reg_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n26, Q => 
                           data_out_24_port, QN => n_1630);
   reg_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n26, Q => 
                           data_out_23_port, QN => n_1631);
   reg_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n26, Q => 
                           data_out_22_port, QN => n_1632);
   reg_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n26, Q => 
                           data_out_21_port, QN => n_1633);
   reg_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n26, Q => 
                           data_out_20_port, QN => n_1634);
   reg_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n26, Q => 
                           data_out_19_port, QN => n_1635);
   reg_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n26, Q => 
                           data_out_18_port, QN => n_1636);
   reg_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n26, Q => 
                           data_out_17_port, QN => n_1637);
   reg_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n26, Q => 
                           data_out_16_port, QN => n_1638);
   reg_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n24, Q => 
                           data_out_15_port, QN => n48);
   reg_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n24, Q => 
                           data_out_14_port, QN => n47);
   reg_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n24, Q => 
                           data_out_13_port, QN => n46);
   reg_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n24, Q => 
                           data_out_12_port, QN => n45);
   reg_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n24, Q => 
                           data_out_11_port, QN => n44);
   reg_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n24, Q => 
                           data_out_10_port, QN => n43);
   reg_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n24, Q => 
                           data_out_9_port, QN => n42);
   reg_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n24, Q => 
                           data_out_8_port, QN => n41);
   reg_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n24, Q => 
                           data_out_7_port, QN => n40);
   reg_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n24, Q => 
                           data_out_6_port, QN => n39);
   reg_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n24, Q => 
                           data_out_5_port, QN => n38);
   reg_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n25, Q => 
                           data_out_4_port, QN => n37);
   reg_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n25, Q => 
                           data_out_3_port, QN => n36);
   reg_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n25, Q => 
                           data_out_2_port, QN => n35);
   reg_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n25, Q => 
                           data_out_1_port, QN => n34);
   reg_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n25, Q => 
                           data_out_0_port, QN => n33);
   reg_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n28, Q => 
                           data_out_27_port, QN => n_1639);
   U2 : BUF_X1 port map( A => n17, Z => n22);
   U3 : BUF_X1 port map( A => n28, Z => n27);
   U4 : BUF_X1 port map( A => n22, Z => n19);
   U5 : BUF_X1 port map( A => n22, Z => n20);
   U6 : BUF_X1 port map( A => n22, Z => n21);
   U7 : BUF_X1 port map( A => n27, Z => n24);
   U8 : BUF_X1 port map( A => n27, Z => n25);
   U9 : BUF_X1 port map( A => n27, Z => n26);
   U10 : BUF_X1 port map( A => n23, Z => n18);
   U11 : BUF_X1 port map( A => n17, Z => n23);
   U12 : INV_X1 port map( A => reset, ZN => n28);
   U13 : BUF_X1 port map( A => enable, Z => n17);
   U14 : OAI21_X1 port map( B1 => n34, B2 => n19, A => n2, ZN => n66);
   U15 : NAND2_X1 port map( A1 => data_in(1), A2 => n19, ZN => n2);
   U16 : OAI21_X1 port map( B1 => n35, B2 => n19, A => n3, ZN => n67);
   U17 : NAND2_X1 port map( A1 => data_in(2), A2 => n19, ZN => n3);
   U18 : OAI21_X1 port map( B1 => n36, B2 => n19, A => n4, ZN => n68);
   U19 : NAND2_X1 port map( A1 => data_in(3), A2 => n19, ZN => n4);
   U20 : OAI21_X1 port map( B1 => n33, B2 => n19, A => n1, ZN => n65);
   U21 : NAND2_X1 port map( A1 => n20, A2 => data_in(0), ZN => n1);
   U22 : OAI21_X1 port map( B1 => n48, B2 => n20, A => n16, ZN => n80);
   U23 : NAND2_X1 port map( A1 => data_in(15), A2 => n18, ZN => n16);
   U24 : OAI21_X1 port map( B1 => n42, B2 => n20, A => n10, ZN => n74);
   U25 : NAND2_X1 port map( A1 => data_in(9), A2 => n18, ZN => n10);
   U26 : OAI21_X1 port map( B1 => n43, B2 => n20, A => n11, ZN => n75);
   U27 : NAND2_X1 port map( A1 => data_in(10), A2 => n18, ZN => n11);
   U28 : OAI21_X1 port map( B1 => n44, B2 => n20, A => n12, ZN => n76);
   U29 : NAND2_X1 port map( A1 => data_in(11), A2 => n18, ZN => n12);
   U30 : OAI21_X1 port map( B1 => n45, B2 => n20, A => n13, ZN => n77);
   U31 : NAND2_X1 port map( A1 => data_in(12), A2 => n18, ZN => n13);
   U32 : OAI21_X1 port map( B1 => n46, B2 => n20, A => n14, ZN => n78);
   U33 : NAND2_X1 port map( A1 => data_in(13), A2 => n18, ZN => n14);
   U34 : OAI21_X1 port map( B1 => n47, B2 => n20, A => n15, ZN => n79);
   U35 : NAND2_X1 port map( A1 => data_in(14), A2 => n18, ZN => n15);
   U36 : OAI21_X1 port map( B1 => n37, B2 => n19, A => n5, ZN => n69);
   U37 : NAND2_X1 port map( A1 => data_in(4), A2 => n18, ZN => n5);
   U38 : OAI21_X1 port map( B1 => n38, B2 => n19, A => n6, ZN => n70);
   U39 : NAND2_X1 port map( A1 => data_in(5), A2 => n18, ZN => n6);
   U40 : OAI21_X1 port map( B1 => n39, B2 => n19, A => n7, ZN => n71);
   U41 : NAND2_X1 port map( A1 => data_in(6), A2 => n18, ZN => n7);
   U42 : OAI21_X1 port map( B1 => n40, B2 => n19, A => n8, ZN => n72);
   U43 : NAND2_X1 port map( A1 => data_in(7), A2 => n18, ZN => n8);
   U44 : OAI21_X1 port map( B1 => n41, B2 => n19, A => n9, ZN => n73);
   U45 : NAND2_X1 port map( A1 => data_in(8), A2 => n18, ZN => n9);
   U46 : MUX2_X1 port map( A => data_out_16_port, B => data_in(16), S => n21, Z
                           => n81);
   U47 : MUX2_X1 port map( A => data_out_17_port, B => data_in(17), S => n21, Z
                           => n82);
   U48 : MUX2_X1 port map( A => data_out_18_port, B => data_in(18), S => n21, Z
                           => n83);
   U49 : MUX2_X1 port map( A => data_out_19_port, B => data_in(19), S => n21, Z
                           => n84);
   U50 : MUX2_X1 port map( A => data_out_20_port, B => data_in(20), S => n21, Z
                           => n85);
   U51 : MUX2_X1 port map( A => data_out_21_port, B => data_in(21), S => n21, Z
                           => n86);
   U52 : MUX2_X1 port map( A => data_out_22_port, B => data_in(22), S => n21, Z
                           => n87);
   U53 : MUX2_X1 port map( A => data_out_23_port, B => data_in(23), S => n21, Z
                           => n88);
   U54 : MUX2_X1 port map( A => data_out_24_port, B => data_in(24), S => n21, Z
                           => n89);
   U55 : MUX2_X1 port map( A => data_out_25_port, B => data_in(25), S => n21, Z
                           => n90);
   U56 : MUX2_X1 port map( A => data_out_26_port, B => data_in(26), S => n20, Z
                           => n91);
   U57 : MUX2_X1 port map( A => data_out_27_port, B => data_in(27), S => n20, Z
                           => n92);
   U58 : MUX2_X1 port map( A => data_out_28_port, B => data_in(28), S => n20, Z
                           => n93);
   U59 : MUX2_X1 port map( A => data_out_29_port, B => data_in(29), S => n20, Z
                           => n94);
   U60 : MUX2_X1 port map( A => data_out_30_port, B => data_in(30), S => n20, Z
                           => n95);
   U61 : MUX2_X1 port map( A => data_out_31_port, B => data_in(31), S => n20, Z
                           => n97);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector (31 
         downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out std_logic_vector (31 
         downto 0);  BMP : inout std_logic;  STALL : out std_logic_vector (1 
         downto 0);  ID_EN, RF_RD, SIGND, IMM_SEL, BPR_EN : in std_logic;  
         ALU_OPCODE : in std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, ALUB_SEL,
         UCB_EN, MEM_EN, MEM_DATA_SEL : in std_logic;  LD_SEL : in 
         std_logic_vector (2 downto 0);  ALR2_SEL : in std_logic;  CWB_SEL : in
         std_logic_vector (1 downto 0);  WB_SEL, RF_WR : in std_logic;  
         RF_MUX_SEL : in std_logic_vector (1 downto 0));

end Datapath;

architecture SYN_BEHAVIORAL of Datapath is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RF_NBIT32_NREG32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component CWBU
      port( CLOCK : in std_logic;  ALU_OP : in std_logic_vector (0 to 4);  PSW 
            : in std_logic_vector (6 downto 0);  COND_SEL : out 
            std_logic_vector (1 downto 0);  CWB_SEL : in std_logic_vector (1 
            downto 0);  CWB_MUW_SEL : out std_logic_vector (1 downto 0));
   end component;
   
   component BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0
      port( clock, rst : in std_logic;  address : in std_logic_vector (31 
            downto 0);  d_in, w_en : in std_logic;  d_out : out std_logic);
   end component;
   
   component HDU_IR_SIZE32
      port( clk, rst : in std_logic;  IR : in std_logic_vector (31 downto 0);  
            STALL_CODE : out std_logic_vector (1 downto 0);  IF_STALL, ID_STALL
            , EX_STALL, MEM_STALL, WB_STALL : out std_logic);
   end component;
   
   component FWDU_IR_SIZE32
      port( CLOCK, RESET, EN : in std_logic;  IR : in std_logic_vector (31 
            downto 0);  FWD_A, FWD_B : out std_logic_vector (1 downto 0);  
            FWD_B2 : out std_logic;  ZDU_SEL : out std_logic_vector (1 downto 
            0));
   end component;
   
   component ALU_NBIT32
      port( CLOCK : in std_logic;  AluOpcode : in std_logic_vector (0 to 4);  A
            , B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            ALU_out : out std_logic_vector (31 downto 0);  Cout : out std_logic
            ;  COND : out std_logic_vector (5 downto 0));
   end component;
   
   component MUX3to1_NBIT5
      port( A, B, C : in std_logic_vector (4 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (4 downto 
            0));
   end component;
   
   component MUX2to1_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX4to1_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT2
      port( A, B, C, SEL : in std_logic_vector (1 downto 0);  Y : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component MUX2to1_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX5to1_NBIT32_0
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX2to1_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX3to1_NBIT32_1
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT32_2
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX3to1_NBIT32_3
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX2to1_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_8
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX2to1_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX3to1_NBIT32_0
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component PC_adder_1
      port( A, B : in std_logic_vector (31 downto 0);  Sum : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component PC_adder_0
      port( A, B : in std_logic_vector (31 downto 0);  Sum : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_4
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_5
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT7
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (6 downto 0);  data_out : out std_logic_vector (6 downto 0));
   end component;
   
   component REG_NBIT32_6
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_7
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_8
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_9
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_10
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component FFD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component REG_NBIT32_11
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_12
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component FFD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component REG_NBIT32_13
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_14
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_15
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_16
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_17
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_NBIT32_0
      port( clk, reset, enable : in std_logic;  data_in : in std_logic_vector 
            (31 downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IRAM_ADDR_31_port, IRAM_ADDR_30_port, 
      IRAM_ADDR_29_port, IRAM_ADDR_28_port, IRAM_ADDR_27_port, 
      IRAM_ADDR_26_port, IRAM_ADDR_25_port, IRAM_ADDR_24_port, 
      IRAM_ADDR_23_port, IRAM_ADDR_22_port, IRAM_ADDR_21_port, 
      IRAM_ADDR_20_port, IRAM_ADDR_19_port, IRAM_ADDR_18_port, 
      IRAM_ADDR_17_port, IRAM_ADDR_16_port, IRAM_ADDR_15_port, 
      IRAM_ADDR_14_port, IRAM_ADDR_13_port, IRAM_ADDR_12_port, 
      IRAM_ADDR_11_port, IRAM_ADDR_10_port, IRAM_ADDR_9_port, IRAM_ADDR_8_port,
      IRAM_ADDR_7_port, IRAM_ADDR_6_port, IRAM_ADDR_5_port, IRAM_ADDR_4_port, 
      IRAM_ADDR_3_port, IRAM_ADDR_2_port, IRAM_ADDR_1_port, IRAM_ADDR_0_port, 
      DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port, NPC_in_31_port, 
      NPC_in_30_port, NPC_in_29_port, NPC_in_28_port, NPC_in_27_port, 
      NPC_in_26_port, NPC_in_25_port, NPC_in_24_port, NPC_in_23_port, 
      NPC_in_22_port, NPC_in_21_port, NPC_in_20_port, NPC_in_19_port, 
      NPC_in_18_port, NPC_in_17_port, NPC_in_16_port, NPC_in_15_port, 
      NPC_in_14_port, NPC_in_13_port, NPC_in_12_port, NPC_in_11_port, 
      NPC_in_10_port, NPC_in_9_port, NPC_in_8_port, NPC_in_7_port, 
      NPC_in_6_port, NPC_in_5_port, NPC_in_4_port, NPC_in_3_port, NPC_in_2_port
      , NPC_in_1_port, NPC_in_0_port, PC_out_31_port, PC_out_30_port, 
      PC_out_29_port, PC_out_28_port, PC_out_27_port, PC_out_26_port, 
      PC_out_25_port, PC_out_24_port, PC_out_23_port, PC_out_22_port, 
      PC_out_21_port, PC_out_20_port, PC_out_19_port, PC_out_18_port, 
      PC_out_17_port, PC_out_16_port, PC_out_15_port, PC_out_14_port, 
      PC_out_13_port, PC_out_12_port, PC_out_11_port, PC_out_10_port, 
      PC_out_9_port, PC_out_8_port, PC_out_7_port, PC_out_6_port, PC_out_5_port
      , PC_out_4_port, PC_out_3_port, PC_out_2_port, PC_out_1_port, 
      PC_out_0_port, IR_out_31_port, IR_out_30_port, IR_out_29_port, 
      IR_out_28_port, IR_out_27_port, IR_out_26_port, IR_out_25_port, 
      IR_out_24_port, IR_out_23_port, IR_out_22_port, IR_out_21_port, 
      IR_out_20_port, IR_out_19_port, IR_out_18_port, IR_out_17_port, 
      IR_out_16_port, IR_out_15_port, IR_out_14_port, IR_out_13_port, 
      IR_out_12_port, IR_out_11_port, IR_out_10_port, IR_out_9_port, 
      IR_out_8_port, IR_out_7_port, IR_out_6_port, IR_out_5_port, IR_out_4_port
      , IR_out_3_port, IR_out_2_port, IR_out_1_port, IR_out_0_port, 
      NPC_out_31_port, NPC_out_30_port, NPC_out_29_port, NPC_out_28_port, 
      NPC_out_27_port, NPC_out_26_port, NPC_out_25_port, NPC_out_24_port, 
      NPC_out_23_port, NPC_out_22_port, NPC_out_21_port, NPC_out_20_port, 
      NPC_out_19_port, NPC_out_18_port, NPC_out_17_port, NPC_out_16_port, 
      NPC_out_15_port, NPC_out_14_port, NPC_out_13_port, NPC_out_12_port, 
      NPC_out_11_port, NPC_out_10_port, NPC_out_9_port, NPC_out_8_port, 
      NPC_out_7_port, NPC_out_6_port, NPC_out_5_port, NPC_out_4_port, 
      NPC_out_3_port, NPC_out_2_port, NPC_out_1_port, NPC_out_0_port, ID_ENABLE
      , PC2_out_31_port, PC2_out_30_port, PC2_out_29_port, PC2_out_28_port, 
      PC2_out_27_port, PC2_out_26_port, PC2_out_25_port, PC2_out_24_port, 
      PC2_out_23_port, PC2_out_22_port, PC2_out_21_port, PC2_out_20_port, 
      PC2_out_19_port, PC2_out_18_port, PC2_out_17_port, PC2_out_16_port, 
      PC2_out_15_port, PC2_out_14_port, PC2_out_13_port, PC2_out_12_port, 
      PC2_out_11_port, PC2_out_10_port, PC2_out_9_port, PC2_out_8_port, 
      PC2_out_7_port, PC2_out_6_port, PC2_out_5_port, PC2_out_4_port, 
      PC2_out_3_port, PC2_out_2_port, PC2_out_1_port, PC2_out_0_port, 
      RIMM_out_31_port, RIMM_out_30_port, RIMM_out_29_port, RIMM_out_28_port, 
      RIMM_out_27_port, RIMM_out_26_port, RIMM_out_25_port, RIMM_out_24_port, 
      RIMM_out_23_port, RIMM_out_22_port, RIMM_out_21_port, RIMM_out_20_port, 
      RIMM_out_19_port, RIMM_out_18_port, RIMM_out_17_port, RIMM_out_16_port, 
      RIMM_out_15_port, RIMM_out_14_port, RIMM_out_13_port, RIMM_out_12_port, 
      RIMM_out_11_port, RIMM_out_10_port, RIMM_out_9_port, RIMM_out_8_port, 
      RIMM_out_7_port, RIMM_out_6_port, RIMM_out_5_port, RIMM_out_4_port, 
      RIMM_out_3_port, RIMM_out_2_port, RIMM_out_1_port, RIMM_out_0_port, 
      RWB1_out_31_port, RWB1_out_30_port, RWB1_out_29_port, RWB1_out_28_port, 
      RWB1_out_27_port, RWB1_out_26_port, RWB1_out_25_port, RWB1_out_24_port, 
      RWB1_out_23_port, RWB1_out_22_port, RWB1_out_21_port, RWB1_out_20_port, 
      RWB1_out_19_port, RWB1_out_18_port, RWB1_out_17_port, RWB1_out_16_port, 
      RWB1_out_15_port, RWB1_out_14_port, RWB1_out_13_port, RWB1_out_12_port, 
      RWB1_out_11_port, RWB1_out_10_port, RWB1_out_9_port, RWB1_out_8_port, 
      RWB1_out_7_port, RWB1_out_6_port, RWB1_out_5_port, RWB1_out_4_port, 
      RWB1_out_3_port, RWB1_out_2_port, RWB1_out_1_port, RWB1_out_0_port, 
      BHT_out, PRD_OUT, NPC2_out_31_port, NPC2_out_30_port, NPC2_out_29_port, 
      NPC2_out_28_port, NPC2_out_27_port, NPC2_out_26_port, NPC2_out_25_port, 
      NPC2_out_24_port, NPC2_out_23_port, NPC2_out_22_port, NPC2_out_21_port, 
      NPC2_out_20_port, NPC2_out_19_port, NPC2_out_18_port, NPC2_out_17_port, 
      NPC2_out_16_port, NPC2_out_15_port, NPC2_out_14_port, NPC2_out_13_port, 
      NPC2_out_12_port, NPC2_out_11_port, NPC2_out_10_port, NPC2_out_9_port, 
      NPC2_out_8_port, NPC2_out_7_port, NPC2_out_6_port, NPC2_out_5_port, 
      NPC2_out_4_port, NPC2_out_3_port, NPC2_out_2_port, NPC2_out_1_port, 
      NPC2_out_0_port, JADDER_out_31_port, JADDER_out_30_port, 
      JADDER_out_29_port, JADDER_out_28_port, JADDER_out_27_port, 
      JADDER_out_26_port, JADDER_out_25_port, JADDER_out_24_port, 
      JADDER_out_23_port, JADDER_out_22_port, JADDER_out_21_port, 
      JADDER_out_20_port, JADDER_out_19_port, JADDER_out_18_port, 
      JADDER_out_17_port, JADDER_out_16_port, JADDER_out_15_port, 
      JADDER_out_14_port, JADDER_out_13_port, JADDER_out_12_port, 
      JADDER_out_11_port, JADDER_out_10_port, JADDER_out_9_port, 
      JADDER_out_8_port, JADDER_out_7_port, JADDER_out_6_port, 
      JADDER_out_5_port, JADDER_out_4_port, JADDER_out_3_port, 
      JADDER_out_2_port, JADDER_out_1_port, JADDER_out_0_port, 
      JADDER2_out_31_port, JADDER2_out_30_port, JADDER2_out_29_port, 
      JADDER2_out_28_port, JADDER2_out_27_port, JADDER2_out_26_port, 
      JADDER2_out_25_port, JADDER2_out_24_port, JADDER2_out_23_port, 
      JADDER2_out_22_port, JADDER2_out_21_port, JADDER2_out_20_port, 
      JADDER2_out_19_port, JADDER2_out_18_port, JADDER2_out_17_port, 
      JADDER2_out_16_port, JADDER2_out_15_port, JADDER2_out_14_port, 
      JADDER2_out_13_port, JADDER2_out_12_port, JADDER2_out_11_port, 
      JADDER2_out_10_port, JADDER2_out_9_port, JADDER2_out_8_port, 
      JADDER2_out_7_port, JADDER2_out_6_port, JADDER2_out_5_port, 
      JADDER2_out_4_port, JADDER2_out_3_port, JADDER2_out_2_port, 
      JADDER2_out_1_port, JADDER2_out_0_port, BPR_EN2, EX_ENABLE, 
      PC3_out_31_port, PC3_out_30_port, PC3_out_29_port, PC3_out_28_port, 
      PC3_out_27_port, PC3_out_26_port, PC3_out_25_port, PC3_out_24_port, 
      PC3_out_23_port, PC3_out_22_port, PC3_out_21_port, PC3_out_20_port, 
      PC3_out_19_port, PC3_out_18_port, PC3_out_17_port, PC3_out_16_port, 
      PC3_out_15_port, PC3_out_14_port, PC3_out_13_port, PC3_out_12_port, 
      PC3_out_11_port, PC3_out_10_port, PC3_out_9_port, PC3_out_8_port, 
      PC3_out_7_port, PC3_out_6_port, PC3_out_5_port, PC3_out_4_port, 
      PC3_out_3_port, PC3_out_2_port, PC3_out_1_port, PC3_out_0_port, 
      RWB2_out_31_port, RWB2_out_30_port, RWB2_out_29_port, RWB2_out_28_port, 
      RWB2_out_27_port, RWB2_out_26_port, RWB2_out_25_port, RWB2_out_24_port, 
      RWB2_out_23_port, RWB2_out_22_port, RWB2_out_21_port, RWB2_out_20_port, 
      RWB2_out_19_port, RWB2_out_18_port, RWB2_out_17_port, RWB2_out_16_port, 
      RWB2_out_15_port, RWB2_out_14_port, RWB2_out_13_port, RWB2_out_12_port, 
      RWB2_out_11_port, RWB2_out_10_port, RWB2_out_9_port, RWB2_out_8_port, 
      RWB2_out_7_port, RWB2_out_6_port, RWB2_out_5_port, RWB2_out_4_port, 
      RWB2_out_3_port, RWB2_out_2_port, RWB2_out_1_port, RWB2_out_0_port, 
      RB_out_31_port, RB_out_30_port, RB_out_29_port, RB_out_28_port, 
      RB_out_27_port, RB_out_26_port, RB_out_25_port, RB_out_24_port, 
      RB_out_23_port, RB_out_22_port, RB_out_21_port, RB_out_20_port, 
      RB_out_19_port, RB_out_18_port, RB_out_17_port, RB_out_16_port, 
      RB_out_15_port, RB_out_14_port, RB_out_13_port, RB_out_12_port, 
      RB_out_11_port, RB_out_10_port, RB_out_9_port, RB_out_8_port, 
      RB_out_7_port, RB_out_6_port, RB_out_5_port, RB_out_4_port, RB_out_3_port
      , RB_out_2_port, RB_out_1_port, RB_out_0_port, B2_out_31_port, 
      B2_out_30_port, B2_out_29_port, B2_out_28_port, B2_out_27_port, 
      B2_out_26_port, B2_out_25_port, B2_out_24_port, B2_out_23_port, 
      B2_out_22_port, B2_out_21_port, B2_out_20_port, B2_out_19_port, 
      B2_out_18_port, B2_out_17_port, B2_out_16_port, B2_out_15_port, 
      B2_out_14_port, B2_out_13_port, B2_out_12_port, B2_out_11_port, 
      B2_out_10_port, B2_out_9_port, B2_out_8_port, B2_out_7_port, 
      B2_out_6_port, B2_out_5_port, B2_out_4_port, B2_out_3_port, B2_out_2_port
      , B2_out_1_port, B2_out_0_port, ALR_in_31_port, ALR_in_30_port, 
      ALR_in_29_port, ALR_in_28_port, ALR_in_27_port, ALR_in_26_port, 
      ALR_in_25_port, ALR_in_24_port, ALR_in_23_port, ALR_in_22_port, 
      ALR_in_21_port, ALR_in_20_port, ALR_in_19_port, ALR_in_18_port, 
      ALR_in_17_port, ALR_in_16_port, ALR_in_15_port, ALR_in_14_port, 
      ALR_in_13_port, ALR_in_12_port, ALR_in_11_port, ALR_in_10_port, 
      ALR_in_9_port, ALR_in_8_port, ALR_in_7_port, ALR_in_6_port, ALR_in_5_port
      , ALR_in_4_port, ALR_in_3_port, ALR_in_2_port, ALR_in_1_port, 
      ALR_in_0_port, NPC3_out_31_port, NPC3_out_30_port, NPC3_out_29_port, 
      NPC3_out_28_port, NPC3_out_27_port, NPC3_out_26_port, NPC3_out_25_port, 
      NPC3_out_24_port, NPC3_out_23_port, NPC3_out_22_port, NPC3_out_21_port, 
      NPC3_out_20_port, NPC3_out_19_port, NPC3_out_18_port, NPC3_out_17_port, 
      NPC3_out_16_port, NPC3_out_15_port, NPC3_out_14_port, NPC3_out_13_port, 
      NPC3_out_12_port, NPC3_out_11_port, NPC3_out_10_port, NPC3_out_9_port, 
      NPC3_out_8_port, NPC3_out_7_port, NPC3_out_6_port, NPC3_out_5_port, 
      NPC3_out_4_port, NPC3_out_3_port, NPC3_out_2_port, NPC3_out_1_port, 
      NPC3_out_0_port, PSW_in_6_port, PSW_in_5_port, PSW_in_4_port, 
      PSW_in_3_port, PSW_in_2_port, PSW_in_1_port, PSW_in_0_port, 
      PSW_out_6_port, PSW_out_5_port, PSW_out_4_port, PSW_out_3_port, 
      PSW_out_2_port, PSW_out_1_port, PSW_out_0_port, MEM_ENABLE, 
      ALR2_in_31_port, ALR2_in_30_port, ALR2_in_29_port, ALR2_in_28_port, 
      ALR2_in_27_port, ALR2_in_26_port, ALR2_in_25_port, ALR2_in_24_port, 
      ALR2_in_23_port, ALR2_in_22_port, ALR2_in_21_port, ALR2_in_20_port, 
      ALR2_in_19_port, ALR2_in_18_port, ALR2_in_17_port, ALR2_in_16_port, 
      ALR2_in_15_port, ALR2_in_14_port, ALR2_in_13_port, ALR2_in_12_port, 
      ALR2_in_11_port, ALR2_in_10_port, ALR2_in_9_port, ALR2_in_8_port, 
      ALR2_in_7_port, ALR2_in_6_port, ALR2_in_5_port, ALR2_in_4_port, 
      ALR2_in_3_port, ALR2_in_2_port, ALR2_in_1_port, ALR2_in_0_port, 
      ALR2_out_31_port, ALR2_out_30_port, ALR2_out_29_port, ALR2_out_28_port, 
      ALR2_out_27_port, ALR2_out_26_port, ALR2_out_25_port, ALR2_out_24_port, 
      ALR2_out_23_port, ALR2_out_22_port, ALR2_out_21_port, ALR2_out_20_port, 
      ALR2_out_19_port, ALR2_out_18_port, ALR2_out_17_port, ALR2_out_16_port, 
      ALR2_out_15_port, ALR2_out_14_port, ALR2_out_13_port, ALR2_out_12_port, 
      ALR2_out_11_port, ALR2_out_10_port, ALR2_out_9_port, ALR2_out_8_port, 
      ALR2_out_7_port, ALR2_out_6_port, ALR2_out_5_port, ALR2_out_4_port, 
      ALR2_out_3_port, ALR2_out_2_port, ALR2_out_1_port, ALR2_out_0_port, 
      RWB3_out_20_port, RWB3_out_19_port, RWB3_out_18_port, RWB3_out_17_port, 
      RWB3_out_16_port, RWB3_out_15_port, RWB3_out_14_port, RWB3_out_13_port, 
      RWB3_out_12_port, RWB3_out_11_port, IMM_out_31_port, IMM_out_30_port, 
      IMM_out_29_port, IMM_out_28_port, IMM_out_27_port, IMM_out_26_port, 
      IMM_out_25_port, IMM_out_24_port, IMM_out_23_port, IMM_out_22_port, 
      IMM_out_21_port, IMM_out_20_port, IMM_out_19_port, IMM_out_18_port, 
      IMM_out_17_port, IMM_out_16_port, IMM_out_15_port, IMM_out_14_port, 
      IMM_out_13_port, IMM_out_12_port, IMM_out_11_port, IMM_out_10_port, 
      IMM_out_9_port, IMM_out_8_port, IMM_out_7_port, IMM_out_6_port, 
      IMM_out_5_port, IMM_out_4_port, IMM_out_3_port, IMM_out_2_port, 
      IMM_out_1_port, IMM_out_0_port, PC_SEL_1_port, PC_MUX_out_31_port, 
      PC_MUX_out_30_port, PC_MUX_out_29_port, PC_MUX_out_28_port, 
      PC_MUX_out_27_port, PC_MUX_out_26_port, PC_MUX_out_25_port, 
      PC_MUX_out_24_port, PC_MUX_out_23_port, PC_MUX_out_22_port, 
      PC_MUX_out_21_port, PC_MUX_out_20_port, PC_MUX_out_19_port, 
      PC_MUX_out_18_port, PC_MUX_out_17_port, PC_MUX_out_16_port, 
      PC_MUX_out_15_port, PC_MUX_out_14_port, PC_MUX_out_13_port, 
      PC_MUX_out_12_port, PC_MUX_out_11_port, PC_MUX_out_10_port, 
      PC_MUX_out_9_port, PC_MUX_out_8_port, PC_MUX_out_7_port, 
      PC_MUX_out_6_port, PC_MUX_out_5_port, PC_MUX_out_4_port, 
      PC_MUX_out_3_port, PC_MUX_out_2_port, PC_MUX_out_1_port, 
      PC_MUX_out_0_port, IRAMMUX_SEL, BHT_in_31_port, BHT_in_30_port, 
      BHT_in_29_port, BHT_in_28_port, BHT_in_27_port, BHT_in_26_port, 
      BHT_in_25_port, BHT_in_24_port, BHT_in_23_port, BHT_in_22_port, 
      BHT_in_21_port, BHT_in_20_port, BHT_in_19_port, BHT_in_18_port, 
      BHT_in_17_port, BHT_in_16_port, BHT_in_15_port, BHT_in_14_port, 
      BHT_in_13_port, BHT_in_12_port, BHT_in_11_port, BHT_in_10_port, 
      BHT_in_9_port, BHT_in_8_port, BHT_in_7_port, BHT_in_6_port, BHT_in_5_port
      , BHT_in_4_port, BHT_in_3_port, BHT_in_2_port, BHT_in_1_port, 
      BHT_in_0_port, FWDA_OUT_31_port, FWDA_OUT_30_port, FWDA_OUT_29_port, 
      FWDA_OUT_28_port, FWDA_OUT_27_port, FWDA_OUT_26_port, FWDA_OUT_25_port, 
      FWDA_OUT_24_port, FWDA_OUT_23_port, FWDA_OUT_22_port, FWDA_OUT_21_port, 
      FWDA_OUT_20_port, FWDA_OUT_19_port, FWDA_OUT_18_port, FWDA_OUT_17_port, 
      FWDA_OUT_16_port, FWDA_OUT_15_port, FWDA_OUT_14_port, FWDA_OUT_13_port, 
      FWDA_OUT_12_port, FWDA_OUT_11_port, FWDA_OUT_10_port, FWDA_OUT_9_port, 
      FWDA_OUT_8_port, FWDA_OUT_7_port, FWDA_OUT_6_port, FWDA_OUT_5_port, 
      FWDA_OUT_4_port, FWDA_OUT_3_port, FWDA_OUT_2_port, FWDA_OUT_1_port, 
      FWDA_OUT_0_port, A_in_31_port, A_in_30_port, A_in_29_port, A_in_28_port, 
      A_in_27_port, A_in_26_port, A_in_25_port, A_in_24_port, A_in_23_port, 
      A_in_22_port, A_in_21_port, A_in_20_port, A_in_19_port, A_in_18_port, 
      A_in_17_port, A_in_16_port, A_in_15_port, A_in_14_port, A_in_13_port, 
      A_in_12_port, A_in_11_port, A_in_10_port, A_in_9_port, A_in_8_port, 
      A_in_7_port, A_in_6_port, A_in_5_port, A_in_4_port, A_in_3_port, 
      A_in_2_port, A_in_1_port, A_in_0_port, FWDB_OUT_31_port, FWDB_OUT_30_port
      , FWDB_OUT_29_port, FWDB_OUT_28_port, FWDB_OUT_27_port, FWDB_OUT_26_port,
      FWDB_OUT_25_port, FWDB_OUT_24_port, FWDB_OUT_23_port, FWDB_OUT_22_port, 
      FWDB_OUT_21_port, FWDB_OUT_20_port, FWDB_OUT_19_port, FWDB_OUT_18_port, 
      FWDB_OUT_17_port, FWDB_OUT_16_port, FWDB_OUT_15_port, FWDB_OUT_14_port, 
      FWDB_OUT_13_port, FWDB_OUT_12_port, FWDB_OUT_11_port, FWDB_OUT_10_port, 
      FWDB_OUT_9_port, FWDB_OUT_8_port, FWDB_OUT_7_port, FWDB_OUT_6_port, 
      FWDB_OUT_5_port, FWDB_OUT_4_port, FWDB_OUT_3_port, FWDB_OUT_2_port, 
      FWDB_OUT_1_port, FWDB_OUT_0_port, B_in_31_port, B_in_30_port, 
      B_in_29_port, B_in_28_port, B_in_27_port, B_in_26_port, B_in_25_port, 
      B_in_24_port, B_in_23_port, B_in_22_port, B_in_21_port, B_in_20_port, 
      B_in_19_port, B_in_18_port, B_in_17_port, B_in_16_port, B_in_15_port, 
      B_in_14_port, B_in_13_port, B_in_12_port, B_in_11_port, B_in_10_port, 
      B_in_9_port, B_in_8_port, B_in_7_port, B_in_6_port, B_in_5_port, 
      B_in_4_port, B_in_3_port, B_in_2_port, B_in_1_port, B_in_0_port, 
      RA_out_31_port, RA_out_30_port, RA_out_29_port, RA_out_28_port, 
      RA_out_27_port, RA_out_26_port, RA_out_25_port, RA_out_24_port, 
      RA_out_23_port, RA_out_22_port, RA_out_21_port, RA_out_20_port, 
      RA_out_19_port, RA_out_18_port, RA_out_17_port, RA_out_16_port, 
      RA_out_15_port, RA_out_14_port, RA_out_13_port, RA_out_12_port, 
      RA_out_11_port, RA_out_10_port, RA_out_9_port, RA_out_8_port, 
      RA_out_7_port, RA_out_6_port, RA_out_5_port, RA_out_4_port, RA_out_3_port
      , RA_out_2_port, RA_out_1_port, RA_out_0_port, WB_in_31_port, 
      WB_in_30_port, WB_in_29_port, WB_in_28_port, WB_in_27_port, WB_in_26_port
      , WB_in_25_port, WB_in_24_port, WB_in_23_port, WB_in_22_port, 
      WB_in_21_port, WB_in_20_port, WB_in_19_port, WB_in_18_port, WB_in_17_port
      , WB_in_16_port, WB_in_15_port, WB_in_14_port, WB_in_13_port, 
      WB_in_12_port, WB_in_11_port, WB_in_10_port, WB_in_9_port, WB_in_8_port, 
      WB_in_7_port, WB_in_6_port, WB_in_5_port, WB_in_4_port, WB_in_3_port, 
      WB_in_2_port, WB_in_1_port, WB_in_0_port, FWDA_SEL_1_port, 
      FWDA_SEL_0_port, FWDB_SEL_1_port, FWDB_SEL_0_port, CWB_MUX2_out_31_port, 
      CWB_MUX2_out_30_port, CWB_MUX2_out_29_port, CWB_MUX2_out_28_port, 
      CWB_MUX2_out_27_port, CWB_MUX2_out_26_port, CWB_MUX2_out_25_port, 
      CWB_MUX2_out_24_port, CWB_MUX2_out_23_port, CWB_MUX2_out_22_port, 
      CWB_MUX2_out_21_port, CWB_MUX2_out_20_port, CWB_MUX2_out_19_port, 
      CWB_MUX2_out_18_port, CWB_MUX2_out_17_port, CWB_MUX2_out_16_port, 
      CWB_MUX2_out_15_port, CWB_MUX2_out_14_port, CWB_MUX2_out_13_port, 
      CWB_MUX2_out_12_port, CWB_MUX2_out_11_port, CWB_MUX2_out_10_port, 
      CWB_MUX2_out_9_port, CWB_MUX2_out_8_port, CWB_MUX2_out_7_port, 
      CWB_MUX2_out_6_port, CWB_MUX2_out_5_port, CWB_MUX2_out_4_port, 
      CWB_MUX2_out_3_port, CWB_MUX2_out_2_port, CWB_MUX2_out_1_port, 
      CWB_MUX2_out_0_port, ZDU_SEL_1_port, ZDU_SEL_0_port, ZDU_MUX_out_30_port,
      ZDU_MUX_out_29_port, ZDU_MUX_out_28_port, ZDU_MUX_out_27_port, 
      ZDU_MUX_out_26_port, ZDU_MUX_out_25_port, ZDU_MUX_out_24_port, 
      ZDU_MUX_out_23_port, ZDU_MUX_out_22_port, ZDU_MUX_out_21_port, 
      ZDU_MUX_out_20_port, ZDU_MUX_out_19_port, ZDU_MUX_out_18_port, 
      ZDU_MUX_out_17_port, ZDU_MUX_out_16_port, ZDU_MUX_out_15_port, 
      ZDU_MUX_out_14_port, ZDU_MUX_out_13_port, ZDU_MUX_out_12_port, 
      ZDU_MUX_out_11_port, ZDU_MUX_out_10_port, ZDU_MUX_out_9_port, 
      ZDU_MUX_out_8_port, ZDU_MUX_out_7_port, ZDU_MUX_out_6_port, 
      ZDU_MUX_out_5_port, ZDU_MUX_out_4_port, ZDU_MUX_out_3_port, 
      ZDU_MUX_out_2_port, ZDU_MUX_out_1_port, ZDU_MUX_out_0_port, 
      B2_MUX_out_31_port, B2_MUX_out_30_port, B2_MUX_out_29_port, 
      B2_MUX_out_28_port, B2_MUX_out_27_port, B2_MUX_out_26_port, 
      B2_MUX_out_25_port, B2_MUX_out_24_port, B2_MUX_out_23_port, 
      B2_MUX_out_22_port, B2_MUX_out_21_port, B2_MUX_out_20_port, 
      B2_MUX_out_19_port, B2_MUX_out_18_port, B2_MUX_out_17_port, 
      B2_MUX_out_16_port, B2_MUX_out_15_port, B2_MUX_out_14_port, 
      B2_MUX_out_13_port, B2_MUX_out_12_port, B2_MUX_out_11_port, 
      B2_MUX_out_10_port, B2_MUX_out_9_port, B2_MUX_out_8_port, 
      B2_MUX_out_7_port, B2_MUX_out_6_port, B2_MUX_out_5_port, 
      B2_MUX_out_4_port, B2_MUX_out_3_port, B2_MUX_out_2_port, 
      B2_MUX_out_1_port, B2_MUX_out_0_port, LMD_out_31_port, LMD_out_30_port, 
      LMD_out_29_port, LMD_out_28_port, LMD_out_27_port, LMD_out_26_port, 
      LMD_out_25_port, LMD_out_24_port, LMD_out_23_port, LMD_out_22_port, 
      LMD_out_21_port, LMD_out_20_port, LMD_out_19_port, LMD_out_18_port, 
      LMD_out_17_port, LMD_out_16_port, LMD_out_15_port, LMD_out_14_port, 
      LMD_out_13_port, LMD_out_12_port, LMD_out_11_port, LMD_out_10_port, 
      LMD_out_9_port, LMD_out_8_port, LMD_out_7_port, LMD_out_6_port, 
      LMD_out_5_port, LMD_out_4_port, LMD_out_3_port, LMD_out_2_port, 
      LMD_out_1_port, LMD_out_0_port, CWB_out_1_port, CWB_out_0_port, 
      CWB_MUX_SEL_1_port, CWB_MUX_SEL_0_port, CWB2_SEL_1_port, CWB2_SEL_0_port,
      FWDB2_SEL, RF_MUX_out_4_port, RF_MUX_out_3_port, RF_MUX_out_2_port, 
      RF_MUX_out_1_port, RF_MUX_out_0_port, IF_STALL, EX_STALL, MEM_STALL, 
      ZDU_out, RF_RD_en, N14, n13, n14_port, n15, n16, n17, n18, n1, n2, n3, n4
      , n5, n6, n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664 : 
      std_logic;

begin
   IRAM_ADDR <= ( IRAM_ADDR_31_port, IRAM_ADDR_30_port, IRAM_ADDR_29_port, 
      IRAM_ADDR_28_port, IRAM_ADDR_27_port, IRAM_ADDR_26_port, 
      IRAM_ADDR_25_port, IRAM_ADDR_24_port, IRAM_ADDR_23_port, 
      IRAM_ADDR_22_port, IRAM_ADDR_21_port, IRAM_ADDR_20_port, 
      IRAM_ADDR_19_port, IRAM_ADDR_18_port, IRAM_ADDR_17_port, 
      IRAM_ADDR_16_port, IRAM_ADDR_15_port, IRAM_ADDR_14_port, 
      IRAM_ADDR_13_port, IRAM_ADDR_12_port, IRAM_ADDR_11_port, 
      IRAM_ADDR_10_port, IRAM_ADDR_9_port, IRAM_ADDR_8_port, IRAM_ADDR_7_port, 
      IRAM_ADDR_6_port, IRAM_ADDR_5_port, IRAM_ADDR_4_port, IRAM_ADDR_3_port, 
      IRAM_ADDR_2_port, IRAM_ADDR_1_port, IRAM_ADDR_0_port );
   DATA_ADDR <= ( DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RegPC : REG_NBIT32_0 port map( clk => CLK, reset => n7, enable => n11, 
                           data_in(31) => NPC_in_31_port, data_in(30) => 
                           NPC_in_30_port, data_in(29) => NPC_in_29_port, 
                           data_in(28) => NPC_in_28_port, data_in(27) => 
                           NPC_in_27_port, data_in(26) => NPC_in_26_port, 
                           data_in(25) => NPC_in_25_port, data_in(24) => 
                           NPC_in_24_port, data_in(23) => NPC_in_23_port, 
                           data_in(22) => NPC_in_22_port, data_in(21) => 
                           NPC_in_21_port, data_in(20) => NPC_in_20_port, 
                           data_in(19) => NPC_in_19_port, data_in(18) => 
                           NPC_in_18_port, data_in(17) => NPC_in_17_port, 
                           data_in(16) => NPC_in_16_port, data_in(15) => 
                           NPC_in_15_port, data_in(14) => NPC_in_14_port, 
                           data_in(13) => NPC_in_13_port, data_in(12) => 
                           NPC_in_12_port, data_in(11) => NPC_in_11_port, 
                           data_in(10) => NPC_in_10_port, data_in(9) => 
                           NPC_in_9_port, data_in(8) => NPC_in_8_port, 
                           data_in(7) => NPC_in_7_port, data_in(6) => 
                           NPC_in_6_port, data_in(5) => NPC_in_5_port, 
                           data_in(4) => NPC_in_4_port, data_in(3) => 
                           NPC_in_3_port, data_in(2) => NPC_in_2_port, 
                           data_in(1) => NPC_in_1_port, data_in(0) => 
                           NPC_in_0_port, data_out(31) => PC_out_31_port, 
                           data_out(30) => PC_out_30_port, data_out(29) => 
                           PC_out_29_port, data_out(28) => PC_out_28_port, 
                           data_out(27) => PC_out_27_port, data_out(26) => 
                           PC_out_26_port, data_out(25) => PC_out_25_port, 
                           data_out(24) => PC_out_24_port, data_out(23) => 
                           PC_out_23_port, data_out(22) => PC_out_22_port, 
                           data_out(21) => PC_out_21_port, data_out(20) => 
                           PC_out_20_port, data_out(19) => PC_out_19_port, 
                           data_out(18) => PC_out_18_port, data_out(17) => 
                           PC_out_17_port, data_out(16) => PC_out_16_port, 
                           data_out(15) => PC_out_15_port, data_out(14) => 
                           PC_out_14_port, data_out(13) => PC_out_13_port, 
                           data_out(12) => PC_out_12_port, data_out(11) => 
                           PC_out_11_port, data_out(10) => PC_out_10_port, 
                           data_out(9) => PC_out_9_port, data_out(8) => 
                           PC_out_8_port, data_out(7) => PC_out_7_port, 
                           data_out(6) => PC_out_6_port, data_out(5) => 
                           PC_out_5_port, data_out(4) => PC_out_4_port, 
                           data_out(3) => PC_out_3_port, data_out(2) => 
                           PC_out_2_port, data_out(1) => PC_out_1_port, 
                           data_out(0) => PC_out_0_port);
   RegIR : REG_NBIT32_17 port map( clk => CLK, reset => n9, enable => n11, 
                           data_in(31) => IRAM_OUT(31), data_in(30) => 
                           IRAM_OUT(30), data_in(29) => IRAM_OUT(29), 
                           data_in(28) => IRAM_OUT(28), data_in(27) => 
                           IRAM_OUT(27), data_in(26) => IRAM_OUT(26), 
                           data_in(25) => IRAM_OUT(25), data_in(24) => 
                           IRAM_OUT(24), data_in(23) => IRAM_OUT(23), 
                           data_in(22) => IRAM_OUT(22), data_in(21) => 
                           IRAM_OUT(21), data_in(20) => IRAM_OUT(20), 
                           data_in(19) => IRAM_OUT(19), data_in(18) => 
                           IRAM_OUT(18), data_in(17) => IRAM_OUT(17), 
                           data_in(16) => IRAM_OUT(16), data_in(15) => 
                           IRAM_OUT(15), data_in(14) => IRAM_OUT(14), 
                           data_in(13) => IRAM_OUT(13), data_in(12) => 
                           IRAM_OUT(12), data_in(11) => IRAM_OUT(11), 
                           data_in(10) => IRAM_OUT(10), data_in(9) => 
                           IRAM_OUT(9), data_in(8) => IRAM_OUT(8), data_in(7) 
                           => IRAM_OUT(7), data_in(6) => IRAM_OUT(6), 
                           data_in(5) => IRAM_OUT(5), data_in(4) => IRAM_OUT(4)
                           , data_in(3) => IRAM_OUT(3), data_in(2) => 
                           IRAM_OUT(2), data_in(1) => IRAM_OUT(1), data_in(0) 
                           => IRAM_OUT(0), data_out(31) => IR_out_31_port, 
                           data_out(30) => IR_out_30_port, data_out(29) => 
                           IR_out_29_port, data_out(28) => IR_out_28_port, 
                           data_out(27) => IR_out_27_port, data_out(26) => 
                           IR_out_26_port, data_out(25) => IR_out_25_port, 
                           data_out(24) => IR_out_24_port, data_out(23) => 
                           IR_out_23_port, data_out(22) => IR_out_22_port, 
                           data_out(21) => IR_out_21_port, data_out(20) => 
                           IR_out_20_port, data_out(19) => IR_out_19_port, 
                           data_out(18) => IR_out_18_port, data_out(17) => 
                           IR_out_17_port, data_out(16) => IR_out_16_port, 
                           data_out(15) => IR_out_15_port, data_out(14) => 
                           IR_out_14_port, data_out(13) => IR_out_13_port, 
                           data_out(12) => IR_out_12_port, data_out(11) => 
                           IR_out_11_port, data_out(10) => IR_out_10_port, 
                           data_out(9) => IR_out_9_port, data_out(8) => 
                           IR_out_8_port, data_out(7) => IR_out_7_port, 
                           data_out(6) => IR_out_6_port, data_out(5) => 
                           IR_out_5_port, data_out(4) => IR_out_4_port, 
                           data_out(3) => IR_out_3_port, data_out(2) => 
                           IR_out_2_port, data_out(1) => IR_out_1_port, 
                           data_out(0) => IR_out_0_port);
   RegNPC : REG_NBIT32_16 port map( clk => CLK, reset => n8, enable => n11, 
                           data_in(31) => NPC_in_31_port, data_in(30) => 
                           NPC_in_30_port, data_in(29) => NPC_in_29_port, 
                           data_in(28) => NPC_in_28_port, data_in(27) => 
                           NPC_in_27_port, data_in(26) => NPC_in_26_port, 
                           data_in(25) => NPC_in_25_port, data_in(24) => 
                           NPC_in_24_port, data_in(23) => NPC_in_23_port, 
                           data_in(22) => NPC_in_22_port, data_in(21) => 
                           NPC_in_21_port, data_in(20) => NPC_in_20_port, 
                           data_in(19) => NPC_in_19_port, data_in(18) => 
                           NPC_in_18_port, data_in(17) => NPC_in_17_port, 
                           data_in(16) => NPC_in_16_port, data_in(15) => 
                           NPC_in_15_port, data_in(14) => NPC_in_14_port, 
                           data_in(13) => NPC_in_13_port, data_in(12) => 
                           NPC_in_12_port, data_in(11) => NPC_in_11_port, 
                           data_in(10) => NPC_in_10_port, data_in(9) => 
                           NPC_in_9_port, data_in(8) => NPC_in_8_port, 
                           data_in(7) => NPC_in_7_port, data_in(6) => 
                           NPC_in_6_port, data_in(5) => NPC_in_5_port, 
                           data_in(4) => NPC_in_4_port, data_in(3) => 
                           NPC_in_3_port, data_in(2) => NPC_in_2_port, 
                           data_in(1) => NPC_in_1_port, data_in(0) => 
                           NPC_in_0_port, data_out(31) => NPC_out_31_port, 
                           data_out(30) => NPC_out_30_port, data_out(29) => 
                           NPC_out_29_port, data_out(28) => NPC_out_28_port, 
                           data_out(27) => NPC_out_27_port, data_out(26) => 
                           NPC_out_26_port, data_out(25) => NPC_out_25_port, 
                           data_out(24) => NPC_out_24_port, data_out(23) => 
                           NPC_out_23_port, data_out(22) => NPC_out_22_port, 
                           data_out(21) => NPC_out_21_port, data_out(20) => 
                           NPC_out_20_port, data_out(19) => NPC_out_19_port, 
                           data_out(18) => NPC_out_18_port, data_out(17) => 
                           NPC_out_17_port, data_out(16) => NPC_out_16_port, 
                           data_out(15) => NPC_out_15_port, data_out(14) => 
                           NPC_out_14_port, data_out(13) => NPC_out_13_port, 
                           data_out(12) => NPC_out_12_port, data_out(11) => 
                           NPC_out_11_port, data_out(10) => NPC_out_10_port, 
                           data_out(9) => NPC_out_9_port, data_out(8) => 
                           NPC_out_8_port, data_out(7) => NPC_out_7_port, 
                           data_out(6) => NPC_out_6_port, data_out(5) => 
                           NPC_out_5_port, data_out(4) => NPC_out_4_port, 
                           data_out(3) => NPC_out_3_port, data_out(2) => 
                           NPC_out_2_port, data_out(1) => NPC_out_1_port, 
                           data_out(0) => NPC_out_0_port);
   RegPC2 : REG_NBIT32_15 port map( clk => CLK, reset => n9, enable => n21, 
                           data_in(31) => PC_out_31_port, data_in(30) => 
                           PC_out_30_port, data_in(29) => PC_out_29_port, 
                           data_in(28) => PC_out_28_port, data_in(27) => 
                           PC_out_27_port, data_in(26) => PC_out_26_port, 
                           data_in(25) => PC_out_25_port, data_in(24) => 
                           PC_out_24_port, data_in(23) => PC_out_23_port, 
                           data_in(22) => PC_out_22_port, data_in(21) => 
                           PC_out_21_port, data_in(20) => PC_out_20_port, 
                           data_in(19) => PC_out_19_port, data_in(18) => 
                           PC_out_18_port, data_in(17) => PC_out_17_port, 
                           data_in(16) => PC_out_16_port, data_in(15) => 
                           PC_out_15_port, data_in(14) => PC_out_14_port, 
                           data_in(13) => PC_out_13_port, data_in(12) => 
                           PC_out_12_port, data_in(11) => PC_out_11_port, 
                           data_in(10) => PC_out_10_port, data_in(9) => 
                           PC_out_9_port, data_in(8) => PC_out_8_port, 
                           data_in(7) => PC_out_7_port, data_in(6) => 
                           PC_out_6_port, data_in(5) => PC_out_5_port, 
                           data_in(4) => PC_out_4_port, data_in(3) => 
                           PC_out_3_port, data_in(2) => PC_out_2_port, 
                           data_in(1) => PC_out_1_port, data_in(0) => 
                           PC_out_0_port, data_out(31) => PC2_out_31_port, 
                           data_out(30) => PC2_out_30_port, data_out(29) => 
                           PC2_out_29_port, data_out(28) => PC2_out_28_port, 
                           data_out(27) => PC2_out_27_port, data_out(26) => 
                           PC2_out_26_port, data_out(25) => PC2_out_25_port, 
                           data_out(24) => PC2_out_24_port, data_out(23) => 
                           PC2_out_23_port, data_out(22) => PC2_out_22_port, 
                           data_out(21) => PC2_out_21_port, data_out(20) => 
                           PC2_out_20_port, data_out(19) => PC2_out_19_port, 
                           data_out(18) => PC2_out_18_port, data_out(17) => 
                           PC2_out_17_port, data_out(16) => PC2_out_16_port, 
                           data_out(15) => PC2_out_15_port, data_out(14) => 
                           PC2_out_14_port, data_out(13) => PC2_out_13_port, 
                           data_out(12) => PC2_out_12_port, data_out(11) => 
                           PC2_out_11_port, data_out(10) => PC2_out_10_port, 
                           data_out(9) => PC2_out_9_port, data_out(8) => 
                           PC2_out_8_port, data_out(7) => PC2_out_7_port, 
                           data_out(6) => PC2_out_6_port, data_out(5) => 
                           PC2_out_5_port, data_out(4) => PC2_out_4_port, 
                           data_out(3) => PC2_out_3_port, data_out(2) => 
                           PC2_out_2_port, data_out(1) => PC2_out_1_port, 
                           data_out(0) => PC2_out_0_port);
   RegIMM : REG_NBIT32_14 port map( clk => CLK, reset => n10, enable => n21, 
                           data_in(31) => N14, data_in(30) => N14, data_in(29) 
                           => N14, data_in(28) => N14, data_in(27) => N14, 
                           data_in(26) => N14, data_in(25) => N14, data_in(24) 
                           => N14, data_in(23) => N14, data_in(22) => N14, 
                           data_in(21) => N14, data_in(20) => N14, data_in(19) 
                           => N14, data_in(18) => N14, data_in(17) => N14, 
                           data_in(16) => N14, data_in(15) => IR_out_15_port, 
                           data_in(14) => IR_out_14_port, data_in(13) => 
                           IR_out_13_port, data_in(12) => IR_out_12_port, 
                           data_in(11) => IR_out_11_port, data_in(10) => 
                           IR_out_10_port, data_in(9) => IR_out_9_port, 
                           data_in(8) => IR_out_8_port, data_in(7) => 
                           IR_out_7_port, data_in(6) => IR_out_6_port, 
                           data_in(5) => IR_out_5_port, data_in(4) => 
                           IR_out_4_port, data_in(3) => IR_out_3_port, 
                           data_in(2) => IR_out_2_port, data_in(1) => 
                           IR_out_1_port, data_in(0) => IR_out_0_port, 
                           data_out(31) => RIMM_out_31_port, data_out(30) => 
                           RIMM_out_30_port, data_out(29) => RIMM_out_29_port, 
                           data_out(28) => RIMM_out_28_port, data_out(27) => 
                           RIMM_out_27_port, data_out(26) => RIMM_out_26_port, 
                           data_out(25) => RIMM_out_25_port, data_out(24) => 
                           RIMM_out_24_port, data_out(23) => RIMM_out_23_port, 
                           data_out(22) => RIMM_out_22_port, data_out(21) => 
                           RIMM_out_21_port, data_out(20) => RIMM_out_20_port, 
                           data_out(19) => RIMM_out_19_port, data_out(18) => 
                           RIMM_out_18_port, data_out(17) => RIMM_out_17_port, 
                           data_out(16) => RIMM_out_16_port, data_out(15) => 
                           RIMM_out_15_port, data_out(14) => RIMM_out_14_port, 
                           data_out(13) => RIMM_out_13_port, data_out(12) => 
                           RIMM_out_12_port, data_out(11) => RIMM_out_11_port, 
                           data_out(10) => RIMM_out_10_port, data_out(9) => 
                           RIMM_out_9_port, data_out(8) => RIMM_out_8_port, 
                           data_out(7) => RIMM_out_7_port, data_out(6) => 
                           RIMM_out_6_port, data_out(5) => RIMM_out_5_port, 
                           data_out(4) => RIMM_out_4_port, data_out(3) => 
                           RIMM_out_3_port, data_out(2) => RIMM_out_2_port, 
                           data_out(1) => RIMM_out_1_port, data_out(0) => 
                           RIMM_out_0_port);
   RegWB1 : REG_NBIT32_13 port map( clk => CLK, reset => n8, enable => n21, 
                           data_in(31) => IR_out_31_port, data_in(30) => 
                           IR_out_30_port, data_in(29) => IR_out_29_port, 
                           data_in(28) => IR_out_28_port, data_in(27) => 
                           IR_out_27_port, data_in(26) => IR_out_26_port, 
                           data_in(25) => IR_out_25_port, data_in(24) => 
                           IR_out_24_port, data_in(23) => IR_out_23_port, 
                           data_in(22) => IR_out_22_port, data_in(21) => 
                           IR_out_21_port, data_in(20) => IR_out_20_port, 
                           data_in(19) => IR_out_19_port, data_in(18) => 
                           IR_out_18_port, data_in(17) => IR_out_17_port, 
                           data_in(16) => IR_out_16_port, data_in(15) => 
                           IR_out_15_port, data_in(14) => IR_out_14_port, 
                           data_in(13) => IR_out_13_port, data_in(12) => 
                           IR_out_12_port, data_in(11) => IR_out_11_port, 
                           data_in(10) => IR_out_10_port, data_in(9) => 
                           IR_out_9_port, data_in(8) => IR_out_8_port, 
                           data_in(7) => IR_out_7_port, data_in(6) => 
                           IR_out_6_port, data_in(5) => IR_out_5_port, 
                           data_in(4) => IR_out_4_port, data_in(3) => 
                           IR_out_3_port, data_in(2) => IR_out_2_port, 
                           data_in(1) => IR_out_1_port, data_in(0) => 
                           IR_out_0_port, data_out(31) => RWB1_out_31_port, 
                           data_out(30) => RWB1_out_30_port, data_out(29) => 
                           RWB1_out_29_port, data_out(28) => RWB1_out_28_port, 
                           data_out(27) => RWB1_out_27_port, data_out(26) => 
                           RWB1_out_26_port, data_out(25) => RWB1_out_25_port, 
                           data_out(24) => RWB1_out_24_port, data_out(23) => 
                           RWB1_out_23_port, data_out(22) => RWB1_out_22_port, 
                           data_out(21) => RWB1_out_21_port, data_out(20) => 
                           RWB1_out_20_port, data_out(19) => RWB1_out_19_port, 
                           data_out(18) => RWB1_out_18_port, data_out(17) => 
                           RWB1_out_17_port, data_out(16) => RWB1_out_16_port, 
                           data_out(15) => RWB1_out_15_port, data_out(14) => 
                           RWB1_out_14_port, data_out(13) => RWB1_out_13_port, 
                           data_out(12) => RWB1_out_12_port, data_out(11) => 
                           RWB1_out_11_port, data_out(10) => RWB1_out_10_port, 
                           data_out(9) => RWB1_out_9_port, data_out(8) => 
                           RWB1_out_8_port, data_out(7) => RWB1_out_7_port, 
                           data_out(6) => RWB1_out_6_port, data_out(5) => 
                           RWB1_out_5_port, data_out(4) => RWB1_out_4_port, 
                           data_out(3) => RWB1_out_3_port, data_out(2) => 
                           RWB1_out_2_port, data_out(1) => RWB1_out_1_port, 
                           data_out(0) => RWB1_out_0_port);
   F_PRD : FFD_0 port map( D => BHT_out, CK => CLK, RESET => n6, ENABLE => n21,
                           Q => PRD_OUT);
   RegNPC2 : REG_NBIT32_12 port map( clk => CLK, reset => n10, enable => n21, 
                           data_in(31) => NPC_out_31_port, data_in(30) => 
                           NPC_out_30_port, data_in(29) => NPC_out_29_port, 
                           data_in(28) => NPC_out_28_port, data_in(27) => 
                           NPC_out_27_port, data_in(26) => NPC_out_26_port, 
                           data_in(25) => NPC_out_25_port, data_in(24) => 
                           NPC_out_24_port, data_in(23) => NPC_out_23_port, 
                           data_in(22) => NPC_out_22_port, data_in(21) => 
                           NPC_out_21_port, data_in(20) => NPC_out_20_port, 
                           data_in(19) => NPC_out_19_port, data_in(18) => 
                           NPC_out_18_port, data_in(17) => NPC_out_17_port, 
                           data_in(16) => NPC_out_16_port, data_in(15) => 
                           NPC_out_15_port, data_in(14) => NPC_out_14_port, 
                           data_in(13) => NPC_out_13_port, data_in(12) => 
                           NPC_out_12_port, data_in(11) => NPC_out_11_port, 
                           data_in(10) => NPC_out_10_port, data_in(9) => 
                           NPC_out_9_port, data_in(8) => NPC_out_8_port, 
                           data_in(7) => NPC_out_7_port, data_in(6) => 
                           NPC_out_6_port, data_in(5) => NPC_out_5_port, 
                           data_in(4) => NPC_out_4_port, data_in(3) => 
                           NPC_out_3_port, data_in(2) => NPC_out_2_port, 
                           data_in(1) => NPC_out_1_port, data_in(0) => 
                           NPC_out_0_port, data_out(31) => NPC2_out_31_port, 
                           data_out(30) => NPC2_out_30_port, data_out(29) => 
                           NPC2_out_29_port, data_out(28) => NPC2_out_28_port, 
                           data_out(27) => NPC2_out_27_port, data_out(26) => 
                           NPC2_out_26_port, data_out(25) => NPC2_out_25_port, 
                           data_out(24) => NPC2_out_24_port, data_out(23) => 
                           NPC2_out_23_port, data_out(22) => NPC2_out_22_port, 
                           data_out(21) => NPC2_out_21_port, data_out(20) => 
                           NPC2_out_20_port, data_out(19) => NPC2_out_19_port, 
                           data_out(18) => NPC2_out_18_port, data_out(17) => 
                           NPC2_out_17_port, data_out(16) => NPC2_out_16_port, 
                           data_out(15) => NPC2_out_15_port, data_out(14) => 
                           NPC2_out_14_port, data_out(13) => NPC2_out_13_port, 
                           data_out(12) => NPC2_out_12_port, data_out(11) => 
                           NPC2_out_11_port, data_out(10) => NPC2_out_10_port, 
                           data_out(9) => NPC2_out_9_port, data_out(8) => 
                           NPC2_out_8_port, data_out(7) => NPC2_out_7_port, 
                           data_out(6) => NPC2_out_6_port, data_out(5) => 
                           NPC2_out_5_port, data_out(4) => NPC2_out_4_port, 
                           data_out(3) => NPC2_out_3_port, data_out(2) => 
                           NPC2_out_2_port, data_out(1) => NPC2_out_1_port, 
                           data_out(0) => NPC2_out_0_port);
   RegJADD2 : REG_NBIT32_11 port map( clk => CLK, reset => n8, enable => n21, 
                           data_in(31) => JADDER_out_31_port, data_in(30) => 
                           JADDER_out_30_port, data_in(29) => 
                           JADDER_out_29_port, data_in(28) => 
                           JADDER_out_28_port, data_in(27) => 
                           JADDER_out_27_port, data_in(26) => 
                           JADDER_out_26_port, data_in(25) => 
                           JADDER_out_25_port, data_in(24) => 
                           JADDER_out_24_port, data_in(23) => 
                           JADDER_out_23_port, data_in(22) => 
                           JADDER_out_22_port, data_in(21) => 
                           JADDER_out_21_port, data_in(20) => 
                           JADDER_out_20_port, data_in(19) => 
                           JADDER_out_19_port, data_in(18) => 
                           JADDER_out_18_port, data_in(17) => 
                           JADDER_out_17_port, data_in(16) => 
                           JADDER_out_16_port, data_in(15) => 
                           JADDER_out_15_port, data_in(14) => 
                           JADDER_out_14_port, data_in(13) => 
                           JADDER_out_13_port, data_in(12) => 
                           JADDER_out_12_port, data_in(11) => 
                           JADDER_out_11_port, data_in(10) => 
                           JADDER_out_10_port, data_in(9) => JADDER_out_9_port,
                           data_in(8) => JADDER_out_8_port, data_in(7) => 
                           JADDER_out_7_port, data_in(6) => JADDER_out_6_port, 
                           data_in(5) => JADDER_out_5_port, data_in(4) => 
                           JADDER_out_4_port, data_in(3) => JADDER_out_3_port, 
                           data_in(2) => JADDER_out_2_port, data_in(1) => 
                           JADDER_out_1_port, data_in(0) => JADDER_out_0_port, 
                           data_out(31) => JADDER2_out_31_port, data_out(30) =>
                           JADDER2_out_30_port, data_out(29) => 
                           JADDER2_out_29_port, data_out(28) => 
                           JADDER2_out_28_port, data_out(27) => 
                           JADDER2_out_27_port, data_out(26) => 
                           JADDER2_out_26_port, data_out(25) => 
                           JADDER2_out_25_port, data_out(24) => 
                           JADDER2_out_24_port, data_out(23) => 
                           JADDER2_out_23_port, data_out(22) => 
                           JADDER2_out_22_port, data_out(21) => 
                           JADDER2_out_21_port, data_out(20) => 
                           JADDER2_out_20_port, data_out(19) => 
                           JADDER2_out_19_port, data_out(18) => 
                           JADDER2_out_18_port, data_out(17) => 
                           JADDER2_out_17_port, data_out(16) => 
                           JADDER2_out_16_port, data_out(15) => 
                           JADDER2_out_15_port, data_out(14) => 
                           JADDER2_out_14_port, data_out(13) => 
                           JADDER2_out_13_port, data_out(12) => 
                           JADDER2_out_12_port, data_out(11) => 
                           JADDER2_out_11_port, data_out(10) => 
                           JADDER2_out_10_port, data_out(9) => 
                           JADDER2_out_9_port, data_out(8) => 
                           JADDER2_out_8_port, data_out(7) => 
                           JADDER2_out_7_port, data_out(6) => 
                           JADDER2_out_6_port, data_out(5) => 
                           JADDER2_out_5_port, data_out(4) => 
                           JADDER2_out_4_port, data_out(3) => 
                           JADDER2_out_3_port, data_out(2) => 
                           JADDER2_out_2_port, data_out(1) => 
                           JADDER2_out_1_port, data_out(0) => 
                           JADDER2_out_0_port);
   F_JR : FFD_1 port map( D => BPR_EN, CK => CLK, RESET => n7, ENABLE => n21, Q
                           => BPR_EN2);
   RegPC3 : REG_NBIT32_10 port map( clk => CLK, reset => n9, enable => n19, 
                           data_in(31) => PC2_out_31_port, data_in(30) => 
                           PC2_out_30_port, data_in(29) => PC2_out_29_port, 
                           data_in(28) => PC2_out_28_port, data_in(27) => 
                           PC2_out_27_port, data_in(26) => PC2_out_26_port, 
                           data_in(25) => PC2_out_25_port, data_in(24) => 
                           PC2_out_24_port, data_in(23) => PC2_out_23_port, 
                           data_in(22) => PC2_out_22_port, data_in(21) => 
                           PC2_out_21_port, data_in(20) => PC2_out_20_port, 
                           data_in(19) => PC2_out_19_port, data_in(18) => 
                           PC2_out_18_port, data_in(17) => PC2_out_17_port, 
                           data_in(16) => PC2_out_16_port, data_in(15) => 
                           PC2_out_15_port, data_in(14) => PC2_out_14_port, 
                           data_in(13) => PC2_out_13_port, data_in(12) => 
                           PC2_out_12_port, data_in(11) => PC2_out_11_port, 
                           data_in(10) => PC2_out_10_port, data_in(9) => 
                           PC2_out_9_port, data_in(8) => PC2_out_8_port, 
                           data_in(7) => PC2_out_7_port, data_in(6) => 
                           PC2_out_6_port, data_in(5) => PC2_out_5_port, 
                           data_in(4) => PC2_out_4_port, data_in(3) => 
                           PC2_out_3_port, data_in(2) => PC2_out_2_port, 
                           data_in(1) => n2, data_in(0) => n1, data_out(31) => 
                           PC3_out_31_port, data_out(30) => PC3_out_30_port, 
                           data_out(29) => PC3_out_29_port, data_out(28) => 
                           PC3_out_28_port, data_out(27) => PC3_out_27_port, 
                           data_out(26) => PC3_out_26_port, data_out(25) => 
                           PC3_out_25_port, data_out(24) => PC3_out_24_port, 
                           data_out(23) => PC3_out_23_port, data_out(22) => 
                           PC3_out_22_port, data_out(21) => PC3_out_21_port, 
                           data_out(20) => PC3_out_20_port, data_out(19) => 
                           PC3_out_19_port, data_out(18) => PC3_out_18_port, 
                           data_out(17) => PC3_out_17_port, data_out(16) => 
                           PC3_out_16_port, data_out(15) => PC3_out_15_port, 
                           data_out(14) => PC3_out_14_port, data_out(13) => 
                           PC3_out_13_port, data_out(12) => PC3_out_12_port, 
                           data_out(11) => PC3_out_11_port, data_out(10) => 
                           PC3_out_10_port, data_out(9) => PC3_out_9_port, 
                           data_out(8) => PC3_out_8_port, data_out(7) => 
                           PC3_out_7_port, data_out(6) => PC3_out_6_port, 
                           data_out(5) => PC3_out_5_port, data_out(4) => 
                           PC3_out_4_port, data_out(3) => PC3_out_3_port, 
                           data_out(2) => PC3_out_2_port, data_out(1) => 
                           PC3_out_1_port, data_out(0) => PC3_out_0_port);
   RegWB2 : REG_NBIT32_9 port map( clk => CLK, reset => n5, enable => n19, 
                           data_in(31) => RWB1_out_31_port, data_in(30) => 
                           RWB1_out_30_port, data_in(29) => RWB1_out_29_port, 
                           data_in(28) => RWB1_out_28_port, data_in(27) => 
                           RWB1_out_27_port, data_in(26) => RWB1_out_26_port, 
                           data_in(25) => RWB1_out_25_port, data_in(24) => 
                           RWB1_out_24_port, data_in(23) => RWB1_out_23_port, 
                           data_in(22) => RWB1_out_22_port, data_in(21) => 
                           RWB1_out_21_port, data_in(20) => RWB1_out_20_port, 
                           data_in(19) => RWB1_out_19_port, data_in(18) => 
                           RWB1_out_18_port, data_in(17) => RWB1_out_17_port, 
                           data_in(16) => RWB1_out_16_port, data_in(15) => 
                           RWB1_out_15_port, data_in(14) => RWB1_out_14_port, 
                           data_in(13) => RWB1_out_13_port, data_in(12) => 
                           RWB1_out_12_port, data_in(11) => RWB1_out_11_port, 
                           data_in(10) => RWB1_out_10_port, data_in(9) => 
                           RWB1_out_9_port, data_in(8) => RWB1_out_8_port, 
                           data_in(7) => RWB1_out_7_port, data_in(6) => 
                           RWB1_out_6_port, data_in(5) => RWB1_out_5_port, 
                           data_in(4) => RWB1_out_4_port, data_in(3) => 
                           RWB1_out_3_port, data_in(2) => RWB1_out_2_port, 
                           data_in(1) => RWB1_out_1_port, data_in(0) => 
                           RWB1_out_0_port, data_out(31) => RWB2_out_31_port, 
                           data_out(30) => RWB2_out_30_port, data_out(29) => 
                           RWB2_out_29_port, data_out(28) => RWB2_out_28_port, 
                           data_out(27) => RWB2_out_27_port, data_out(26) => 
                           RWB2_out_26_port, data_out(25) => RWB2_out_25_port, 
                           data_out(24) => RWB2_out_24_port, data_out(23) => 
                           RWB2_out_23_port, data_out(22) => RWB2_out_22_port, 
                           data_out(21) => RWB2_out_21_port, data_out(20) => 
                           RWB2_out_20_port, data_out(19) => RWB2_out_19_port, 
                           data_out(18) => RWB2_out_18_port, data_out(17) => 
                           RWB2_out_17_port, data_out(16) => RWB2_out_16_port, 
                           data_out(15) => RWB2_out_15_port, data_out(14) => 
                           RWB2_out_14_port, data_out(13) => RWB2_out_13_port, 
                           data_out(12) => RWB2_out_12_port, data_out(11) => 
                           RWB2_out_11_port, data_out(10) => RWB2_out_10_port, 
                           data_out(9) => RWB2_out_9_port, data_out(8) => 
                           RWB2_out_8_port, data_out(7) => RWB2_out_7_port, 
                           data_out(6) => RWB2_out_6_port, data_out(5) => 
                           RWB2_out_5_port, data_out(4) => RWB2_out_4_port, 
                           data_out(3) => RWB2_out_3_port, data_out(2) => 
                           RWB2_out_2_port, data_out(1) => RWB2_out_1_port, 
                           data_out(0) => RWB2_out_0_port);
   RegB2 : REG_NBIT32_8 port map( clk => CLK, reset => n6, enable => n19, 
                           data_in(31) => RB_out_31_port, data_in(30) => 
                           RB_out_30_port, data_in(29) => RB_out_29_port, 
                           data_in(28) => RB_out_28_port, data_in(27) => 
                           RB_out_27_port, data_in(26) => RB_out_26_port, 
                           data_in(25) => RB_out_25_port, data_in(24) => 
                           RB_out_24_port, data_in(23) => RB_out_23_port, 
                           data_in(22) => RB_out_22_port, data_in(21) => 
                           RB_out_21_port, data_in(20) => RB_out_20_port, 
                           data_in(19) => RB_out_19_port, data_in(18) => 
                           RB_out_18_port, data_in(17) => RB_out_17_port, 
                           data_in(16) => RB_out_16_port, data_in(15) => 
                           RB_out_15_port, data_in(14) => RB_out_14_port, 
                           data_in(13) => RB_out_13_port, data_in(12) => 
                           RB_out_12_port, data_in(11) => RB_out_11_port, 
                           data_in(10) => RB_out_10_port, data_in(9) => 
                           RB_out_9_port, data_in(8) => RB_out_8_port, 
                           data_in(7) => RB_out_7_port, data_in(6) => 
                           RB_out_6_port, data_in(5) => RB_out_5_port, 
                           data_in(4) => RB_out_4_port, data_in(3) => 
                           RB_out_3_port, data_in(2) => RB_out_2_port, 
                           data_in(1) => RB_out_1_port, data_in(0) => 
                           RB_out_0_port, data_out(31) => B2_out_31_port, 
                           data_out(30) => B2_out_30_port, data_out(29) => 
                           B2_out_29_port, data_out(28) => B2_out_28_port, 
                           data_out(27) => B2_out_27_port, data_out(26) => 
                           B2_out_26_port, data_out(25) => B2_out_25_port, 
                           data_out(24) => B2_out_24_port, data_out(23) => 
                           B2_out_23_port, data_out(22) => B2_out_22_port, 
                           data_out(21) => B2_out_21_port, data_out(20) => 
                           B2_out_20_port, data_out(19) => B2_out_19_port, 
                           data_out(18) => B2_out_18_port, data_out(17) => 
                           B2_out_17_port, data_out(16) => B2_out_16_port, 
                           data_out(15) => B2_out_15_port, data_out(14) => 
                           B2_out_14_port, data_out(13) => B2_out_13_port, 
                           data_out(12) => B2_out_12_port, data_out(11) => 
                           B2_out_11_port, data_out(10) => B2_out_10_port, 
                           data_out(9) => B2_out_9_port, data_out(8) => 
                           B2_out_8_port, data_out(7) => B2_out_7_port, 
                           data_out(6) => B2_out_6_port, data_out(5) => 
                           B2_out_5_port, data_out(4) => B2_out_4_port, 
                           data_out(3) => B2_out_3_port, data_out(2) => 
                           B2_out_2_port, data_out(1) => B2_out_1_port, 
                           data_out(0) => B2_out_0_port);
   RegALR : REG_NBIT32_7 port map( clk => CLK, reset => n5, enable => n19, 
                           data_in(31) => ALR_in_31_port, data_in(30) => 
                           ALR_in_30_port, data_in(29) => ALR_in_29_port, 
                           data_in(28) => ALR_in_28_port, data_in(27) => 
                           ALR_in_27_port, data_in(26) => ALR_in_26_port, 
                           data_in(25) => ALR_in_25_port, data_in(24) => 
                           ALR_in_24_port, data_in(23) => ALR_in_23_port, 
                           data_in(22) => ALR_in_22_port, data_in(21) => 
                           ALR_in_21_port, data_in(20) => ALR_in_20_port, 
                           data_in(19) => ALR_in_19_port, data_in(18) => 
                           ALR_in_18_port, data_in(17) => ALR_in_17_port, 
                           data_in(16) => ALR_in_16_port, data_in(15) => 
                           ALR_in_15_port, data_in(14) => ALR_in_14_port, 
                           data_in(13) => ALR_in_13_port, data_in(12) => 
                           ALR_in_12_port, data_in(11) => ALR_in_11_port, 
                           data_in(10) => ALR_in_10_port, data_in(9) => 
                           ALR_in_9_port, data_in(8) => ALR_in_8_port, 
                           data_in(7) => ALR_in_7_port, data_in(6) => 
                           ALR_in_6_port, data_in(5) => ALR_in_5_port, 
                           data_in(4) => ALR_in_4_port, data_in(3) => 
                           ALR_in_3_port, data_in(2) => ALR_in_2_port, 
                           data_in(1) => ALR_in_1_port, data_in(0) => 
                           ALR_in_0_port, data_out(31) => DATA_ADDR_31_port, 
                           data_out(30) => DATA_ADDR_30_port, data_out(29) => 
                           DATA_ADDR_29_port, data_out(28) => DATA_ADDR_28_port
                           , data_out(27) => DATA_ADDR_27_port, data_out(26) =>
                           DATA_ADDR_26_port, data_out(25) => DATA_ADDR_25_port
                           , data_out(24) => DATA_ADDR_24_port, data_out(23) =>
                           DATA_ADDR_23_port, data_out(22) => DATA_ADDR_22_port
                           , data_out(21) => DATA_ADDR_21_port, data_out(20) =>
                           DATA_ADDR_20_port, data_out(19) => DATA_ADDR_19_port
                           , data_out(18) => DATA_ADDR_18_port, data_out(17) =>
                           DATA_ADDR_17_port, data_out(16) => DATA_ADDR_16_port
                           , data_out(15) => DATA_ADDR_15_port, data_out(14) =>
                           DATA_ADDR_14_port, data_out(13) => DATA_ADDR_13_port
                           , data_out(12) => DATA_ADDR_12_port, data_out(11) =>
                           DATA_ADDR_11_port, data_out(10) => DATA_ADDR_10_port
                           , data_out(9) => DATA_ADDR_9_port, data_out(8) => 
                           DATA_ADDR_8_port, data_out(7) => DATA_ADDR_7_port, 
                           data_out(6) => DATA_ADDR_6_port, data_out(5) => 
                           DATA_ADDR_5_port, data_out(4) => DATA_ADDR_4_port, 
                           data_out(3) => DATA_ADDR_3_port, data_out(2) => 
                           DATA_ADDR_2_port, data_out(1) => DATA_ADDR_1_port, 
                           data_out(0) => DATA_ADDR_0_port);
   RegNPC3 : REG_NBIT32_6 port map( clk => CLK, reset => n6, enable => n19, 
                           data_in(31) => NPC2_out_31_port, data_in(30) => 
                           NPC2_out_30_port, data_in(29) => NPC2_out_29_port, 
                           data_in(28) => NPC2_out_28_port, data_in(27) => 
                           NPC2_out_27_port, data_in(26) => NPC2_out_26_port, 
                           data_in(25) => NPC2_out_25_port, data_in(24) => 
                           NPC2_out_24_port, data_in(23) => NPC2_out_23_port, 
                           data_in(22) => NPC2_out_22_port, data_in(21) => 
                           NPC2_out_21_port, data_in(20) => NPC2_out_20_port, 
                           data_in(19) => NPC2_out_19_port, data_in(18) => 
                           NPC2_out_18_port, data_in(17) => NPC2_out_17_port, 
                           data_in(16) => NPC2_out_16_port, data_in(15) => 
                           NPC2_out_15_port, data_in(14) => NPC2_out_14_port, 
                           data_in(13) => NPC2_out_13_port, data_in(12) => 
                           NPC2_out_12_port, data_in(11) => NPC2_out_11_port, 
                           data_in(10) => NPC2_out_10_port, data_in(9) => 
                           NPC2_out_9_port, data_in(8) => NPC2_out_8_port, 
                           data_in(7) => NPC2_out_7_port, data_in(6) => 
                           NPC2_out_6_port, data_in(5) => NPC2_out_5_port, 
                           data_in(4) => NPC2_out_4_port, data_in(3) => 
                           NPC2_out_3_port, data_in(2) => NPC2_out_2_port, 
                           data_in(1) => NPC2_out_1_port, data_in(0) => 
                           NPC2_out_0_port, data_out(31) => NPC3_out_31_port, 
                           data_out(30) => NPC3_out_30_port, data_out(29) => 
                           NPC3_out_29_port, data_out(28) => NPC3_out_28_port, 
                           data_out(27) => NPC3_out_27_port, data_out(26) => 
                           NPC3_out_26_port, data_out(25) => NPC3_out_25_port, 
                           data_out(24) => NPC3_out_24_port, data_out(23) => 
                           NPC3_out_23_port, data_out(22) => NPC3_out_22_port, 
                           data_out(21) => NPC3_out_21_port, data_out(20) => 
                           NPC3_out_20_port, data_out(19) => NPC3_out_19_port, 
                           data_out(18) => NPC3_out_18_port, data_out(17) => 
                           NPC3_out_17_port, data_out(16) => NPC3_out_16_port, 
                           data_out(15) => NPC3_out_15_port, data_out(14) => 
                           NPC3_out_14_port, data_out(13) => NPC3_out_13_port, 
                           data_out(12) => NPC3_out_12_port, data_out(11) => 
                           NPC3_out_11_port, data_out(10) => NPC3_out_10_port, 
                           data_out(9) => NPC3_out_9_port, data_out(8) => 
                           NPC3_out_8_port, data_out(7) => NPC3_out_7_port, 
                           data_out(6) => NPC3_out_6_port, data_out(5) => 
                           NPC3_out_5_port, data_out(4) => NPC3_out_4_port, 
                           data_out(3) => NPC3_out_3_port, data_out(2) => 
                           NPC3_out_2_port, data_out(1) => NPC3_out_1_port, 
                           data_out(0) => NPC3_out_0_port);
   RegPSW : REG_NBIT7 port map( clk => CLK, reset => n6, enable => n19, 
                           data_in(6) => PSW_in_6_port, data_in(5) => 
                           PSW_in_5_port, data_in(4) => PSW_in_4_port, 
                           data_in(3) => PSW_in_3_port, data_in(2) => 
                           PSW_in_2_port, data_in(1) => PSW_in_1_port, 
                           data_in(0) => PSW_in_0_port, data_out(6) => 
                           PSW_out_6_port, data_out(5) => PSW_out_5_port, 
                           data_out(4) => PSW_out_4_port, data_out(3) => 
                           PSW_out_3_port, data_out(2) => PSW_out_2_port, 
                           data_out(1) => PSW_out_1_port, data_out(0) => 
                           PSW_out_0_port);
   RegALR2 : REG_NBIT32_5 port map( clk => CLK, reset => n7, enable => n12, 
                           data_in(31) => ALR2_in_31_port, data_in(30) => 
                           ALR2_in_30_port, data_in(29) => ALR2_in_29_port, 
                           data_in(28) => ALR2_in_28_port, data_in(27) => 
                           ALR2_in_27_port, data_in(26) => ALR2_in_26_port, 
                           data_in(25) => ALR2_in_25_port, data_in(24) => 
                           ALR2_in_24_port, data_in(23) => ALR2_in_23_port, 
                           data_in(22) => ALR2_in_22_port, data_in(21) => 
                           ALR2_in_21_port, data_in(20) => ALR2_in_20_port, 
                           data_in(19) => ALR2_in_19_port, data_in(18) => 
                           ALR2_in_18_port, data_in(17) => ALR2_in_17_port, 
                           data_in(16) => ALR2_in_16_port, data_in(15) => 
                           ALR2_in_15_port, data_in(14) => ALR2_in_14_port, 
                           data_in(13) => ALR2_in_13_port, data_in(12) => 
                           ALR2_in_12_port, data_in(11) => ALR2_in_11_port, 
                           data_in(10) => ALR2_in_10_port, data_in(9) => 
                           ALR2_in_9_port, data_in(8) => ALR2_in_8_port, 
                           data_in(7) => ALR2_in_7_port, data_in(6) => 
                           ALR2_in_6_port, data_in(5) => ALR2_in_5_port, 
                           data_in(4) => ALR2_in_4_port, data_in(3) => 
                           ALR2_in_3_port, data_in(2) => ALR2_in_2_port, 
                           data_in(1) => ALR2_in_1_port, data_in(0) => 
                           ALR2_in_0_port, data_out(31) => ALR2_out_31_port, 
                           data_out(30) => ALR2_out_30_port, data_out(29) => 
                           ALR2_out_29_port, data_out(28) => ALR2_out_28_port, 
                           data_out(27) => ALR2_out_27_port, data_out(26) => 
                           ALR2_out_26_port, data_out(25) => ALR2_out_25_port, 
                           data_out(24) => ALR2_out_24_port, data_out(23) => 
                           ALR2_out_23_port, data_out(22) => ALR2_out_22_port, 
                           data_out(21) => ALR2_out_21_port, data_out(20) => 
                           ALR2_out_20_port, data_out(19) => ALR2_out_19_port, 
                           data_out(18) => ALR2_out_18_port, data_out(17) => 
                           ALR2_out_17_port, data_out(16) => ALR2_out_16_port, 
                           data_out(15) => ALR2_out_15_port, data_out(14) => 
                           ALR2_out_14_port, data_out(13) => ALR2_out_13_port, 
                           data_out(12) => ALR2_out_12_port, data_out(11) => 
                           ALR2_out_11_port, data_out(10) => ALR2_out_10_port, 
                           data_out(9) => ALR2_out_9_port, data_out(8) => 
                           ALR2_out_8_port, data_out(7) => ALR2_out_7_port, 
                           data_out(6) => ALR2_out_6_port, data_out(5) => 
                           ALR2_out_5_port, data_out(4) => ALR2_out_4_port, 
                           data_out(3) => ALR2_out_3_port, data_out(2) => 
                           ALR2_out_2_port, data_out(1) => ALR2_out_1_port, 
                           data_out(0) => ALR2_out_0_port);
   RegWB3 : REG_NBIT32_4 port map( clk => CLK, reset => n5, enable => n12, 
                           data_in(31) => RWB2_out_31_port, data_in(30) => 
                           RWB2_out_30_port, data_in(29) => RWB2_out_29_port, 
                           data_in(28) => RWB2_out_28_port, data_in(27) => 
                           RWB2_out_27_port, data_in(26) => RWB2_out_26_port, 
                           data_in(25) => RWB2_out_25_port, data_in(24) => 
                           RWB2_out_24_port, data_in(23) => RWB2_out_23_port, 
                           data_in(22) => RWB2_out_22_port, data_in(21) => 
                           RWB2_out_21_port, data_in(20) => RWB2_out_20_port, 
                           data_in(19) => RWB2_out_19_port, data_in(18) => 
                           RWB2_out_18_port, data_in(17) => RWB2_out_17_port, 
                           data_in(16) => RWB2_out_16_port, data_in(15) => 
                           RWB2_out_15_port, data_in(14) => RWB2_out_14_port, 
                           data_in(13) => RWB2_out_13_port, data_in(12) => 
                           RWB2_out_12_port, data_in(11) => RWB2_out_11_port, 
                           data_in(10) => RWB2_out_10_port, data_in(9) => 
                           RWB2_out_9_port, data_in(8) => RWB2_out_8_port, 
                           data_in(7) => RWB2_out_7_port, data_in(6) => 
                           RWB2_out_6_port, data_in(5) => RWB2_out_5_port, 
                           data_in(4) => RWB2_out_4_port, data_in(3) => 
                           RWB2_out_3_port, data_in(2) => RWB2_out_2_port, 
                           data_in(1) => RWB2_out_1_port, data_in(0) => 
                           RWB2_out_0_port, data_out(31) => n_1640, 
                           data_out(30) => n_1641, data_out(29) => n_1642, 
                           data_out(28) => n_1643, data_out(27) => n_1644, 
                           data_out(26) => n_1645, data_out(25) => n_1646, 
                           data_out(24) => n_1647, data_out(23) => n_1648, 
                           data_out(22) => n_1649, data_out(21) => n_1650, 
                           data_out(20) => RWB3_out_20_port, data_out(19) => 
                           RWB3_out_19_port, data_out(18) => RWB3_out_18_port, 
                           data_out(17) => RWB3_out_17_port, data_out(16) => 
                           RWB3_out_16_port, data_out(15) => RWB3_out_15_port, 
                           data_out(14) => RWB3_out_14_port, data_out(13) => 
                           RWB3_out_13_port, data_out(12) => RWB3_out_12_port, 
                           data_out(11) => RWB3_out_11_port, data_out(10) => 
                           n_1651, data_out(9) => n_1652, data_out(8) => n_1653
                           , data_out(7) => n_1654, data_out(6) => n_1655, 
                           data_out(5) => n_1656, data_out(4) => n_1657, 
                           data_out(3) => n_1658, data_out(2) => n_1659, 
                           data_out(1) => n_1660, data_out(0) => n_1661);
   AdderPC : PC_adder_0 port map( A(31) => IRAM_ADDR_31_port, A(30) => 
                           IRAM_ADDR_30_port, A(29) => IRAM_ADDR_29_port, A(28)
                           => IRAM_ADDR_28_port, A(27) => IRAM_ADDR_27_port, 
                           A(26) => IRAM_ADDR_26_port, A(25) => 
                           IRAM_ADDR_25_port, A(24) => IRAM_ADDR_24_port, A(23)
                           => IRAM_ADDR_23_port, A(22) => IRAM_ADDR_22_port, 
                           A(21) => IRAM_ADDR_21_port, A(20) => 
                           IRAM_ADDR_20_port, A(19) => IRAM_ADDR_19_port, A(18)
                           => IRAM_ADDR_18_port, A(17) => IRAM_ADDR_17_port, 
                           A(16) => IRAM_ADDR_16_port, A(15) => 
                           IRAM_ADDR_15_port, A(14) => IRAM_ADDR_14_port, A(13)
                           => IRAM_ADDR_13_port, A(12) => IRAM_ADDR_12_port, 
                           A(11) => IRAM_ADDR_11_port, A(10) => 
                           IRAM_ADDR_10_port, A(9) => IRAM_ADDR_9_port, A(8) =>
                           IRAM_ADDR_8_port, A(7) => IRAM_ADDR_7_port, A(6) => 
                           IRAM_ADDR_6_port, A(5) => IRAM_ADDR_5_port, A(4) => 
                           IRAM_ADDR_4_port, A(3) => IRAM_ADDR_3_port, A(2) => 
                           IRAM_ADDR_2_port, A(1) => IRAM_ADDR_1_port, A(0) => 
                           IRAM_ADDR_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, Sum(31) => NPC_in_31_port, Sum(30) =>
                           NPC_in_30_port, Sum(29) => NPC_in_29_port, Sum(28) 
                           => NPC_in_28_port, Sum(27) => NPC_in_27_port, 
                           Sum(26) => NPC_in_26_port, Sum(25) => NPC_in_25_port
                           , Sum(24) => NPC_in_24_port, Sum(23) => 
                           NPC_in_23_port, Sum(22) => NPC_in_22_port, Sum(21) 
                           => NPC_in_21_port, Sum(20) => NPC_in_20_port, 
                           Sum(19) => NPC_in_19_port, Sum(18) => NPC_in_18_port
                           , Sum(17) => NPC_in_17_port, Sum(16) => 
                           NPC_in_16_port, Sum(15) => NPC_in_15_port, Sum(14) 
                           => NPC_in_14_port, Sum(13) => NPC_in_13_port, 
                           Sum(12) => NPC_in_12_port, Sum(11) => NPC_in_11_port
                           , Sum(10) => NPC_in_10_port, Sum(9) => NPC_in_9_port
                           , Sum(8) => NPC_in_8_port, Sum(7) => NPC_in_7_port, 
                           Sum(6) => NPC_in_6_port, Sum(5) => NPC_in_5_port, 
                           Sum(4) => NPC_in_4_port, Sum(3) => NPC_in_3_port, 
                           Sum(2) => NPC_in_2_port, Sum(1) => NPC_in_1_port, 
                           Sum(0) => NPC_in_0_port);
   J_Adder : PC_adder_1 port map( A(31) => PC2_out_31_port, A(30) => 
                           PC2_out_30_port, A(29) => PC2_out_29_port, A(28) => 
                           PC2_out_28_port, A(27) => PC2_out_27_port, A(26) => 
                           PC2_out_26_port, A(25) => PC2_out_25_port, A(24) => 
                           PC2_out_24_port, A(23) => PC2_out_23_port, A(22) => 
                           PC2_out_22_port, A(21) => PC2_out_21_port, A(20) => 
                           PC2_out_20_port, A(19) => PC2_out_19_port, A(18) => 
                           PC2_out_18_port, A(17) => PC2_out_17_port, A(16) => 
                           PC2_out_16_port, A(15) => PC2_out_15_port, A(14) => 
                           PC2_out_14_port, A(13) => PC2_out_13_port, A(12) => 
                           PC2_out_12_port, A(11) => PC2_out_11_port, A(10) => 
                           PC2_out_10_port, A(9) => PC2_out_9_port, A(8) => 
                           PC2_out_8_port, A(7) => PC2_out_7_port, A(6) => 
                           PC2_out_6_port, A(5) => PC2_out_5_port, A(4) => 
                           PC2_out_4_port, A(3) => PC2_out_3_port, A(2) => 
                           PC2_out_2_port, A(1) => n2, A(0) => n1, B(31) => 
                           IMM_out_31_port, B(30) => IMM_out_30_port, B(29) => 
                           IMM_out_29_port, B(28) => IMM_out_28_port, B(27) => 
                           IMM_out_27_port, B(26) => IMM_out_26_port, B(25) => 
                           IMM_out_25_port, B(24) => IMM_out_24_port, B(23) => 
                           IMM_out_23_port, B(22) => IMM_out_22_port, B(21) => 
                           IMM_out_21_port, B(20) => IMM_out_20_port, B(19) => 
                           IMM_out_19_port, B(18) => IMM_out_18_port, B(17) => 
                           IMM_out_17_port, B(16) => IMM_out_16_port, B(15) => 
                           IMM_out_15_port, B(14) => IMM_out_14_port, B(13) => 
                           IMM_out_13_port, B(12) => IMM_out_12_port, B(11) => 
                           IMM_out_11_port, B(10) => IMM_out_10_port, B(9) => 
                           IMM_out_9_port, B(8) => IMM_out_8_port, B(7) => 
                           IMM_out_7_port, B(6) => IMM_out_6_port, B(5) => 
                           IMM_out_5_port, B(4) => IMM_out_4_port, B(3) => 
                           IMM_out_3_port, B(2) => IMM_out_2_port, B(1) => 
                           IMM_out_1_port, B(0) => IMM_out_0_port, Sum(31) => 
                           JADDER_out_31_port, Sum(30) => JADDER_out_30_port, 
                           Sum(29) => JADDER_out_29_port, Sum(28) => 
                           JADDER_out_28_port, Sum(27) => JADDER_out_27_port, 
                           Sum(26) => JADDER_out_26_port, Sum(25) => 
                           JADDER_out_25_port, Sum(24) => JADDER_out_24_port, 
                           Sum(23) => JADDER_out_23_port, Sum(22) => 
                           JADDER_out_22_port, Sum(21) => JADDER_out_21_port, 
                           Sum(20) => JADDER_out_20_port, Sum(19) => 
                           JADDER_out_19_port, Sum(18) => JADDER_out_18_port, 
                           Sum(17) => JADDER_out_17_port, Sum(16) => 
                           JADDER_out_16_port, Sum(15) => JADDER_out_15_port, 
                           Sum(14) => JADDER_out_14_port, Sum(13) => 
                           JADDER_out_13_port, Sum(12) => JADDER_out_12_port, 
                           Sum(11) => JADDER_out_11_port, Sum(10) => 
                           JADDER_out_10_port, Sum(9) => JADDER_out_9_port, 
                           Sum(8) => JADDER_out_8_port, Sum(7) => 
                           JADDER_out_7_port, Sum(6) => JADDER_out_6_port, 
                           Sum(5) => JADDER_out_5_port, Sum(4) => 
                           JADDER_out_4_port, Sum(3) => JADDER_out_3_port, 
                           Sum(2) => JADDER_out_2_port, Sum(1) => 
                           JADDER_out_1_port, Sum(0) => JADDER_out_0_port);
   PCMUX : MUX3to1_NBIT32_0 port map( A(31) => PC_out_31_port, A(30) => 
                           PC_out_30_port, A(29) => PC_out_29_port, A(28) => 
                           PC_out_28_port, A(27) => PC_out_27_port, A(26) => 
                           PC_out_26_port, A(25) => PC_out_25_port, A(24) => 
                           PC_out_24_port, A(23) => PC_out_23_port, A(22) => 
                           PC_out_22_port, A(21) => PC_out_21_port, A(20) => 
                           PC_out_20_port, A(19) => PC_out_19_port, A(18) => 
                           PC_out_18_port, A(17) => PC_out_17_port, A(16) => 
                           PC_out_16_port, A(15) => PC_out_15_port, A(14) => 
                           PC_out_14_port, A(13) => PC_out_13_port, A(12) => 
                           PC_out_12_port, A(11) => PC_out_11_port, A(10) => 
                           PC_out_10_port, A(9) => PC_out_9_port, A(8) => 
                           PC_out_8_port, A(7) => PC_out_7_port, A(6) => 
                           PC_out_6_port, A(5) => PC_out_5_port, A(4) => 
                           PC_out_4_port, A(3) => PC_out_3_port, A(2) => 
                           PC_out_2_port, A(1) => PC_out_1_port, A(0) => 
                           PC_out_0_port, B(31) => JADDER_out_31_port, B(30) =>
                           JADDER_out_30_port, B(29) => JADDER_out_29_port, 
                           B(28) => JADDER_out_28_port, B(27) => 
                           JADDER_out_27_port, B(26) => JADDER_out_26_port, 
                           B(25) => JADDER_out_25_port, B(24) => 
                           JADDER_out_24_port, B(23) => JADDER_out_23_port, 
                           B(22) => JADDER_out_22_port, B(21) => 
                           JADDER_out_21_port, B(20) => JADDER_out_20_port, 
                           B(19) => JADDER_out_19_port, B(18) => 
                           JADDER_out_18_port, B(17) => JADDER_out_17_port, 
                           B(16) => JADDER_out_16_port, B(15) => 
                           JADDER_out_15_port, B(14) => JADDER_out_14_port, 
                           B(13) => JADDER_out_13_port, B(12) => 
                           JADDER_out_12_port, B(11) => JADDER_out_11_port, 
                           B(10) => JADDER_out_10_port, B(9) => 
                           JADDER_out_9_port, B(8) => JADDER_out_8_port, B(7) 
                           => JADDER_out_7_port, B(6) => JADDER_out_6_port, 
                           B(5) => JADDER_out_5_port, B(4) => JADDER_out_4_port
                           , B(3) => JADDER_out_3_port, B(2) => 
                           JADDER_out_2_port, B(1) => JADDER_out_1_port, B(0) 
                           => JADDER_out_0_port, C(31) => JADDER2_out_31_port, 
                           C(30) => JADDER2_out_30_port, C(29) => 
                           JADDER2_out_29_port, C(28) => JADDER2_out_28_port, 
                           C(27) => JADDER2_out_27_port, C(26) => 
                           JADDER2_out_26_port, C(25) => JADDER2_out_25_port, 
                           C(24) => JADDER2_out_24_port, C(23) => 
                           JADDER2_out_23_port, C(22) => JADDER2_out_22_port, 
                           C(21) => JADDER2_out_21_port, C(20) => 
                           JADDER2_out_20_port, C(19) => JADDER2_out_19_port, 
                           C(18) => JADDER2_out_18_port, C(17) => 
                           JADDER2_out_17_port, C(16) => JADDER2_out_16_port, 
                           C(15) => JADDER2_out_15_port, C(14) => 
                           JADDER2_out_14_port, C(13) => JADDER2_out_13_port, 
                           C(12) => JADDER2_out_12_port, C(11) => 
                           JADDER2_out_11_port, C(10) => JADDER2_out_10_port, 
                           C(9) => JADDER2_out_9_port, C(8) => 
                           JADDER2_out_8_port, C(7) => JADDER2_out_7_port, C(6)
                           => JADDER2_out_6_port, C(5) => JADDER2_out_5_port, 
                           C(4) => JADDER2_out_4_port, C(3) => 
                           JADDER2_out_3_port, C(2) => JADDER2_out_2_port, C(1)
                           => JADDER2_out_1_port, C(0) => JADDER2_out_0_port, 
                           SEL(1) => PC_SEL_1_port, SEL(0) => n40, Y(31) => 
                           PC_MUX_out_31_port, Y(30) => PC_MUX_out_30_port, 
                           Y(29) => PC_MUX_out_29_port, Y(28) => 
                           PC_MUX_out_28_port, Y(27) => PC_MUX_out_27_port, 
                           Y(26) => PC_MUX_out_26_port, Y(25) => 
                           PC_MUX_out_25_port, Y(24) => PC_MUX_out_24_port, 
                           Y(23) => PC_MUX_out_23_port, Y(22) => 
                           PC_MUX_out_22_port, Y(21) => PC_MUX_out_21_port, 
                           Y(20) => PC_MUX_out_20_port, Y(19) => 
                           PC_MUX_out_19_port, Y(18) => PC_MUX_out_18_port, 
                           Y(17) => PC_MUX_out_17_port, Y(16) => 
                           PC_MUX_out_16_port, Y(15) => PC_MUX_out_15_port, 
                           Y(14) => PC_MUX_out_14_port, Y(13) => 
                           PC_MUX_out_13_port, Y(12) => PC_MUX_out_12_port, 
                           Y(11) => PC_MUX_out_11_port, Y(10) => 
                           PC_MUX_out_10_port, Y(9) => PC_MUX_out_9_port, Y(8) 
                           => PC_MUX_out_8_port, Y(7) => PC_MUX_out_7_port, 
                           Y(6) => PC_MUX_out_6_port, Y(5) => PC_MUX_out_5_port
                           , Y(4) => PC_MUX_out_4_port, Y(3) => 
                           PC_MUX_out_3_port, Y(2) => PC_MUX_out_2_port, Y(1) 
                           => PC_MUX_out_1_port, Y(0) => PC_MUX_out_0_port);
   IRAMMUX : MUX2to1_NBIT32_0 port map( A(31) => PC_MUX_out_31_port, A(30) => 
                           PC_MUX_out_30_port, A(29) => PC_MUX_out_29_port, 
                           A(28) => PC_MUX_out_28_port, A(27) => 
                           PC_MUX_out_27_port, A(26) => PC_MUX_out_26_port, 
                           A(25) => PC_MUX_out_25_port, A(24) => 
                           PC_MUX_out_24_port, A(23) => PC_MUX_out_23_port, 
                           A(22) => PC_MUX_out_22_port, A(21) => 
                           PC_MUX_out_21_port, A(20) => PC_MUX_out_20_port, 
                           A(19) => PC_MUX_out_19_port, A(18) => 
                           PC_MUX_out_18_port, A(17) => PC_MUX_out_17_port, 
                           A(16) => PC_MUX_out_16_port, A(15) => 
                           PC_MUX_out_15_port, A(14) => PC_MUX_out_14_port, 
                           A(13) => PC_MUX_out_13_port, A(12) => 
                           PC_MUX_out_12_port, A(11) => PC_MUX_out_11_port, 
                           A(10) => PC_MUX_out_10_port, A(9) => 
                           PC_MUX_out_9_port, A(8) => PC_MUX_out_8_port, A(7) 
                           => PC_MUX_out_7_port, A(6) => PC_MUX_out_6_port, 
                           A(5) => PC_MUX_out_5_port, A(4) => PC_MUX_out_4_port
                           , A(3) => PC_MUX_out_3_port, A(2) => 
                           PC_MUX_out_2_port, A(1) => PC_MUX_out_1_port, A(0) 
                           => PC_MUX_out_0_port, B(31) => NPC2_out_31_port, 
                           B(30) => NPC2_out_30_port, B(29) => NPC2_out_29_port
                           , B(28) => NPC2_out_28_port, B(27) => 
                           NPC2_out_27_port, B(26) => NPC2_out_26_port, B(25) 
                           => NPC2_out_25_port, B(24) => NPC2_out_24_port, 
                           B(23) => NPC2_out_23_port, B(22) => NPC2_out_22_port
                           , B(21) => NPC2_out_21_port, B(20) => 
                           NPC2_out_20_port, B(19) => NPC2_out_19_port, B(18) 
                           => NPC2_out_18_port, B(17) => NPC2_out_17_port, 
                           B(16) => NPC2_out_16_port, B(15) => NPC2_out_15_port
                           , B(14) => NPC2_out_14_port, B(13) => 
                           NPC2_out_13_port, B(12) => NPC2_out_12_port, B(11) 
                           => NPC2_out_11_port, B(10) => NPC2_out_10_port, B(9)
                           => NPC2_out_9_port, B(8) => NPC2_out_8_port, B(7) =>
                           NPC2_out_7_port, B(6) => NPC2_out_6_port, B(5) => 
                           NPC2_out_5_port, B(4) => NPC2_out_4_port, B(3) => 
                           NPC2_out_3_port, B(2) => NPC2_out_2_port, B(1) => 
                           NPC2_out_1_port, B(0) => NPC2_out_0_port, SEL => 
                           IRAMMUX_SEL, Y(31) => IRAM_ADDR_31_port, Y(30) => 
                           IRAM_ADDR_30_port, Y(29) => IRAM_ADDR_29_port, Y(28)
                           => IRAM_ADDR_28_port, Y(27) => IRAM_ADDR_27_port, 
                           Y(26) => IRAM_ADDR_26_port, Y(25) => 
                           IRAM_ADDR_25_port, Y(24) => IRAM_ADDR_24_port, Y(23)
                           => IRAM_ADDR_23_port, Y(22) => IRAM_ADDR_22_port, 
                           Y(21) => IRAM_ADDR_21_port, Y(20) => 
                           IRAM_ADDR_20_port, Y(19) => IRAM_ADDR_19_port, Y(18)
                           => IRAM_ADDR_18_port, Y(17) => IRAM_ADDR_17_port, 
                           Y(16) => IRAM_ADDR_16_port, Y(15) => 
                           IRAM_ADDR_15_port, Y(14) => IRAM_ADDR_14_port, Y(13)
                           => IRAM_ADDR_13_port, Y(12) => IRAM_ADDR_12_port, 
                           Y(11) => IRAM_ADDR_11_port, Y(10) => 
                           IRAM_ADDR_10_port, Y(9) => IRAM_ADDR_9_port, Y(8) =>
                           IRAM_ADDR_8_port, Y(7) => IRAM_ADDR_7_port, Y(6) => 
                           IRAM_ADDR_6_port, Y(5) => IRAM_ADDR_5_port, Y(4) => 
                           IRAM_ADDR_4_port, Y(3) => IRAM_ADDR_3_port, Y(2) => 
                           IRAM_ADDR_2_port, Y(1) => IRAM_ADDR_1_port, Y(0) => 
                           IRAM_ADDR_0_port);
   IMMMUX : MUX2to1_NBIT32_8 port map( A(31) => IR_out_15_port, A(30) => 
                           IR_out_15_port, A(29) => IR_out_15_port, A(28) => 
                           IR_out_15_port, A(27) => IR_out_15_port, A(26) => 
                           IR_out_15_port, A(25) => IR_out_15_port, A(24) => 
                           IR_out_15_port, A(23) => IR_out_15_port, A(22) => 
                           IR_out_15_port, A(21) => IR_out_15_port, A(20) => 
                           IR_out_15_port, A(19) => IR_out_15_port, A(18) => 
                           IR_out_15_port, A(17) => IR_out_15_port, A(16) => 
                           IR_out_15_port, A(15) => IR_out_15_port, A(14) => 
                           IR_out_14_port, A(13) => IR_out_13_port, A(12) => 
                           IR_out_12_port, A(11) => IR_out_11_port, A(10) => 
                           IR_out_10_port, A(9) => IR_out_9_port, A(8) => 
                           IR_out_8_port, A(7) => IR_out_7_port, A(6) => 
                           IR_out_6_port, A(5) => IR_out_5_port, A(4) => 
                           IR_out_4_port, A(3) => IR_out_3_port, A(2) => 
                           IR_out_2_port, A(1) => IR_out_1_port, A(0) => 
                           IR_out_0_port, B(31) => IR_out_25_port, B(30) => 
                           IR_out_25_port, B(29) => IR_out_25_port, B(28) => 
                           IR_out_25_port, B(27) => IR_out_25_port, B(26) => 
                           IR_out_25_port, B(25) => IR_out_25_port, B(24) => 
                           IR_out_24_port, B(23) => IR_out_23_port, B(22) => 
                           IR_out_22_port, B(21) => IR_out_21_port, B(20) => 
                           IR_out_20_port, B(19) => IR_out_19_port, B(18) => 
                           IR_out_18_port, B(17) => IR_out_17_port, B(16) => 
                           IR_out_16_port, B(15) => IR_out_15_port, B(14) => 
                           IR_out_14_port, B(13) => IR_out_13_port, B(12) => 
                           IR_out_12_port, B(11) => IR_out_11_port, B(10) => 
                           IR_out_10_port, B(9) => IR_out_9_port, B(8) => 
                           IR_out_8_port, B(7) => IR_out_7_port, B(6) => 
                           IR_out_6_port, B(5) => IR_out_5_port, B(4) => 
                           IR_out_4_port, B(3) => IR_out_3_port, B(2) => 
                           IR_out_2_port, B(1) => IR_out_1_port, B(0) => 
                           IR_out_0_port, SEL => IMM_SEL, Y(31) => 
                           IMM_out_31_port, Y(30) => IMM_out_30_port, Y(29) => 
                           IMM_out_29_port, Y(28) => IMM_out_28_port, Y(27) => 
                           IMM_out_27_port, Y(26) => IMM_out_26_port, Y(25) => 
                           IMM_out_25_port, Y(24) => IMM_out_24_port, Y(23) => 
                           IMM_out_23_port, Y(22) => IMM_out_22_port, Y(21) => 
                           IMM_out_21_port, Y(20) => IMM_out_20_port, Y(19) => 
                           IMM_out_19_port, Y(18) => IMM_out_18_port, Y(17) => 
                           IMM_out_17_port, Y(16) => IMM_out_16_port, Y(15) => 
                           IMM_out_15_port, Y(14) => IMM_out_14_port, Y(13) => 
                           IMM_out_13_port, Y(12) => IMM_out_12_port, Y(11) => 
                           IMM_out_11_port, Y(10) => IMM_out_10_port, Y(9) => 
                           IMM_out_9_port, Y(8) => IMM_out_8_port, Y(7) => 
                           IMM_out_7_port, Y(6) => IMM_out_6_port, Y(5) => 
                           IMM_out_5_port, Y(4) => IMM_out_4_port, Y(3) => 
                           IMM_out_3_port, Y(2) => IMM_out_2_port, Y(1) => 
                           IMM_out_1_port, Y(0) => IMM_out_0_port);
   BHTMUX : MUX2to1_NBIT32_7 port map( A(31) => PC2_out_31_port, A(30) => 
                           PC2_out_30_port, A(29) => PC2_out_29_port, A(28) => 
                           PC2_out_28_port, A(27) => PC2_out_27_port, A(26) => 
                           PC2_out_26_port, A(25) => PC2_out_25_port, A(24) => 
                           PC2_out_24_port, A(23) => PC2_out_23_port, A(22) => 
                           PC2_out_22_port, A(21) => PC2_out_21_port, A(20) => 
                           PC2_out_20_port, A(19) => PC2_out_19_port, A(18) => 
                           PC2_out_18_port, A(17) => PC2_out_17_port, A(16) => 
                           PC2_out_16_port, A(15) => PC2_out_15_port, A(14) => 
                           PC2_out_14_port, A(13) => PC2_out_13_port, A(12) => 
                           PC2_out_12_port, A(11) => PC2_out_11_port, A(10) => 
                           PC2_out_10_port, A(9) => PC2_out_9_port, A(8) => 
                           PC2_out_8_port, A(7) => PC2_out_7_port, A(6) => 
                           PC2_out_6_port, A(5) => PC2_out_5_port, A(4) => 
                           PC2_out_4_port, A(3) => PC2_out_3_port, A(2) => 
                           PC2_out_2_port, A(1) => PC2_out_1_port, A(0) => 
                           PC2_out_0_port, B(31) => PC3_out_31_port, B(30) => 
                           PC3_out_30_port, B(29) => PC3_out_29_port, B(28) => 
                           PC3_out_28_port, B(27) => PC3_out_27_port, B(26) => 
                           PC3_out_26_port, B(25) => PC3_out_25_port, B(24) => 
                           PC3_out_24_port, B(23) => PC3_out_23_port, B(22) => 
                           PC3_out_22_port, B(21) => PC3_out_21_port, B(20) => 
                           PC3_out_20_port, B(19) => PC3_out_19_port, B(18) => 
                           PC3_out_18_port, B(17) => PC3_out_17_port, B(16) => 
                           PC3_out_16_port, B(15) => PC3_out_15_port, B(14) => 
                           PC3_out_14_port, B(13) => PC3_out_13_port, B(12) => 
                           PC3_out_12_port, B(11) => PC3_out_11_port, B(10) => 
                           PC3_out_10_port, B(9) => PC3_out_9_port, B(8) => 
                           PC3_out_8_port, B(7) => PC3_out_7_port, B(6) => 
                           PC3_out_6_port, B(5) => PC3_out_5_port, B(4) => 
                           PC3_out_4_port, B(3) => PC3_out_3_port, B(2) => 
                           PC3_out_2_port, B(1) => PC3_out_1_port, B(0) => 
                           PC3_out_0_port, SEL => BPR_EN2, Y(31) => 
                           BHT_in_31_port, Y(30) => BHT_in_30_port, Y(29) => 
                           BHT_in_29_port, Y(28) => BHT_in_28_port, Y(27) => 
                           BHT_in_27_port, Y(26) => BHT_in_26_port, Y(25) => 
                           BHT_in_25_port, Y(24) => BHT_in_24_port, Y(23) => 
                           BHT_in_23_port, Y(22) => BHT_in_22_port, Y(21) => 
                           BHT_in_21_port, Y(20) => BHT_in_20_port, Y(19) => 
                           BHT_in_19_port, Y(18) => BHT_in_18_port, Y(17) => 
                           BHT_in_17_port, Y(16) => BHT_in_16_port, Y(15) => 
                           BHT_in_15_port, Y(14) => BHT_in_14_port, Y(13) => 
                           BHT_in_13_port, Y(12) => BHT_in_12_port, Y(11) => 
                           BHT_in_11_port, Y(10) => BHT_in_10_port, Y(9) => 
                           BHT_in_9_port, Y(8) => BHT_in_8_port, Y(7) => 
                           BHT_in_7_port, Y(6) => BHT_in_6_port, Y(5) => 
                           BHT_in_5_port, Y(4) => BHT_in_4_port, Y(3) => 
                           BHT_in_3_port, Y(2) => BHT_in_2_port, Y(1) => 
                           BHT_in_1_port, Y(0) => BHT_in_0_port);
   RegAMUX : MUX2to1_NBIT32_6 port map( A(31) => FWDA_OUT_31_port, A(30) => 
                           FWDA_OUT_30_port, A(29) => FWDA_OUT_29_port, A(28) 
                           => FWDA_OUT_28_port, A(27) => FWDA_OUT_27_port, 
                           A(26) => FWDA_OUT_26_port, A(25) => FWDA_OUT_25_port
                           , A(24) => FWDA_OUT_24_port, A(23) => 
                           FWDA_OUT_23_port, A(22) => FWDA_OUT_22_port, A(21) 
                           => FWDA_OUT_21_port, A(20) => FWDA_OUT_20_port, 
                           A(19) => FWDA_OUT_19_port, A(18) => FWDA_OUT_18_port
                           , A(17) => FWDA_OUT_17_port, A(16) => 
                           FWDA_OUT_16_port, A(15) => FWDA_OUT_15_port, A(14) 
                           => FWDA_OUT_14_port, A(13) => FWDA_OUT_13_port, 
                           A(12) => FWDA_OUT_12_port, A(11) => FWDA_OUT_11_port
                           , A(10) => FWDA_OUT_10_port, A(9) => FWDA_OUT_9_port
                           , A(8) => FWDA_OUT_8_port, A(7) => FWDA_OUT_7_port, 
                           A(6) => FWDA_OUT_6_port, A(5) => FWDA_OUT_5_port, 
                           A(4) => FWDA_OUT_4_port, A(3) => FWDA_OUT_3_port, 
                           A(2) => FWDA_OUT_2_port, A(1) => FWDA_OUT_1_port, 
                           A(0) => FWDA_OUT_0_port, B(31) => X_Logic0_port, 
                           B(30) => X_Logic0_port, B(29) => X_Logic0_port, 
                           B(28) => X_Logic0_port, B(27) => X_Logic0_port, 
                           B(26) => X_Logic0_port, B(25) => X_Logic0_port, 
                           B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
                           B(22) => X_Logic0_port, B(21) => X_Logic0_port, 
                           B(20) => X_Logic0_port, B(19) => X_Logic0_port, 
                           B(18) => X_Logic0_port, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => X_Logic0_port, 
                           B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
                           B(12) => X_Logic0_port, B(11) => X_Logic0_port, 
                           B(10) => X_Logic0_port, B(9) => X_Logic0_port, B(8) 
                           => X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => ALUA_SEL, Y(31) => 
                           A_in_31_port, Y(30) => A_in_30_port, Y(29) => 
                           A_in_29_port, Y(28) => A_in_28_port, Y(27) => 
                           A_in_27_port, Y(26) => A_in_26_port, Y(25) => 
                           A_in_25_port, Y(24) => A_in_24_port, Y(23) => 
                           A_in_23_port, Y(22) => A_in_22_port, Y(21) => 
                           A_in_21_port, Y(20) => A_in_20_port, Y(19) => 
                           A_in_19_port, Y(18) => A_in_18_port, Y(17) => 
                           A_in_17_port, Y(16) => A_in_16_port, Y(15) => 
                           A_in_15_port, Y(14) => A_in_14_port, Y(13) => 
                           A_in_13_port, Y(12) => A_in_12_port, Y(11) => 
                           A_in_11_port, Y(10) => A_in_10_port, Y(9) => 
                           A_in_9_port, Y(8) => A_in_8_port, Y(7) => 
                           A_in_7_port, Y(6) => A_in_6_port, Y(5) => 
                           A_in_5_port, Y(4) => A_in_4_port, Y(3) => 
                           A_in_3_port, Y(2) => A_in_2_port, Y(1) => 
                           A_in_1_port, Y(0) => A_in_0_port);
   RegBMUX : MUX2to1_NBIT32_5 port map( A(31) => FWDB_OUT_31_port, A(30) => 
                           FWDB_OUT_30_port, A(29) => FWDB_OUT_29_port, A(28) 
                           => FWDB_OUT_28_port, A(27) => FWDB_OUT_27_port, 
                           A(26) => FWDB_OUT_26_port, A(25) => FWDB_OUT_25_port
                           , A(24) => FWDB_OUT_24_port, A(23) => 
                           FWDB_OUT_23_port, A(22) => FWDB_OUT_22_port, A(21) 
                           => FWDB_OUT_21_port, A(20) => FWDB_OUT_20_port, 
                           A(19) => FWDB_OUT_19_port, A(18) => FWDB_OUT_18_port
                           , A(17) => FWDB_OUT_17_port, A(16) => 
                           FWDB_OUT_16_port, A(15) => FWDB_OUT_15_port, A(14) 
                           => FWDB_OUT_14_port, A(13) => FWDB_OUT_13_port, 
                           A(12) => FWDB_OUT_12_port, A(11) => FWDB_OUT_11_port
                           , A(10) => FWDB_OUT_10_port, A(9) => FWDB_OUT_9_port
                           , A(8) => FWDB_OUT_8_port, A(7) => FWDB_OUT_7_port, 
                           A(6) => FWDB_OUT_6_port, A(5) => FWDB_OUT_5_port, 
                           A(4) => FWDB_OUT_4_port, A(3) => FWDB_OUT_3_port, 
                           A(2) => FWDB_OUT_2_port, A(1) => FWDB_OUT_1_port, 
                           A(0) => FWDB_OUT_0_port, B(31) => RIMM_out_31_port, 
                           B(30) => RIMM_out_30_port, B(29) => RIMM_out_29_port
                           , B(28) => RIMM_out_28_port, B(27) => 
                           RIMM_out_27_port, B(26) => RIMM_out_26_port, B(25) 
                           => RIMM_out_25_port, B(24) => RIMM_out_24_port, 
                           B(23) => RIMM_out_23_port, B(22) => RIMM_out_22_port
                           , B(21) => RIMM_out_21_port, B(20) => 
                           RIMM_out_20_port, B(19) => RIMM_out_19_port, B(18) 
                           => RIMM_out_18_port, B(17) => RIMM_out_17_port, 
                           B(16) => RIMM_out_16_port, B(15) => RIMM_out_15_port
                           , B(14) => RIMM_out_14_port, B(13) => 
                           RIMM_out_13_port, B(12) => RIMM_out_12_port, B(11) 
                           => RIMM_out_11_port, B(10) => RIMM_out_10_port, B(9)
                           => RIMM_out_9_port, B(8) => RIMM_out_8_port, B(7) =>
                           RIMM_out_7_port, B(6) => RIMM_out_6_port, B(5) => 
                           RIMM_out_5_port, B(4) => RIMM_out_4_port, B(3) => 
                           RIMM_out_3_port, B(2) => RIMM_out_2_port, B(1) => 
                           RIMM_out_1_port, B(0) => RIMM_out_0_port, SEL => 
                           ALUB_SEL, Y(31) => B_in_31_port, Y(30) => 
                           B_in_30_port, Y(29) => B_in_29_port, Y(28) => 
                           B_in_28_port, Y(27) => B_in_27_port, Y(26) => 
                           B_in_26_port, Y(25) => B_in_25_port, Y(24) => 
                           B_in_24_port, Y(23) => B_in_23_port, Y(22) => 
                           B_in_22_port, Y(21) => B_in_21_port, Y(20) => 
                           B_in_20_port, Y(19) => B_in_19_port, Y(18) => 
                           B_in_18_port, Y(17) => B_in_17_port, Y(16) => 
                           B_in_16_port, Y(15) => B_in_15_port, Y(14) => 
                           B_in_14_port, Y(13) => B_in_13_port, Y(12) => 
                           B_in_12_port, Y(11) => B_in_11_port, Y(10) => 
                           B_in_10_port, Y(9) => B_in_9_port, Y(8) => 
                           B_in_8_port, Y(7) => B_in_7_port, Y(6) => 
                           B_in_6_port, Y(5) => B_in_5_port, Y(4) => 
                           B_in_4_port, Y(3) => B_in_3_port, Y(2) => 
                           B_in_2_port, Y(1) => B_in_1_port, Y(0) => 
                           B_in_0_port);
   FWDA_MUX : MUX3to1_NBIT32_3 port map( A(31) => RA_out_31_port, A(30) => 
                           RA_out_30_port, A(29) => RA_out_29_port, A(28) => 
                           RA_out_28_port, A(27) => RA_out_27_port, A(26) => 
                           RA_out_26_port, A(25) => RA_out_25_port, A(24) => 
                           RA_out_24_port, A(23) => RA_out_23_port, A(22) => 
                           RA_out_22_port, A(21) => RA_out_21_port, A(20) => 
                           RA_out_20_port, A(19) => RA_out_19_port, A(18) => 
                           RA_out_18_port, A(17) => RA_out_17_port, A(16) => 
                           RA_out_16_port, A(15) => RA_out_15_port, A(14) => 
                           RA_out_14_port, A(13) => RA_out_13_port, A(12) => 
                           RA_out_12_port, A(11) => RA_out_11_port, A(10) => 
                           RA_out_10_port, A(9) => RA_out_9_port, A(8) => 
                           RA_out_8_port, A(7) => RA_out_7_port, A(6) => 
                           RA_out_6_port, A(5) => RA_out_5_port, A(4) => 
                           RA_out_4_port, A(3) => RA_out_3_port, A(2) => 
                           RA_out_2_port, A(1) => RA_out_1_port, A(0) => 
                           RA_out_0_port, B(31) => DATA_ADDR_31_port, B(30) => 
                           DATA_ADDR_30_port, B(29) => DATA_ADDR_29_port, B(28)
                           => DATA_ADDR_28_port, B(27) => DATA_ADDR_27_port, 
                           B(26) => DATA_ADDR_26_port, B(25) => 
                           DATA_ADDR_25_port, B(24) => DATA_ADDR_24_port, B(23)
                           => DATA_ADDR_23_port, B(22) => DATA_ADDR_22_port, 
                           B(21) => DATA_ADDR_21_port, B(20) => 
                           DATA_ADDR_20_port, B(19) => DATA_ADDR_19_port, B(18)
                           => DATA_ADDR_18_port, B(17) => DATA_ADDR_17_port, 
                           B(16) => DATA_ADDR_16_port, B(15) => 
                           DATA_ADDR_15_port, B(14) => DATA_ADDR_14_port, B(13)
                           => DATA_ADDR_13_port, B(12) => DATA_ADDR_12_port, 
                           B(11) => DATA_ADDR_11_port, B(10) => 
                           DATA_ADDR_10_port, B(9) => DATA_ADDR_9_port, B(8) =>
                           DATA_ADDR_8_port, B(7) => DATA_ADDR_7_port, B(6) => 
                           DATA_ADDR_6_port, B(5) => DATA_ADDR_5_port, B(4) => 
                           DATA_ADDR_4_port, B(3) => DATA_ADDR_3_port, B(2) => 
                           DATA_ADDR_2_port, B(1) => DATA_ADDR_1_port, B(0) => 
                           DATA_ADDR_0_port, C(31) => WB_in_31_port, C(30) => 
                           WB_in_30_port, C(29) => WB_in_29_port, C(28) => 
                           WB_in_28_port, C(27) => WB_in_27_port, C(26) => 
                           WB_in_26_port, C(25) => WB_in_25_port, C(24) => 
                           WB_in_24_port, C(23) => WB_in_23_port, C(22) => 
                           WB_in_22_port, C(21) => WB_in_21_port, C(20) => 
                           WB_in_20_port, C(19) => WB_in_19_port, C(18) => 
                           WB_in_18_port, C(17) => WB_in_17_port, C(16) => 
                           WB_in_16_port, C(15) => WB_in_15_port, C(14) => 
                           WB_in_14_port, C(13) => WB_in_13_port, C(12) => 
                           WB_in_12_port, C(11) => WB_in_11_port, C(10) => 
                           WB_in_10_port, C(9) => WB_in_9_port, C(8) => 
                           WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => FWDA_SEL_1_port, SEL(0) => 
                           FWDA_SEL_0_port, Y(31) => FWDA_OUT_31_port, Y(30) =>
                           FWDA_OUT_30_port, Y(29) => FWDA_OUT_29_port, Y(28) 
                           => FWDA_OUT_28_port, Y(27) => FWDA_OUT_27_port, 
                           Y(26) => FWDA_OUT_26_port, Y(25) => FWDA_OUT_25_port
                           , Y(24) => FWDA_OUT_24_port, Y(23) => 
                           FWDA_OUT_23_port, Y(22) => FWDA_OUT_22_port, Y(21) 
                           => FWDA_OUT_21_port, Y(20) => FWDA_OUT_20_port, 
                           Y(19) => FWDA_OUT_19_port, Y(18) => FWDA_OUT_18_port
                           , Y(17) => FWDA_OUT_17_port, Y(16) => 
                           FWDA_OUT_16_port, Y(15) => FWDA_OUT_15_port, Y(14) 
                           => FWDA_OUT_14_port, Y(13) => FWDA_OUT_13_port, 
                           Y(12) => FWDA_OUT_12_port, Y(11) => FWDA_OUT_11_port
                           , Y(10) => FWDA_OUT_10_port, Y(9) => FWDA_OUT_9_port
                           , Y(8) => FWDA_OUT_8_port, Y(7) => FWDA_OUT_7_port, 
                           Y(6) => FWDA_OUT_6_port, Y(5) => FWDA_OUT_5_port, 
                           Y(4) => FWDA_OUT_4_port, Y(3) => FWDA_OUT_3_port, 
                           Y(2) => FWDA_OUT_2_port, Y(1) => FWDA_OUT_1_port, 
                           Y(0) => FWDA_OUT_0_port);
   FWDB_MUX : MUX3to1_NBIT32_2 port map( A(31) => RB_out_31_port, A(30) => 
                           RB_out_30_port, A(29) => RB_out_29_port, A(28) => 
                           RB_out_28_port, A(27) => RB_out_27_port, A(26) => 
                           RB_out_26_port, A(25) => RB_out_25_port, A(24) => 
                           RB_out_24_port, A(23) => RB_out_23_port, A(22) => 
                           RB_out_22_port, A(21) => RB_out_21_port, A(20) => 
                           RB_out_20_port, A(19) => RB_out_19_port, A(18) => 
                           RB_out_18_port, A(17) => RB_out_17_port, A(16) => 
                           RB_out_16_port, A(15) => RB_out_15_port, A(14) => 
                           RB_out_14_port, A(13) => RB_out_13_port, A(12) => 
                           RB_out_12_port, A(11) => RB_out_11_port, A(10) => 
                           RB_out_10_port, A(9) => RB_out_9_port, A(8) => 
                           RB_out_8_port, A(7) => RB_out_7_port, A(6) => 
                           RB_out_6_port, A(5) => RB_out_5_port, A(4) => 
                           RB_out_4_port, A(3) => RB_out_3_port, A(2) => 
                           RB_out_2_port, A(1) => RB_out_1_port, A(0) => 
                           RB_out_0_port, B(31) => DATA_ADDR_31_port, B(30) => 
                           DATA_ADDR_30_port, B(29) => DATA_ADDR_29_port, B(28)
                           => DATA_ADDR_28_port, B(27) => DATA_ADDR_27_port, 
                           B(26) => DATA_ADDR_26_port, B(25) => 
                           DATA_ADDR_25_port, B(24) => DATA_ADDR_24_port, B(23)
                           => DATA_ADDR_23_port, B(22) => DATA_ADDR_22_port, 
                           B(21) => DATA_ADDR_21_port, B(20) => 
                           DATA_ADDR_20_port, B(19) => DATA_ADDR_19_port, B(18)
                           => DATA_ADDR_18_port, B(17) => DATA_ADDR_17_port, 
                           B(16) => DATA_ADDR_16_port, B(15) => 
                           DATA_ADDR_15_port, B(14) => DATA_ADDR_14_port, B(13)
                           => DATA_ADDR_13_port, B(12) => DATA_ADDR_12_port, 
                           B(11) => DATA_ADDR_11_port, B(10) => 
                           DATA_ADDR_10_port, B(9) => DATA_ADDR_9_port, B(8) =>
                           DATA_ADDR_8_port, B(7) => DATA_ADDR_7_port, B(6) => 
                           DATA_ADDR_6_port, B(5) => DATA_ADDR_5_port, B(4) => 
                           DATA_ADDR_4_port, B(3) => DATA_ADDR_3_port, B(2) => 
                           DATA_ADDR_2_port, B(1) => DATA_ADDR_1_port, B(0) => 
                           DATA_ADDR_0_port, C(31) => WB_in_31_port, C(30) => 
                           WB_in_30_port, C(29) => WB_in_29_port, C(28) => 
                           WB_in_28_port, C(27) => WB_in_27_port, C(26) => 
                           WB_in_26_port, C(25) => WB_in_25_port, C(24) => 
                           WB_in_24_port, C(23) => WB_in_23_port, C(22) => 
                           WB_in_22_port, C(21) => WB_in_21_port, C(20) => 
                           WB_in_20_port, C(19) => WB_in_19_port, C(18) => 
                           WB_in_18_port, C(17) => WB_in_17_port, C(16) => 
                           WB_in_16_port, C(15) => WB_in_15_port, C(14) => 
                           WB_in_14_port, C(13) => WB_in_13_port, C(12) => 
                           WB_in_12_port, C(11) => WB_in_11_port, C(10) => 
                           WB_in_10_port, C(9) => WB_in_9_port, C(8) => 
                           WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => FWDB_SEL_1_port, SEL(0) => 
                           FWDB_SEL_0_port, Y(31) => FWDB_OUT_31_port, Y(30) =>
                           FWDB_OUT_30_port, Y(29) => FWDB_OUT_29_port, Y(28) 
                           => FWDB_OUT_28_port, Y(27) => FWDB_OUT_27_port, 
                           Y(26) => FWDB_OUT_26_port, Y(25) => FWDB_OUT_25_port
                           , Y(24) => FWDB_OUT_24_port, Y(23) => 
                           FWDB_OUT_23_port, Y(22) => FWDB_OUT_22_port, Y(21) 
                           => FWDB_OUT_21_port, Y(20) => FWDB_OUT_20_port, 
                           Y(19) => FWDB_OUT_19_port, Y(18) => FWDB_OUT_18_port
                           , Y(17) => FWDB_OUT_17_port, Y(16) => 
                           FWDB_OUT_16_port, Y(15) => FWDB_OUT_15_port, Y(14) 
                           => FWDB_OUT_14_port, Y(13) => FWDB_OUT_13_port, 
                           Y(12) => FWDB_OUT_12_port, Y(11) => FWDB_OUT_11_port
                           , Y(10) => FWDB_OUT_10_port, Y(9) => FWDB_OUT_9_port
                           , Y(8) => FWDB_OUT_8_port, Y(7) => FWDB_OUT_7_port, 
                           Y(6) => FWDB_OUT_6_port, Y(5) => FWDB_OUT_5_port, 
                           Y(4) => FWDB_OUT_4_port, Y(3) => FWDB_OUT_3_port, 
                           Y(2) => FWDB_OUT_2_port, Y(1) => FWDB_OUT_1_port, 
                           Y(0) => FWDB_OUT_0_port);
   ZDU_MUX : MUX3to1_NBIT32_1 port map( A(31) => RA_out_31_port, A(30) => 
                           RA_out_30_port, A(29) => RA_out_29_port, A(28) => 
                           RA_out_28_port, A(27) => RA_out_27_port, A(26) => 
                           RA_out_26_port, A(25) => RA_out_25_port, A(24) => 
                           RA_out_24_port, A(23) => RA_out_23_port, A(22) => 
                           RA_out_22_port, A(21) => RA_out_21_port, A(20) => 
                           RA_out_20_port, A(19) => RA_out_19_port, A(18) => 
                           RA_out_18_port, A(17) => RA_out_17_port, A(16) => 
                           RA_out_16_port, A(15) => RA_out_15_port, A(14) => 
                           RA_out_14_port, A(13) => RA_out_13_port, A(12) => 
                           RA_out_12_port, A(11) => RA_out_11_port, A(10) => 
                           RA_out_10_port, A(9) => RA_out_9_port, A(8) => 
                           RA_out_8_port, A(7) => RA_out_7_port, A(6) => 
                           RA_out_6_port, A(5) => RA_out_5_port, A(4) => 
                           RA_out_4_port, A(3) => RA_out_3_port, A(2) => 
                           RA_out_2_port, A(1) => RA_out_1_port, A(0) => 
                           RA_out_0_port, B(31) => CWB_MUX2_out_31_port, B(30) 
                           => CWB_MUX2_out_30_port, B(29) => 
                           CWB_MUX2_out_29_port, B(28) => CWB_MUX2_out_28_port,
                           B(27) => CWB_MUX2_out_27_port, B(26) => 
                           CWB_MUX2_out_26_port, B(25) => CWB_MUX2_out_25_port,
                           B(24) => CWB_MUX2_out_24_port, B(23) => 
                           CWB_MUX2_out_23_port, B(22) => CWB_MUX2_out_22_port,
                           B(21) => CWB_MUX2_out_21_port, B(20) => 
                           CWB_MUX2_out_20_port, B(19) => CWB_MUX2_out_19_port,
                           B(18) => CWB_MUX2_out_18_port, B(17) => 
                           CWB_MUX2_out_17_port, B(16) => CWB_MUX2_out_16_port,
                           B(15) => CWB_MUX2_out_15_port, B(14) => 
                           CWB_MUX2_out_14_port, B(13) => CWB_MUX2_out_13_port,
                           B(12) => CWB_MUX2_out_12_port, B(11) => 
                           CWB_MUX2_out_11_port, B(10) => CWB_MUX2_out_10_port,
                           B(9) => CWB_MUX2_out_9_port, B(8) => 
                           CWB_MUX2_out_8_port, B(7) => CWB_MUX2_out_7_port, 
                           B(6) => CWB_MUX2_out_6_port, B(5) => 
                           CWB_MUX2_out_5_port, B(4) => CWB_MUX2_out_4_port, 
                           B(3) => CWB_MUX2_out_3_port, B(2) => 
                           CWB_MUX2_out_2_port, B(1) => CWB_MUX2_out_1_port, 
                           B(0) => CWB_MUX2_out_0_port, C(31) => WB_in_31_port,
                           C(30) => WB_in_30_port, C(29) => WB_in_29_port, 
                           C(28) => WB_in_28_port, C(27) => WB_in_27_port, 
                           C(26) => WB_in_26_port, C(25) => WB_in_25_port, 
                           C(24) => WB_in_24_port, C(23) => WB_in_23_port, 
                           C(22) => WB_in_22_port, C(21) => WB_in_21_port, 
                           C(20) => WB_in_20_port, C(19) => WB_in_19_port, 
                           C(18) => WB_in_18_port, C(17) => WB_in_17_port, 
                           C(16) => WB_in_16_port, C(15) => WB_in_15_port, 
                           C(14) => WB_in_14_port, C(13) => WB_in_13_port, 
                           C(12) => WB_in_12_port, C(11) => WB_in_11_port, 
                           C(10) => WB_in_10_port, C(9) => WB_in_9_port, C(8) 
                           => WB_in_8_port, C(7) => WB_in_7_port, C(6) => 
                           WB_in_6_port, C(5) => WB_in_5_port, C(4) => 
                           WB_in_4_port, C(3) => WB_in_3_port, C(2) => 
                           WB_in_2_port, C(1) => WB_in_1_port, C(0) => 
                           WB_in_0_port, SEL(1) => ZDU_SEL_1_port, SEL(0) => 
                           ZDU_SEL_0_port, Y(31) => n_1662, Y(30) => 
                           ZDU_MUX_out_30_port, Y(29) => ZDU_MUX_out_29_port, 
                           Y(28) => ZDU_MUX_out_28_port, Y(27) => 
                           ZDU_MUX_out_27_port, Y(26) => ZDU_MUX_out_26_port, 
                           Y(25) => ZDU_MUX_out_25_port, Y(24) => 
                           ZDU_MUX_out_24_port, Y(23) => ZDU_MUX_out_23_port, 
                           Y(22) => ZDU_MUX_out_22_port, Y(21) => 
                           ZDU_MUX_out_21_port, Y(20) => ZDU_MUX_out_20_port, 
                           Y(19) => ZDU_MUX_out_19_port, Y(18) => 
                           ZDU_MUX_out_18_port, Y(17) => ZDU_MUX_out_17_port, 
                           Y(16) => ZDU_MUX_out_16_port, Y(15) => 
                           ZDU_MUX_out_15_port, Y(14) => ZDU_MUX_out_14_port, 
                           Y(13) => ZDU_MUX_out_13_port, Y(12) => 
                           ZDU_MUX_out_12_port, Y(11) => ZDU_MUX_out_11_port, 
                           Y(10) => ZDU_MUX_out_10_port, Y(9) => 
                           ZDU_MUX_out_9_port, Y(8) => ZDU_MUX_out_8_port, Y(7)
                           => ZDU_MUX_out_7_port, Y(6) => ZDU_MUX_out_6_port, 
                           Y(5) => ZDU_MUX_out_5_port, Y(4) => 
                           ZDU_MUX_out_4_port, Y(3) => ZDU_MUX_out_3_port, Y(2)
                           => ZDU_MUX_out_2_port, Y(1) => ZDU_MUX_out_1_port, 
                           Y(0) => ZDU_MUX_out_0_port);
   MEMDATAMUX : MUX2to1_NBIT32_4 port map( A(31) => ALR2_out_31_port, A(30) => 
                           ALR2_out_30_port, A(29) => ALR2_out_29_port, A(28) 
                           => ALR2_out_28_port, A(27) => ALR2_out_27_port, 
                           A(26) => ALR2_out_26_port, A(25) => ALR2_out_25_port
                           , A(24) => ALR2_out_24_port, A(23) => 
                           ALR2_out_23_port, A(22) => ALR2_out_22_port, A(21) 
                           => ALR2_out_21_port, A(20) => ALR2_out_20_port, 
                           A(19) => ALR2_out_19_port, A(18) => ALR2_out_18_port
                           , A(17) => ALR2_out_17_port, A(16) => 
                           ALR2_out_16_port, A(15) => ALR2_out_15_port, A(14) 
                           => ALR2_out_14_port, A(13) => ALR2_out_13_port, 
                           A(12) => ALR2_out_12_port, A(11) => ALR2_out_11_port
                           , A(10) => ALR2_out_10_port, A(9) => ALR2_out_9_port
                           , A(8) => ALR2_out_8_port, A(7) => ALR2_out_7_port, 
                           A(6) => ALR2_out_6_port, A(5) => ALR2_out_5_port, 
                           A(4) => ALR2_out_4_port, A(3) => ALR2_out_3_port, 
                           A(2) => ALR2_out_2_port, A(1) => ALR2_out_1_port, 
                           A(0) => ALR2_out_0_port, B(31) => B2_MUX_out_31_port
                           , B(30) => B2_MUX_out_30_port, B(29) => 
                           B2_MUX_out_29_port, B(28) => B2_MUX_out_28_port, 
                           B(27) => B2_MUX_out_27_port, B(26) => 
                           B2_MUX_out_26_port, B(25) => B2_MUX_out_25_port, 
                           B(24) => B2_MUX_out_24_port, B(23) => 
                           B2_MUX_out_23_port, B(22) => B2_MUX_out_22_port, 
                           B(21) => B2_MUX_out_21_port, B(20) => 
                           B2_MUX_out_20_port, B(19) => B2_MUX_out_19_port, 
                           B(18) => B2_MUX_out_18_port, B(17) => 
                           B2_MUX_out_17_port, B(16) => B2_MUX_out_16_port, 
                           B(15) => B2_MUX_out_15_port, B(14) => 
                           B2_MUX_out_14_port, B(13) => B2_MUX_out_13_port, 
                           B(12) => B2_MUX_out_12_port, B(11) => 
                           B2_MUX_out_11_port, B(10) => B2_MUX_out_10_port, 
                           B(9) => B2_MUX_out_9_port, B(8) => B2_MUX_out_8_port
                           , B(7) => B2_MUX_out_7_port, B(6) => 
                           B2_MUX_out_6_port, B(5) => B2_MUX_out_5_port, B(4) 
                           => B2_MUX_out_4_port, B(3) => B2_MUX_out_3_port, 
                           B(2) => B2_MUX_out_2_port, B(1) => B2_MUX_out_1_port
                           , B(0) => B2_MUX_out_0_port, SEL => MEM_DATA_SEL, 
                           Y(31) => DATA_OUT(31), Y(30) => DATA_OUT(30), Y(29) 
                           => DATA_OUT(29), Y(28) => DATA_OUT(28), Y(27) => 
                           DATA_OUT(27), Y(26) => DATA_OUT(26), Y(25) => 
                           DATA_OUT(25), Y(24) => DATA_OUT(24), Y(23) => 
                           DATA_OUT(23), Y(22) => DATA_OUT(22), Y(21) => 
                           DATA_OUT(21), Y(20) => DATA_OUT(20), Y(19) => 
                           DATA_OUT(19), Y(18) => DATA_OUT(18), Y(17) => 
                           DATA_OUT(17), Y(16) => DATA_OUT(16), Y(15) => 
                           DATA_OUT(15), Y(14) => DATA_OUT(14), Y(13) => 
                           DATA_OUT(13), Y(12) => DATA_OUT(12), Y(11) => 
                           DATA_OUT(11), Y(10) => DATA_OUT(10), Y(9) => 
                           DATA_OUT(9), Y(8) => DATA_OUT(8), Y(7) => 
                           DATA_OUT(7), Y(6) => DATA_OUT(6), Y(5) => 
                           DATA_OUT(5), Y(4) => DATA_OUT(4), Y(3) => 
                           DATA_OUT(3), Y(2) => DATA_OUT(2), Y(1) => 
                           DATA_OUT(1), Y(0) => DATA_OUT(0));
   LMDMUX : MUX5to1_NBIT32_0 port map( A(31) => n25, A(30) => DATA_IN(6), A(29)
                           => DATA_IN(5), A(28) => DATA_IN(4), A(27) => 
                           DATA_IN(3), A(26) => DATA_IN(2), A(25) => DATA_IN(1)
                           , A(24) => DATA_IN(0), A(23) => DATA_IN(15), A(22) 
                           => DATA_IN(14), A(21) => DATA_IN(13), A(20) => 
                           DATA_IN(12), A(19) => DATA_IN(11), A(18) => 
                           DATA_IN(10), A(17) => DATA_IN(9), A(16) => 
                           DATA_IN(8), A(15) => DATA_IN(23), A(14) => 
                           DATA_IN(22), A(13) => DATA_IN(21), A(12) => 
                           DATA_IN(20), A(11) => DATA_IN(19), A(10) => 
                           DATA_IN(18), A(9) => DATA_IN(17), A(8) => 
                           DATA_IN(16), A(7) => DATA_IN(31), A(6) => 
                           DATA_IN(30), A(5) => DATA_IN(29), A(4) => 
                           DATA_IN(28), A(3) => DATA_IN(27), A(2) => 
                           DATA_IN(26), A(1) => DATA_IN(25), A(0) => 
                           DATA_IN(24), B(31) => n23, B(30) => n23, B(29) => 
                           n23, B(28) => n23, B(27) => n23, B(26) => n23, B(25)
                           => n23, B(24) => n23, B(23) => n23, B(22) => n23, 
                           B(21) => n23, B(20) => n24, B(19) => n24, B(18) => 
                           n24, B(17) => n24, B(16) => n24, B(15) => n24, B(14)
                           => n24, B(13) => n24, B(12) => n24, B(11) => n24, 
                           B(10) => n24, B(9) => n24, B(8) => n25, B(7) => n25,
                           B(6) => DATA_IN(6), B(5) => DATA_IN(5), B(4) => 
                           DATA_IN(4), B(3) => DATA_IN(3), B(2) => DATA_IN(2), 
                           B(1) => DATA_IN(1), B(0) => DATA_IN(0), C(31) => 
                           X_Logic0_port, C(30) => X_Logic0_port, C(29) => 
                           X_Logic0_port, C(28) => X_Logic0_port, C(27) => 
                           X_Logic0_port, C(26) => X_Logic0_port, C(25) => 
                           X_Logic0_port, C(24) => X_Logic0_port, C(23) => 
                           X_Logic0_port, C(22) => X_Logic0_port, C(21) => 
                           X_Logic0_port, C(20) => X_Logic0_port, C(19) => 
                           X_Logic0_port, C(18) => X_Logic0_port, C(17) => 
                           X_Logic0_port, C(16) => X_Logic0_port, C(15) => 
                           X_Logic0_port, C(14) => X_Logic0_port, C(13) => 
                           X_Logic0_port, C(12) => X_Logic0_port, C(11) => 
                           X_Logic0_port, C(10) => X_Logic0_port, C(9) => 
                           X_Logic0_port, C(8) => X_Logic0_port, C(7) => n23, 
                           C(6) => DATA_IN(6), C(5) => DATA_IN(5), C(4) => 
                           DATA_IN(4), C(3) => DATA_IN(3), C(2) => DATA_IN(2), 
                           C(1) => DATA_IN(1), C(0) => DATA_IN(0), D(31) => n25
                           , D(30) => n25, D(29) => n25, D(28) => n25, D(27) =>
                           n25, D(26) => n25, D(25) => n25, D(24) => n26, D(23)
                           => n25, D(22) => n26, D(21) => n26, D(20) => n26, 
                           D(19) => n26, D(18) => n26, D(17) => n26, D(16) => 
                           n26, D(15) => n26, D(14) => DATA_IN(6), D(13) => 
                           DATA_IN(5), D(12) => DATA_IN(4), D(11) => DATA_IN(3)
                           , D(10) => DATA_IN(2), D(9) => DATA_IN(1), D(8) => 
                           DATA_IN(0), D(7) => DATA_IN(15), D(6) => DATA_IN(14)
                           , D(5) => DATA_IN(13), D(4) => DATA_IN(12), D(3) => 
                           DATA_IN(11), D(2) => DATA_IN(10), D(1) => DATA_IN(9)
                           , D(0) => DATA_IN(8), E(31) => X_Logic0_port, E(30) 
                           => X_Logic0_port, E(29) => X_Logic0_port, E(28) => 
                           X_Logic0_port, E(27) => X_Logic0_port, E(26) => 
                           X_Logic0_port, E(25) => X_Logic0_port, E(24) => 
                           X_Logic0_port, E(23) => X_Logic0_port, E(22) => 
                           X_Logic0_port, E(21) => X_Logic0_port, E(20) => 
                           X_Logic0_port, E(19) => X_Logic0_port, E(18) => 
                           X_Logic0_port, E(17) => X_Logic0_port, E(16) => 
                           X_Logic0_port, E(15) => n25, E(14) => DATA_IN(6), 
                           E(13) => DATA_IN(5), E(12) => DATA_IN(4), E(11) => 
                           DATA_IN(3), E(10) => DATA_IN(2), E(9) => DATA_IN(1),
                           E(8) => DATA_IN(0), E(7) => DATA_IN(15), E(6) => 
                           DATA_IN(14), E(5) => DATA_IN(13), E(4) => 
                           DATA_IN(12), E(3) => DATA_IN(11), E(2) => 
                           DATA_IN(10), E(1) => DATA_IN(9), E(0) => DATA_IN(8),
                           SEL(2) => LD_SEL(2), SEL(1) => LD_SEL(1), SEL(0) => 
                           LD_SEL(0), Y(31) => LMD_out_31_port, Y(30) => 
                           LMD_out_30_port, Y(29) => LMD_out_29_port, Y(28) => 
                           LMD_out_28_port, Y(27) => LMD_out_27_port, Y(26) => 
                           LMD_out_26_port, Y(25) => LMD_out_25_port, Y(24) => 
                           LMD_out_24_port, Y(23) => LMD_out_23_port, Y(22) => 
                           LMD_out_22_port, Y(21) => LMD_out_21_port, Y(20) => 
                           LMD_out_20_port, Y(19) => LMD_out_19_port, Y(18) => 
                           LMD_out_18_port, Y(17) => LMD_out_17_port, Y(16) => 
                           LMD_out_16_port, Y(15) => LMD_out_15_port, Y(14) => 
                           LMD_out_14_port, Y(13) => LMD_out_13_port, Y(12) => 
                           LMD_out_12_port, Y(11) => LMD_out_11_port, Y(10) => 
                           LMD_out_10_port, Y(9) => LMD_out_9_port, Y(8) => 
                           LMD_out_8_port, Y(7) => LMD_out_7_port, Y(6) => 
                           LMD_out_6_port, Y(5) => LMD_out_5_port, Y(4) => 
                           LMD_out_4_port, Y(3) => LMD_out_3_port, Y(2) => 
                           LMD_out_2_port, Y(1) => LMD_out_1_port, Y(0) => 
                           LMD_out_0_port);
   ALR2_MUX : MUX2to1_NBIT32_3 port map( A(31) => CWB_MUX2_out_31_port, A(30) 
                           => CWB_MUX2_out_30_port, A(29) => 
                           CWB_MUX2_out_29_port, A(28) => CWB_MUX2_out_28_port,
                           A(27) => CWB_MUX2_out_27_port, A(26) => 
                           CWB_MUX2_out_26_port, A(25) => CWB_MUX2_out_25_port,
                           A(24) => CWB_MUX2_out_24_port, A(23) => 
                           CWB_MUX2_out_23_port, A(22) => CWB_MUX2_out_22_port,
                           A(21) => CWB_MUX2_out_21_port, A(20) => 
                           CWB_MUX2_out_20_port, A(19) => CWB_MUX2_out_19_port,
                           A(18) => CWB_MUX2_out_18_port, A(17) => 
                           CWB_MUX2_out_17_port, A(16) => CWB_MUX2_out_16_port,
                           A(15) => CWB_MUX2_out_15_port, A(14) => 
                           CWB_MUX2_out_14_port, A(13) => CWB_MUX2_out_13_port,
                           A(12) => CWB_MUX2_out_12_port, A(11) => 
                           CWB_MUX2_out_11_port, A(10) => CWB_MUX2_out_10_port,
                           A(9) => CWB_MUX2_out_9_port, A(8) => 
                           CWB_MUX2_out_8_port, A(7) => CWB_MUX2_out_7_port, 
                           A(6) => CWB_MUX2_out_6_port, A(5) => 
                           CWB_MUX2_out_5_port, A(4) => CWB_MUX2_out_4_port, 
                           A(3) => CWB_MUX2_out_3_port, A(2) => 
                           CWB_MUX2_out_2_port, A(1) => CWB_MUX2_out_1_port, 
                           A(0) => CWB_MUX2_out_0_port, B(31) => 
                           NPC3_out_31_port, B(30) => NPC3_out_30_port, B(29) 
                           => NPC3_out_29_port, B(28) => NPC3_out_28_port, 
                           B(27) => NPC3_out_27_port, B(26) => NPC3_out_26_port
                           , B(25) => NPC3_out_25_port, B(24) => 
                           NPC3_out_24_port, B(23) => NPC3_out_23_port, B(22) 
                           => NPC3_out_22_port, B(21) => NPC3_out_21_port, 
                           B(20) => NPC3_out_20_port, B(19) => NPC3_out_19_port
                           , B(18) => NPC3_out_18_port, B(17) => 
                           NPC3_out_17_port, B(16) => NPC3_out_16_port, B(15) 
                           => NPC3_out_15_port, B(14) => NPC3_out_14_port, 
                           B(13) => NPC3_out_13_port, B(12) => NPC3_out_12_port
                           , B(11) => NPC3_out_11_port, B(10) => 
                           NPC3_out_10_port, B(9) => NPC3_out_9_port, B(8) => 
                           NPC3_out_8_port, B(7) => NPC3_out_7_port, B(6) => 
                           NPC3_out_6_port, B(5) => NPC3_out_5_port, B(4) => 
                           NPC3_out_4_port, B(3) => NPC3_out_3_port, B(2) => 
                           NPC3_out_2_port, B(1) => NPC3_out_1_port, B(0) => 
                           NPC3_out_0_port, SEL => ALR2_SEL, Y(31) => 
                           ALR2_in_31_port, Y(30) => ALR2_in_30_port, Y(29) => 
                           ALR2_in_29_port, Y(28) => ALR2_in_28_port, Y(27) => 
                           ALR2_in_27_port, Y(26) => ALR2_in_26_port, Y(25) => 
                           ALR2_in_25_port, Y(24) => ALR2_in_24_port, Y(23) => 
                           ALR2_in_23_port, Y(22) => ALR2_in_22_port, Y(21) => 
                           ALR2_in_21_port, Y(20) => ALR2_in_20_port, Y(19) => 
                           ALR2_in_19_port, Y(18) => ALR2_in_18_port, Y(17) => 
                           ALR2_in_17_port, Y(16) => ALR2_in_16_port, Y(15) => 
                           ALR2_in_15_port, Y(14) => ALR2_in_14_port, Y(13) => 
                           ALR2_in_13_port, Y(12) => ALR2_in_12_port, Y(11) => 
                           ALR2_in_11_port, Y(10) => ALR2_in_10_port, Y(9) => 
                           ALR2_in_9_port, Y(8) => ALR2_in_8_port, Y(7) => 
                           ALR2_in_7_port, Y(6) => ALR2_in_6_port, Y(5) => 
                           ALR2_in_5_port, Y(4) => ALR2_in_4_port, Y(3) => 
                           ALR2_in_3_port, Y(2) => ALR2_in_2_port, Y(1) => 
                           ALR2_in_1_port, Y(0) => ALR2_in_0_port);
   CWB_MUX1 : MUX3to1_NBIT2 port map( A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, C(1) => CWB_out_1_port, C(0) => 
                           CWB_out_0_port, SEL(1) => CWB_MUX_SEL_1_port, SEL(0)
                           => CWB_MUX_SEL_0_port, Y(1) => CWB2_SEL_1_port, Y(0)
                           => CWB2_SEL_0_port);
   CWB_MUX2 : MUX4to1_NBIT32_0 port map( A(31) => DATA_ADDR_31_port, A(30) => 
                           DATA_ADDR_30_port, A(29) => DATA_ADDR_29_port, A(28)
                           => DATA_ADDR_28_port, A(27) => DATA_ADDR_27_port, 
                           A(26) => DATA_ADDR_26_port, A(25) => 
                           DATA_ADDR_25_port, A(24) => DATA_ADDR_24_port, A(23)
                           => DATA_ADDR_23_port, A(22) => DATA_ADDR_22_port, 
                           A(21) => DATA_ADDR_21_port, A(20) => 
                           DATA_ADDR_20_port, A(19) => DATA_ADDR_19_port, A(18)
                           => DATA_ADDR_18_port, A(17) => DATA_ADDR_17_port, 
                           A(16) => DATA_ADDR_16_port, A(15) => 
                           DATA_ADDR_15_port, A(14) => DATA_ADDR_14_port, A(13)
                           => DATA_ADDR_13_port, A(12) => DATA_ADDR_12_port, 
                           A(11) => DATA_ADDR_11_port, A(10) => 
                           DATA_ADDR_10_port, A(9) => DATA_ADDR_9_port, A(8) =>
                           DATA_ADDR_8_port, A(7) => DATA_ADDR_7_port, A(6) => 
                           DATA_ADDR_6_port, A(5) => DATA_ADDR_5_port, A(4) => 
                           DATA_ADDR_4_port, A(3) => DATA_ADDR_3_port, A(2) => 
                           DATA_ADDR_2_port, A(1) => DATA_ADDR_1_port, A(0) => 
                           DATA_ADDR_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, C(31) => X_Logic0_port, C(30) => 
                           X_Logic0_port, C(29) => X_Logic0_port, C(28) => 
                           X_Logic0_port, C(27) => X_Logic0_port, C(26) => 
                           X_Logic0_port, C(25) => X_Logic0_port, C(24) => 
                           X_Logic0_port, C(23) => X_Logic0_port, C(22) => 
                           X_Logic0_port, C(21) => X_Logic0_port, C(20) => 
                           X_Logic0_port, C(19) => X_Logic0_port, C(18) => 
                           X_Logic0_port, C(17) => X_Logic0_port, C(16) => 
                           X_Logic0_port, C(15) => X_Logic0_port, C(14) => 
                           X_Logic0_port, C(13) => X_Logic0_port, C(12) => 
                           X_Logic0_port, C(11) => X_Logic0_port, C(10) => 
                           X_Logic0_port, C(9) => X_Logic0_port, C(8) => 
                           X_Logic0_port, C(7) => X_Logic0_port, C(6) => 
                           X_Logic0_port, C(5) => X_Logic0_port, C(4) => 
                           X_Logic0_port, C(3) => X_Logic0_port, C(2) => 
                           X_Logic0_port, C(1) => X_Logic0_port, C(0) => 
                           X_Logic0_port, D(31) => DATA_ADDR_15_port, D(30) => 
                           DATA_ADDR_14_port, D(29) => DATA_ADDR_13_port, D(28)
                           => DATA_ADDR_12_port, D(27) => DATA_ADDR_11_port, 
                           D(26) => DATA_ADDR_10_port, D(25) => 
                           DATA_ADDR_9_port, D(24) => DATA_ADDR_8_port, D(23) 
                           => DATA_ADDR_7_port, D(22) => DATA_ADDR_6_port, 
                           D(21) => DATA_ADDR_5_port, D(20) => DATA_ADDR_4_port
                           , D(19) => DATA_ADDR_3_port, D(18) => 
                           DATA_ADDR_2_port, D(17) => DATA_ADDR_1_port, D(16) 
                           => DATA_ADDR_0_port, D(15) => X_Logic0_port, D(14) 
                           => X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, SEL(1) => CWB2_SEL_1_port, SEL(0) => 
                           CWB2_SEL_0_port, Y(31) => CWB_MUX2_out_31_port, 
                           Y(30) => CWB_MUX2_out_30_port, Y(29) => 
                           CWB_MUX2_out_29_port, Y(28) => CWB_MUX2_out_28_port,
                           Y(27) => CWB_MUX2_out_27_port, Y(26) => 
                           CWB_MUX2_out_26_port, Y(25) => CWB_MUX2_out_25_port,
                           Y(24) => CWB_MUX2_out_24_port, Y(23) => 
                           CWB_MUX2_out_23_port, Y(22) => CWB_MUX2_out_22_port,
                           Y(21) => CWB_MUX2_out_21_port, Y(20) => 
                           CWB_MUX2_out_20_port, Y(19) => CWB_MUX2_out_19_port,
                           Y(18) => CWB_MUX2_out_18_port, Y(17) => 
                           CWB_MUX2_out_17_port, Y(16) => CWB_MUX2_out_16_port,
                           Y(15) => CWB_MUX2_out_15_port, Y(14) => 
                           CWB_MUX2_out_14_port, Y(13) => CWB_MUX2_out_13_port,
                           Y(12) => CWB_MUX2_out_12_port, Y(11) => 
                           CWB_MUX2_out_11_port, Y(10) => CWB_MUX2_out_10_port,
                           Y(9) => CWB_MUX2_out_9_port, Y(8) => 
                           CWB_MUX2_out_8_port, Y(7) => CWB_MUX2_out_7_port, 
                           Y(6) => CWB_MUX2_out_6_port, Y(5) => 
                           CWB_MUX2_out_5_port, Y(4) => CWB_MUX2_out_4_port, 
                           Y(3) => CWB_MUX2_out_3_port, Y(2) => 
                           CWB_MUX2_out_2_port, Y(1) => CWB_MUX2_out_1_port, 
                           Y(0) => CWB_MUX2_out_0_port);
   B2_MUX : MUX2to1_NBIT32_2 port map( A(31) => B2_out_31_port, A(30) => 
                           B2_out_30_port, A(29) => B2_out_29_port, A(28) => 
                           B2_out_28_port, A(27) => B2_out_27_port, A(26) => 
                           B2_out_26_port, A(25) => B2_out_25_port, A(24) => 
                           B2_out_24_port, A(23) => B2_out_23_port, A(22) => 
                           B2_out_22_port, A(21) => B2_out_21_port, A(20) => 
                           B2_out_20_port, A(19) => B2_out_19_port, A(18) => 
                           B2_out_18_port, A(17) => B2_out_17_port, A(16) => 
                           B2_out_16_port, A(15) => B2_out_15_port, A(14) => 
                           B2_out_14_port, A(13) => B2_out_13_port, A(12) => 
                           B2_out_12_port, A(11) => B2_out_11_port, A(10) => 
                           B2_out_10_port, A(9) => B2_out_9_port, A(8) => 
                           B2_out_8_port, A(7) => B2_out_7_port, A(6) => 
                           B2_out_6_port, A(5) => B2_out_5_port, A(4) => 
                           B2_out_4_port, A(3) => B2_out_3_port, A(2) => 
                           B2_out_2_port, A(1) => B2_out_1_port, A(0) => 
                           B2_out_0_port, B(31) => WB_in_31_port, B(30) => 
                           WB_in_30_port, B(29) => WB_in_29_port, B(28) => 
                           WB_in_28_port, B(27) => WB_in_27_port, B(26) => 
                           WB_in_26_port, B(25) => WB_in_25_port, B(24) => 
                           WB_in_24_port, B(23) => WB_in_23_port, B(22) => 
                           WB_in_22_port, B(21) => WB_in_21_port, B(20) => 
                           WB_in_20_port, B(19) => WB_in_19_port, B(18) => 
                           WB_in_18_port, B(17) => WB_in_17_port, B(16) => 
                           WB_in_16_port, B(15) => WB_in_15_port, B(14) => 
                           WB_in_14_port, B(13) => WB_in_13_port, B(12) => 
                           WB_in_12_port, B(11) => WB_in_11_port, B(10) => 
                           WB_in_10_port, B(9) => WB_in_9_port, B(8) => 
                           WB_in_8_port, B(7) => WB_in_7_port, B(6) => 
                           WB_in_6_port, B(5) => WB_in_5_port, B(4) => 
                           WB_in_4_port, B(3) => WB_in_3_port, B(2) => 
                           WB_in_2_port, B(1) => WB_in_1_port, B(0) => 
                           WB_in_0_port, SEL => FWDB2_SEL, Y(31) => 
                           B2_MUX_out_31_port, Y(30) => B2_MUX_out_30_port, 
                           Y(29) => B2_MUX_out_29_port, Y(28) => 
                           B2_MUX_out_28_port, Y(27) => B2_MUX_out_27_port, 
                           Y(26) => B2_MUX_out_26_port, Y(25) => 
                           B2_MUX_out_25_port, Y(24) => B2_MUX_out_24_port, 
                           Y(23) => B2_MUX_out_23_port, Y(22) => 
                           B2_MUX_out_22_port, Y(21) => B2_MUX_out_21_port, 
                           Y(20) => B2_MUX_out_20_port, Y(19) => 
                           B2_MUX_out_19_port, Y(18) => B2_MUX_out_18_port, 
                           Y(17) => B2_MUX_out_17_port, Y(16) => 
                           B2_MUX_out_16_port, Y(15) => B2_MUX_out_15_port, 
                           Y(14) => B2_MUX_out_14_port, Y(13) => 
                           B2_MUX_out_13_port, Y(12) => B2_MUX_out_12_port, 
                           Y(11) => B2_MUX_out_11_port, Y(10) => 
                           B2_MUX_out_10_port, Y(9) => B2_MUX_out_9_port, Y(8) 
                           => B2_MUX_out_8_port, Y(7) => B2_MUX_out_7_port, 
                           Y(6) => B2_MUX_out_6_port, Y(5) => B2_MUX_out_5_port
                           , Y(4) => B2_MUX_out_4_port, Y(3) => 
                           B2_MUX_out_3_port, Y(2) => B2_MUX_out_2_port, Y(1) 
                           => B2_MUX_out_1_port, Y(0) => B2_MUX_out_0_port);
   WBMUX : MUX2to1_NBIT32_1 port map( A(31) => ALR2_out_31_port, A(30) => 
                           ALR2_out_30_port, A(29) => ALR2_out_29_port, A(28) 
                           => ALR2_out_28_port, A(27) => ALR2_out_27_port, 
                           A(26) => ALR2_out_26_port, A(25) => ALR2_out_25_port
                           , A(24) => ALR2_out_24_port, A(23) => 
                           ALR2_out_23_port, A(22) => ALR2_out_22_port, A(21) 
                           => ALR2_out_21_port, A(20) => ALR2_out_20_port, 
                           A(19) => ALR2_out_19_port, A(18) => ALR2_out_18_port
                           , A(17) => ALR2_out_17_port, A(16) => 
                           ALR2_out_16_port, A(15) => ALR2_out_15_port, A(14) 
                           => ALR2_out_14_port, A(13) => ALR2_out_13_port, 
                           A(12) => ALR2_out_12_port, A(11) => ALR2_out_11_port
                           , A(10) => ALR2_out_10_port, A(9) => ALR2_out_9_port
                           , A(8) => ALR2_out_8_port, A(7) => ALR2_out_7_port, 
                           A(6) => ALR2_out_6_port, A(5) => ALR2_out_5_port, 
                           A(4) => ALR2_out_4_port, A(3) => ALR2_out_3_port, 
                           A(2) => ALR2_out_2_port, A(1) => ALR2_out_1_port, 
                           A(0) => ALR2_out_0_port, B(31) => LMD_out_31_port, 
                           B(30) => LMD_out_30_port, B(29) => LMD_out_29_port, 
                           B(28) => LMD_out_28_port, B(27) => LMD_out_27_port, 
                           B(26) => LMD_out_26_port, B(25) => LMD_out_25_port, 
                           B(24) => LMD_out_24_port, B(23) => LMD_out_23_port, 
                           B(22) => LMD_out_22_port, B(21) => LMD_out_21_port, 
                           B(20) => LMD_out_20_port, B(19) => LMD_out_19_port, 
                           B(18) => LMD_out_18_port, B(17) => LMD_out_17_port, 
                           B(16) => LMD_out_16_port, B(15) => LMD_out_15_port, 
                           B(14) => LMD_out_14_port, B(13) => LMD_out_13_port, 
                           B(12) => LMD_out_12_port, B(11) => LMD_out_11_port, 
                           B(10) => LMD_out_10_port, B(9) => LMD_out_9_port, 
                           B(8) => LMD_out_8_port, B(7) => LMD_out_7_port, B(6)
                           => LMD_out_6_port, B(5) => LMD_out_5_port, B(4) => 
                           LMD_out_4_port, B(3) => LMD_out_3_port, B(2) => 
                           LMD_out_2_port, B(1) => LMD_out_1_port, B(0) => 
                           LMD_out_0_port, SEL => WB_SEL, Y(31) => 
                           WB_in_31_port, Y(30) => WB_in_30_port, Y(29) => 
                           WB_in_29_port, Y(28) => WB_in_28_port, Y(27) => 
                           WB_in_27_port, Y(26) => WB_in_26_port, Y(25) => 
                           WB_in_25_port, Y(24) => WB_in_24_port, Y(23) => 
                           WB_in_23_port, Y(22) => WB_in_22_port, Y(21) => 
                           WB_in_21_port, Y(20) => WB_in_20_port, Y(19) => 
                           WB_in_19_port, Y(18) => WB_in_18_port, Y(17) => 
                           WB_in_17_port, Y(16) => WB_in_16_port, Y(15) => 
                           WB_in_15_port, Y(14) => WB_in_14_port, Y(13) => 
                           WB_in_13_port, Y(12) => WB_in_12_port, Y(11) => 
                           WB_in_11_port, Y(10) => WB_in_10_port, Y(9) => 
                           WB_in_9_port, Y(8) => WB_in_8_port, Y(7) => 
                           WB_in_7_port, Y(6) => WB_in_6_port, Y(5) => 
                           WB_in_5_port, Y(4) => WB_in_4_port, Y(3) => 
                           WB_in_3_port, Y(2) => WB_in_2_port, Y(1) => 
                           WB_in_1_port, Y(0) => WB_in_0_port);
   RF_MUX_ADDR : MUX3to1_NBIT5 port map( A(4) => RWB3_out_15_port, A(3) => 
                           RWB3_out_14_port, A(2) => RWB3_out_13_port, A(1) => 
                           RWB3_out_12_port, A(0) => RWB3_out_11_port, B(4) => 
                           RWB3_out_20_port, B(3) => RWB3_out_19_port, B(2) => 
                           RWB3_out_18_port, B(1) => RWB3_out_17_port, B(0) => 
                           RWB3_out_16_port, C(4) => X_Logic1_port, C(3) => 
                           X_Logic1_port, C(2) => X_Logic1_port, C(1) => 
                           X_Logic1_port, C(0) => X_Logic1_port, SEL(1) => 
                           RF_MUX_SEL(1), SEL(0) => RF_MUX_SEL(0), Y(4) => 
                           RF_MUX_out_4_port, Y(3) => RF_MUX_out_3_port, Y(2) 
                           => RF_MUX_out_2_port, Y(1) => RF_MUX_out_1_port, 
                           Y(0) => RF_MUX_out_0_port);
   ALU1 : ALU_NBIT32 port map( CLOCK => CLK, AluOpcode(0) => ALU_OPCODE(0), 
                           AluOpcode(1) => ALU_OPCODE(1), AluOpcode(2) => 
                           ALU_OPCODE(2), AluOpcode(3) => ALU_OPCODE(3), 
                           AluOpcode(4) => ALU_OPCODE(4), A(31) => A_in_31_port
                           , A(30) => A_in_30_port, A(29) => A_in_29_port, 
                           A(28) => A_in_28_port, A(27) => A_in_27_port, A(26) 
                           => A_in_26_port, A(25) => A_in_25_port, A(24) => 
                           A_in_24_port, A(23) => A_in_23_port, A(22) => 
                           A_in_22_port, A(21) => A_in_21_port, A(20) => 
                           A_in_20_port, A(19) => A_in_19_port, A(18) => 
                           A_in_18_port, A(17) => A_in_17_port, A(16) => 
                           A_in_16_port, A(15) => A_in_15_port, A(14) => 
                           A_in_14_port, A(13) => A_in_13_port, A(12) => 
                           A_in_12_port, A(11) => A_in_11_port, A(10) => 
                           A_in_10_port, A(9) => A_in_9_port, A(8) => 
                           A_in_8_port, A(7) => A_in_7_port, A(6) => 
                           A_in_6_port, A(5) => A_in_5_port, A(4) => 
                           A_in_4_port, A(3) => A_in_3_port, A(2) => 
                           A_in_2_port, A(1) => A_in_1_port, A(0) => 
                           A_in_0_port, B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Cin => PSW_out_6_port, ALU_out(31) => 
                           ALR_in_31_port, ALU_out(30) => ALR_in_30_port, 
                           ALU_out(29) => ALR_in_29_port, ALU_out(28) => 
                           ALR_in_28_port, ALU_out(27) => ALR_in_27_port, 
                           ALU_out(26) => ALR_in_26_port, ALU_out(25) => 
                           ALR_in_25_port, ALU_out(24) => ALR_in_24_port, 
                           ALU_out(23) => ALR_in_23_port, ALU_out(22) => 
                           ALR_in_22_port, ALU_out(21) => ALR_in_21_port, 
                           ALU_out(20) => ALR_in_20_port, ALU_out(19) => 
                           ALR_in_19_port, ALU_out(18) => ALR_in_18_port, 
                           ALU_out(17) => ALR_in_17_port, ALU_out(16) => 
                           ALR_in_16_port, ALU_out(15) => ALR_in_15_port, 
                           ALU_out(14) => ALR_in_14_port, ALU_out(13) => 
                           ALR_in_13_port, ALU_out(12) => ALR_in_12_port, 
                           ALU_out(11) => ALR_in_11_port, ALU_out(10) => 
                           ALR_in_10_port, ALU_out(9) => ALR_in_9_port, 
                           ALU_out(8) => ALR_in_8_port, ALU_out(7) => 
                           ALR_in_7_port, ALU_out(6) => ALR_in_6_port, 
                           ALU_out(5) => ALR_in_5_port, ALU_out(4) => 
                           ALR_in_4_port, ALU_out(3) => ALR_in_3_port, 
                           ALU_out(2) => ALR_in_2_port, ALU_out(1) => 
                           ALR_in_1_port, ALU_out(0) => ALR_in_0_port, Cout => 
                           PSW_in_6_port, COND(5) => PSW_in_5_port, COND(4) => 
                           PSW_in_4_port, COND(3) => PSW_in_3_port, COND(2) => 
                           PSW_in_2_port, COND(1) => PSW_in_1_port, COND(0) => 
                           PSW_in_0_port);
   FWD1 : FWDU_IR_SIZE32 port map( CLOCK => CLK, RESET => n5, EN => n41, IR(31)
                           => IR_out_31_port, IR(30) => IR_out_30_port, IR(29) 
                           => IR_out_29_port, IR(28) => IR_out_28_port, IR(27) 
                           => IR_out_27_port, IR(26) => IR_out_26_port, IR(25) 
                           => IR_out_25_port, IR(24) => IR_out_24_port, IR(23) 
                           => IR_out_23_port, IR(22) => IR_out_22_port, IR(21) 
                           => IR_out_21_port, IR(20) => IR_out_20_port, IR(19) 
                           => IR_out_19_port, IR(18) => IR_out_18_port, IR(17) 
                           => IR_out_17_port, IR(16) => IR_out_16_port, IR(15) 
                           => IR_out_15_port, IR(14) => IR_out_14_port, IR(13) 
                           => IR_out_13_port, IR(12) => IR_out_12_port, IR(11) 
                           => IR_out_11_port, IR(10) => IR_out_10_port, IR(9) 
                           => IR_out_9_port, IR(8) => IR_out_8_port, IR(7) => 
                           IR_out_7_port, IR(6) => IR_out_6_port, IR(5) => 
                           IR_out_5_port, IR(4) => IR_out_4_port, IR(3) => 
                           IR_out_3_port, IR(2) => IR_out_2_port, IR(1) => 
                           IR_out_1_port, IR(0) => IR_out_0_port, FWD_A(1) => 
                           FWDA_SEL_1_port, FWD_A(0) => FWDA_SEL_0_port, 
                           FWD_B(1) => FWDB_SEL_1_port, FWD_B(0) => 
                           FWDB_SEL_0_port, FWD_B2 => FWDB2_SEL, ZDU_SEL(1) => 
                           ZDU_SEL_1_port, ZDU_SEL(0) => ZDU_SEL_0_port);
   HDU1 : HDU_IR_SIZE32 port map( clk => CLK, rst => n7, IR(31) => 
                           IR_out_31_port, IR(30) => IR_out_30_port, IR(29) => 
                           IR_out_29_port, IR(28) => IR_out_28_port, IR(27) => 
                           IR_out_27_port, IR(26) => IR_out_26_port, IR(25) => 
                           IR_out_25_port, IR(24) => IR_out_24_port, IR(23) => 
                           IR_out_23_port, IR(22) => IR_out_22_port, IR(21) => 
                           IR_out_21_port, IR(20) => IR_out_20_port, IR(19) => 
                           IR_out_19_port, IR(18) => IR_out_18_port, IR(17) => 
                           IR_out_17_port, IR(16) => IR_out_16_port, IR(15) => 
                           IR_out_15_port, IR(14) => IR_out_14_port, IR(13) => 
                           IR_out_13_port, IR(12) => IR_out_12_port, IR(11) => 
                           IR_out_11_port, IR(10) => IR_out_10_port, IR(9) => 
                           IR_out_9_port, IR(8) => IR_out_8_port, IR(7) => 
                           IR_out_7_port, IR(6) => IR_out_6_port, IR(5) => 
                           IR_out_5_port, IR(4) => IR_out_4_port, IR(3) => 
                           IR_out_3_port, IR(2) => IR_out_2_port, IR(1) => 
                           IR_out_1_port, IR(0) => IR_out_0_port, STALL_CODE(1)
                           => STALL(1), STALL_CODE(0) => STALL(0), IF_STALL => 
                           IF_STALL, ID_STALL => n_1663, EX_STALL => EX_STALL, 
                           MEM_STALL => MEM_STALL, WB_STALL => n_1664);
   BHT1 : BHT_NBIT32_N_ENTRIES8_WORD_OFFSET0 port map( clock => CLK, rst => n10
                           , address(31) => BHT_in_31_port, address(30) => 
                           BHT_in_30_port, address(29) => BHT_in_29_port, 
                           address(28) => BHT_in_28_port, address(27) => 
                           BHT_in_27_port, address(26) => BHT_in_26_port, 
                           address(25) => BHT_in_25_port, address(24) => 
                           BHT_in_24_port, address(23) => BHT_in_23_port, 
                           address(22) => BHT_in_22_port, address(21) => 
                           BHT_in_21_port, address(20) => BHT_in_20_port, 
                           address(19) => BHT_in_19_port, address(18) => 
                           BHT_in_18_port, address(17) => BHT_in_17_port, 
                           address(16) => BHT_in_16_port, address(15) => 
                           BHT_in_15_port, address(14) => BHT_in_14_port, 
                           address(13) => BHT_in_13_port, address(12) => 
                           BHT_in_12_port, address(11) => BHT_in_11_port, 
                           address(10) => BHT_in_10_port, address(9) => 
                           BHT_in_9_port, address(8) => BHT_in_8_port, 
                           address(7) => BHT_in_7_port, address(6) => 
                           BHT_in_6_port, address(5) => BHT_in_5_port, 
                           address(4) => BHT_in_4_port, address(3) => 
                           BHT_in_3_port, address(2) => BHT_in_2_port, 
                           address(1) => BHT_in_1_port, address(0) => 
                           BHT_in_0_port, d_in => ZDU_out, w_en => n3, d_out =>
                           BHT_out);
   CWBU1 : CWBU port map( CLOCK => CLK, ALU_OP(0) => ALU_OPCODE(0), ALU_OP(1) 
                           => ALU_OPCODE(1), ALU_OP(2) => ALU_OPCODE(2), 
                           ALU_OP(3) => ALU_OPCODE(3), ALU_OP(4) => 
                           ALU_OPCODE(4), PSW(6) => PSW_out_6_port, PSW(5) => 
                           PSW_out_5_port, PSW(4) => PSW_out_4_port, PSW(3) => 
                           PSW_out_3_port, PSW(2) => PSW_out_2_port, PSW(1) => 
                           PSW_out_1_port, PSW(0) => PSW_out_0_port, 
                           COND_SEL(1) => CWB_out_1_port, COND_SEL(0) => 
                           CWB_out_0_port, CWB_SEL(1) => CWB_SEL(1), CWB_SEL(0)
                           => CWB_SEL(0), CWB_MUW_SEL(1) => CWB_MUX_SEL_1_port,
                           CWB_MUW_SEL(0) => CWB_MUX_SEL_0_port);
   RF1 : RF_NBIT32_NREG32 port map( CLK => CLK, RESET => n5, ENABLE => 
                           X_Logic1_port, RD1 => RF_RD_en, RD2 => RF_RD_en, WR 
                           => RF_WR, ADD_WR(4) => RF_MUX_out_4_port, ADD_WR(3) 
                           => RF_MUX_out_3_port, ADD_WR(2) => RF_MUX_out_2_port
                           , ADD_WR(1) => RF_MUX_out_1_port, ADD_WR(0) => 
                           RF_MUX_out_0_port, ADD_RD1(4) => IR_out_25_port, 
                           ADD_RD1(3) => IR_out_24_port, ADD_RD1(2) => 
                           IR_out_23_port, ADD_RD1(1) => IR_out_22_port, 
                           ADD_RD1(0) => IR_out_21_port, ADD_RD2(4) => 
                           IR_out_20_port, ADD_RD2(3) => IR_out_19_port, 
                           ADD_RD2(2) => IR_out_18_port, ADD_RD2(1) => 
                           IR_out_17_port, ADD_RD2(0) => IR_out_16_port, 
                           DATAIN(31) => WB_in_31_port, DATAIN(30) => 
                           WB_in_30_port, DATAIN(29) => WB_in_29_port, 
                           DATAIN(28) => WB_in_28_port, DATAIN(27) => 
                           WB_in_27_port, DATAIN(26) => WB_in_26_port, 
                           DATAIN(25) => WB_in_25_port, DATAIN(24) => 
                           WB_in_24_port, DATAIN(23) => WB_in_23_port, 
                           DATAIN(22) => WB_in_22_port, DATAIN(21) => 
                           WB_in_21_port, DATAIN(20) => WB_in_20_port, 
                           DATAIN(19) => WB_in_19_port, DATAIN(18) => 
                           WB_in_18_port, DATAIN(17) => WB_in_17_port, 
                           DATAIN(16) => WB_in_16_port, DATAIN(15) => 
                           WB_in_15_port, DATAIN(14) => WB_in_14_port, 
                           DATAIN(13) => WB_in_13_port, DATAIN(12) => 
                           WB_in_12_port, DATAIN(11) => WB_in_11_port, 
                           DATAIN(10) => WB_in_10_port, DATAIN(9) => 
                           WB_in_9_port, DATAIN(8) => WB_in_8_port, DATAIN(7) 
                           => WB_in_7_port, DATAIN(6) => WB_in_6_port, 
                           DATAIN(5) => WB_in_5_port, DATAIN(4) => WB_in_4_port
                           , DATAIN(3) => WB_in_3_port, DATAIN(2) => 
                           WB_in_2_port, DATAIN(1) => WB_in_1_port, DATAIN(0) 
                           => WB_in_0_port, OUT1(31) => RA_out_31_port, 
                           OUT1(30) => RA_out_30_port, OUT1(29) => 
                           RA_out_29_port, OUT1(28) => RA_out_28_port, OUT1(27)
                           => RA_out_27_port, OUT1(26) => RA_out_26_port, 
                           OUT1(25) => RA_out_25_port, OUT1(24) => 
                           RA_out_24_port, OUT1(23) => RA_out_23_port, OUT1(22)
                           => RA_out_22_port, OUT1(21) => RA_out_21_port, 
                           OUT1(20) => RA_out_20_port, OUT1(19) => 
                           RA_out_19_port, OUT1(18) => RA_out_18_port, OUT1(17)
                           => RA_out_17_port, OUT1(16) => RA_out_16_port, 
                           OUT1(15) => RA_out_15_port, OUT1(14) => 
                           RA_out_14_port, OUT1(13) => RA_out_13_port, OUT1(12)
                           => RA_out_12_port, OUT1(11) => RA_out_11_port, 
                           OUT1(10) => RA_out_10_port, OUT1(9) => RA_out_9_port
                           , OUT1(8) => RA_out_8_port, OUT1(7) => RA_out_7_port
                           , OUT1(6) => RA_out_6_port, OUT1(5) => RA_out_5_port
                           , OUT1(4) => RA_out_4_port, OUT1(3) => RA_out_3_port
                           , OUT1(2) => RA_out_2_port, OUT1(1) => RA_out_1_port
                           , OUT1(0) => RA_out_0_port, OUT2(31) => 
                           RB_out_31_port, OUT2(30) => RB_out_30_port, OUT2(29)
                           => RB_out_29_port, OUT2(28) => RB_out_28_port, 
                           OUT2(27) => RB_out_27_port, OUT2(26) => 
                           RB_out_26_port, OUT2(25) => RB_out_25_port, OUT2(24)
                           => RB_out_24_port, OUT2(23) => RB_out_23_port, 
                           OUT2(22) => RB_out_22_port, OUT2(21) => 
                           RB_out_21_port, OUT2(20) => RB_out_20_port, OUT2(19)
                           => RB_out_19_port, OUT2(18) => RB_out_18_port, 
                           OUT2(17) => RB_out_17_port, OUT2(16) => 
                           RB_out_16_port, OUT2(15) => RB_out_15_port, OUT2(14)
                           => RB_out_14_port, OUT2(13) => RB_out_13_port, 
                           OUT2(12) => RB_out_12_port, OUT2(11) => 
                           RB_out_11_port, OUT2(10) => RB_out_10_port, OUT2(9) 
                           => RB_out_9_port, OUT2(8) => RB_out_8_port, OUT2(7) 
                           => RB_out_7_port, OUT2(6) => RB_out_6_port, OUT2(5) 
                           => RB_out_5_port, OUT2(4) => RB_out_4_port, OUT2(3) 
                           => RB_out_3_port, OUT2(2) => RB_out_2_port, OUT2(1) 
                           => RB_out_1_port, OUT2(0) => RB_out_0_port);
   U3 : AND4_X1 port map( A1 => n15, A2 => n16, A3 => n13, A4 => n14_port, ZN 
                           => n36);
   U4 : AND2_X1 port map( A1 => SIGND, A2 => IR_out_15_port, ZN => N14);
   U5 : CLKBUF_X1 port map( A => PC2_out_0_port, Z => n1);
   U6 : CLKBUF_X1 port map( A => PC2_out_1_port, Z => n2);
   U7 : XNOR2_X1 port map( A => n38, B => n32, ZN => n39);
   U8 : CLKBUF_X1 port map( A => BPR_EN2, Z => n3);
   U9 : BUF_X1 port map( A => n31, Z => n8);
   U10 : BUF_X1 port map( A => n31, Z => n9);
   U11 : BUF_X1 port map( A => n30, Z => n5);
   U12 : BUF_X1 port map( A => n31, Z => n10);
   U13 : BUF_X1 port map( A => n30, Z => n7);
   U14 : BUF_X1 port map( A => n30, Z => n6);
   U15 : BUF_X1 port map( A => n41, Z => n11);
   U16 : BUF_X1 port map( A => n29, Z => n30);
   U17 : BUF_X1 port map( A => n29, Z => n31);
   U18 : BUF_X1 port map( A => n22, Z => n27);
   U19 : BUF_X1 port map( A => MEM_ENABLE, Z => n12);
   U20 : BUF_X1 port map( A => ID_ENABLE, Z => n21);
   U21 : BUF_X1 port map( A => EX_ENABLE, Z => n19);
   U22 : BUF_X1 port map( A => n27, Z => n24);
   U23 : BUF_X1 port map( A => n27, Z => n25);
   U24 : BUF_X1 port map( A => n27, Z => n26);
   U25 : INV_X1 port map( A => IF_STALL, ZN => n41);
   U26 : BUF_X1 port map( A => n28, Z => n23);
   U27 : BUF_X1 port map( A => n22, Z => n28);
   U28 : XNOR2_X1 port map( A => n4, B => RWB1_out_26_port, ZN => n38);
   U29 : AND4_X1 port map( A1 => n36, A2 => n35, A3 => n34, A4 => n33, ZN => n4
                           );
   U30 : NOR2_X1 port map( A1 => MEM_STALL, A2 => n43, ZN => MEM_ENABLE);
   U31 : INV_X1 port map( A => MEM_EN, ZN => n43);
   U32 : OR4_X1 port map( A1 => ZDU_MUX_out_13_port, A2 => ZDU_MUX_out_12_port,
                           A3 => ZDU_MUX_out_15_port, A4 => ZDU_MUX_out_14_port
                           , ZN => n17);
   U33 : NOR4_X1 port map( A1 => ZDU_MUX_out_2_port, A2 => ZDU_MUX_out_29_port,
                           A3 => ZDU_MUX_out_28_port, A4 => ZDU_MUX_out_27_port
                           , ZN => n14_port);
   U34 : NOR4_X1 port map( A1 => ZDU_MUX_out_26_port, A2 => ZDU_MUX_out_25_port
                           , A3 => ZDU_MUX_out_24_port, A4 => 
                           ZDU_MUX_out_23_port, ZN => n13);
   U35 : NOR4_X1 port map( A1 => ZDU_MUX_out_9_port, A2 => ZDU_MUX_out_8_port, 
                           A3 => ZDU_MUX_out_7_port, A4 => ZDU_MUX_out_6_port, 
                           ZN => n16);
   U36 : NOR4_X1 port map( A1 => ZDU_MUX_out_5_port, A2 => ZDU_MUX_out_4_port, 
                           A3 => ZDU_MUX_out_3_port, A4 => ZDU_MUX_out_30_port,
                           ZN => n15);
   U37 : INV_X1 port map( A => n18, ZN => n40);
   U38 : NOR2_X1 port map( A1 => EX_STALL, A2 => n42, ZN => EX_ENABLE);
   U39 : INV_X1 port map( A => EX_EN, ZN => n42);
   U40 : AND2_X1 port map( A1 => ID_EN, A2 => n11, ZN => ID_ENABLE);
   U41 : AND2_X1 port map( A1 => RF_RD, A2 => n11, ZN => RF_RD_en);
   U42 : BUF_X1 port map( A => RST, Z => n29);
   U43 : BUF_X1 port map( A => DATA_IN(7), Z => n22);
   U44 : INV_X1 port map( A => n3, ZN => n20);
   U45 : AOI21_X1 port map( B1 => BPR_EN, B2 => BHT_out, A => UCB_EN, ZN => n18
                           );
   U46 : INV_X1 port map( A => BMP, ZN => n37);
   U47 : INV_X1 port map( A => PRD_OUT, ZN => n32);
   U48 : NOR2_X1 port map( A1 => n37, A2 => n32, ZN => IRAMMUX_SEL);
   U49 : NOR4_X1 port map( A1 => ZDU_MUX_out_19_port, A2 => ZDU_MUX_out_20_port
                           , A3 => ZDU_MUX_out_21_port, A4 => 
                           ZDU_MUX_out_22_port, ZN => n35);
   U50 : NOR4_X1 port map( A1 => ZDU_MUX_out_11_port, A2 => ZDU_MUX_out_16_port
                           , A3 => ZDU_MUX_out_17_port, A4 => 
                           ZDU_MUX_out_18_port, ZN => n34);
   U51 : NOR4_X1 port map( A1 => n17, A2 => ZDU_MUX_out_0_port, A3 => 
                           ZDU_MUX_out_1_port, A4 => ZDU_MUX_out_10_port, ZN =>
                           n33);
   U52 : INV_X1 port map( A => n38, ZN => ZDU_out);
   U53 : NOR3_X1 port map( A1 => n40, A2 => PRD_OUT, A3 => n37, ZN => 
                           PC_SEL_1_port);
   U54 : NOR2_X1 port map( A1 => n39, A2 => n20, ZN => BMP);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26 is

   port( Clk, Rst : in std_logic;  STALL : in std_logic_vector (1 downto 0);  
         IR_IN : in std_logic_vector (31 downto 0);  BMP : in std_logic;  ID_EN
         , RF_RD, SIGND, IMM_SEL, BPR_EN, UCB_EN : out std_logic;  ALU_OPCODE :
         out std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, ALUB_SEL, MEM_EN, 
         MEM_DATA_SEL, MEM_RD, MEM_WR, CS, MEM_BLC0, MEM_BLC1, LD_SEL0, LD_SEL1
         , LD_SEL2, ALR2_SEL, CWB_SEL0, CWB_SEL1, WB_SEL, RF_WR, RF_MUX_SEL0, 
         RF_MUX_SEL1 : out std_logic);

end CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26;

architecture SYN_dlx_cu_hw of 
   CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal ALU_OPCODE_4_port, ALU_OPCODE_3_port, ALU_OPCODE_2_port, 
      ALU_OPCODE_1_port, ALU_OPCODE_0_port, MEM_EN_port, MEM_DATA_SEL_port, 
      MEM_RD_port, MEM_WR_port, CS_port, MEM_BLC0_port, MEM_BLC1_port, 
      LD_SEL0_port, LD_SEL1_port, LD_SEL2_port, ALR2_SEL_port, CWB_SEL0_port, 
      CWB_SEL1_port, WB_SEL_port, RF_WR_port, RF_MUX_SEL0_port, 
      RF_MUX_SEL1_port, cw3_16_port, cw3_14_port, cw3_13_port, cw3_12_port, 
      cw3_11_port, cw3_10_port, cw3_9_port, cw3_8_port, cw3_7_port, cw3_0_port,
      cw4_3_port, cw4_2_port, cw4_1_port, cw4_0_port, aluOpcode1_4_port, 
      aluOpcode1_3_port, aluOpcode1_2_port, aluOpcode1_1_port, 
      aluOpcode1_0_port, N86, n3, n4, n6, n10, n12, n14, n16, n18, n20, n22, 
      n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n45, n46, n47, n48
      , n49, n50, n51, n52, n53, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86_port, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n189, n190, n191, n192, n1, n2, n5, n7, n8, n9, n11, n13, n15, n17, n19, 
      n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n54, n55, n56
      , n57, n58, n59, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, 
      n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, 
      n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, 
      n_1690, n_1691 : std_logic;

begin
   ALU_OPCODE <= ( ALU_OPCODE_4_port, ALU_OPCODE_3_port, ALU_OPCODE_2_port, 
      ALU_OPCODE_1_port, ALU_OPCODE_0_port );
   MEM_EN <= MEM_EN_port;
   MEM_DATA_SEL <= MEM_DATA_SEL_port;
   MEM_RD <= MEM_RD_port;
   MEM_WR <= MEM_WR_port;
   CS <= CS_port;
   MEM_BLC0 <= MEM_BLC0_port;
   MEM_BLC1 <= MEM_BLC1_port;
   LD_SEL0 <= LD_SEL0_port;
   LD_SEL1 <= LD_SEL1_port;
   LD_SEL2 <= LD_SEL2_port;
   ALR2_SEL <= ALR2_SEL_port;
   CWB_SEL0 <= CWB_SEL0_port;
   CWB_SEL1 <= CWB_SEL1_port;
   WB_SEL <= WB_SEL_port;
   RF_WR <= RF_WR_port;
   RF_MUX_SEL0 <= RF_MUX_SEL0_port;
   RF_MUX_SEL1 <= RF_MUX_SEL1_port;
   
   cw4_reg_16_inst : DFFR_X1 port map( D => n10, CK => Clk, RN => n11, Q => 
                           MEM_EN_port, QN => n_1665);
   cw4_reg_15_inst : DFFR_X1 port map( D => n12, CK => Clk, RN => n11, Q => 
                           MEM_DATA_SEL_port, QN => n_1666);
   cw4_reg_14_inst : DFFR_X1 port map( D => n14, CK => Clk, RN => n11, Q => 
                           MEM_RD_port, QN => n_1667);
   cw4_reg_13_inst : DFFR_X1 port map( D => n16, CK => Clk, RN => n11, Q => 
                           MEM_WR_port, QN => n_1668);
   cw4_reg_12_inst : DFFR_X1 port map( D => n18, CK => Clk, RN => n11, Q => 
                           CS_port, QN => n_1669);
   cw4_reg_11_inst : DFFR_X1 port map( D => n20, CK => Clk, RN => n11, Q => 
                           MEM_BLC0_port, QN => n_1670);
   cw4_reg_10_inst : DFFR_X1 port map( D => n22, CK => Clk, RN => n11, Q => 
                           MEM_BLC1_port, QN => n_1671);
   cw4_reg_9_inst : DFFR_X1 port map( D => n24, CK => Clk, RN => n11, Q => 
                           LD_SEL0_port, QN => n_1672);
   cw4_reg_8_inst : DFFR_X1 port map( D => n26, CK => Clk, RN => n11, Q => 
                           LD_SEL1_port, QN => n_1673);
   cw4_reg_7_inst : DFFR_X1 port map( D => n28, CK => Clk, RN => n9, Q => 
                           LD_SEL2_port, QN => n_1674);
   cw4_reg_6_inst : DFFR_X1 port map( D => n30, CK => Clk, RN => n9, Q => 
                           ALR2_SEL_port, QN => n_1675);
   cw4_reg_5_inst : DFFR_X1 port map( D => n32, CK => Clk, RN => n9, Q => 
                           CWB_SEL0_port, QN => n_1676);
   cw4_reg_4_inst : DFFR_X1 port map( D => n34, CK => Clk, RN => n9, Q => 
                           CWB_SEL1_port, QN => n_1677);
   cw4_reg_3_inst : DFFR_X1 port map( D => n36, CK => Clk, RN => n9, Q => 
                           cw4_3_port, QN => n_1678);
   cw4_reg_2_inst : DFFR_X1 port map( D => n38, CK => Clk, RN => n9, Q => 
                           cw4_2_port, QN => n_1679);
   cw4_reg_1_inst : DFFR_X1 port map( D => n40, CK => Clk, RN => n9, Q => 
                           cw4_1_port, QN => n_1680);
   cw4_reg_0_inst : DFFR_X1 port map( D => n42, CK => Clk, RN => n9, Q => 
                           cw4_0_port, QN => n_1681);
   cw5_reg_3_inst : DFFR_X1 port map( D => n44, CK => Clk, RN => n9, Q => 
                           WB_SEL_port, QN => n_1682);
   cw5_reg_2_inst : DFFR_X1 port map( D => n45, CK => Clk, RN => n9, Q => 
                           RF_WR_port, QN => n_1683);
   cw5_reg_1_inst : DFFR_X1 port map( D => n46, CK => Clk, RN => n9, Q => 
                           RF_MUX_SEL0_port, QN => n_1684);
   cw5_reg_0_inst : DFFR_X1 port map( D => n47, CK => Clk, RN => n8, Q => 
                           RF_MUX_SEL1_port, QN => n_1685);
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => n192, CK => Clk, RN => n8, Q 
                           => aluOpcode1_4_port, QN => n48);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => n49, CK => Clk, RN => n8, Q 
                           => aluOpcode1_3_port, QN => n_1686);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => n191, CK => Clk, RN => n8, Q 
                           => aluOpcode1_2_port, QN => n50);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => n4, CK => Clk, RN => n8, Q =>
                           ALU_OPCODE_2_port, QN => n_1687);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => n190, CK => Clk, RN => n8, Q 
                           => aluOpcode1_1_port, QN => n51);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => n189, CK => Clk, RN => n8, Q 
                           => aluOpcode1_0_port, QN => n52);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => n6, CK => Clk, RN => n8, Q =>
                           ALU_OPCODE_0_port, QN => n_1688);
   UCB_EN <= '0';
   BPR_EN <= '0';
   IMM_SEL <= '0';
   SIGND <= '0';
   RF_RD <= '0';
   ID_EN <= '0';
   U199 : NAND3_X1 port map( A1 => n133, A2 => n105, A3 => n120, ZN => n114);
   U200 : NAND3_X1 port map( A1 => n112, A2 => n142, A3 => n143, ZN => n85);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => n3, CK => Clk, RN => n8, Q =>
                           ALU_OPCODE_3_port, QN => n_1689);
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => n2, CK => Clk, RN => n17, Q 
                           => ALU_OPCODE_4_port, QN => n_1690);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => n1, CK => Clk, RN => n17, Q 
                           => ALU_OPCODE_1_port, QN => n_1691);
   U3 : AOI22_X1 port map( A1 => n148, A2 => cw3_0_port, B1 => n53, B2 => 
                           cw4_0_port, ZN => n152);
   U4 : AOI22_X1 port map( A1 => n5, A2 => cw3_7_port, B1 => n53, B2 => 
                           LD_SEL2_port, ZN => n159);
   U5 : AOI22_X1 port map( A1 => n148, A2 => cw3_8_port, B1 => n53, B2 => 
                           LD_SEL1_port, ZN => n160);
   U6 : AOI22_X1 port map( A1 => n5, A2 => cw3_9_port, B1 => n53, B2 => 
                           LD_SEL0_port, ZN => n161);
   U7 : AOI22_X1 port map( A1 => n5, A2 => cw3_10_port, B1 => n53, B2 => 
                           MEM_BLC1_port, ZN => n162);
   U8 : AOI22_X1 port map( A1 => n5, A2 => cw3_11_port, B1 => n53, B2 => 
                           MEM_BLC0_port, ZN => n163);
   U9 : AOI22_X1 port map( A1 => n5, A2 => cw3_12_port, B1 => n53, B2 => 
                           CS_port, ZN => n164);
   U10 : AOI22_X1 port map( A1 => n5, A2 => cw3_13_port, B1 => n53, B2 => 
                           MEM_WR_port, ZN => n165);
   U11 : AOI22_X1 port map( A1 => n5, A2 => cw3_14_port, B1 => n53, B2 => 
                           MEM_RD_port, ZN => n166);
   U12 : NAND2_X2 port map( A1 => n53, A2 => MEM_DATA_SEL_port, ZN => n167);
   U13 : AOI22_X1 port map( A1 => n148, A2 => cw3_16_port, B1 => n53, B2 => 
                           MEM_EN_port, ZN => n168);
   U14 : NAND2_X2 port map( A1 => cw4_1_port, A2 => n53, ZN => n153);
   U15 : NAND2_X2 port map( A1 => n53, A2 => cw4_2_port, ZN => n154);
   U16 : NAND2_X2 port map( A1 => n53, A2 => cw4_3_port, ZN => n155);
   U17 : NAND2_X2 port map( A1 => n53, A2 => CWB_SEL1_port, ZN => n156);
   U18 : NAND2_X2 port map( A1 => n53, A2 => CWB_SEL0_port, ZN => n157);
   U19 : NAND2_X2 port map( A1 => n53, A2 => ALR2_SEL_port, ZN => n158);
   U20 : NOR4_X1 port map( A1 => n27, A2 => n29, A3 => IR_IN(29), A4 => 
                           IR_IN(31), ZN => n91);
   U21 : INV_X1 port map( A => n79, ZN => n1);
   U22 : INV_X1 port map( A => n75, ZN => n2);
   U23 : INV_X1 port map( A => n148, ZN => n53);
   U30 : OAI22_X1 port map( A1 => n101, A2 => n136, B1 => n57, B2 => n100, ZN 
                           => n126);
   U31 : INV_X1 port map( A => n136, ZN => n54);
   U32 : BUF_X1 port map( A => n148, Z => n5);
   U33 : BUF_X1 port map( A => n15, Z => n9);
   U34 : BUF_X1 port map( A => n15, Z => n8);
   U35 : NOR2_X1 port map( A1 => n7, A2 => BMP, ZN => n76);
   U36 : INV_X1 port map( A => BMP, ZN => n74);
   U37 : NOR2_X1 port map( A1 => n31, A2 => n112, ZN => n86_port);
   U38 : AOI22_X1 port map( A1 => n90, A2 => n107, B1 => n123, B2 => n93, ZN =>
                           n120);
   U39 : AOI22_X1 port map( A1 => n89, A2 => n31, B1 => n90, B2 => n91, ZN => 
                           n88);
   U40 : NOR2_X1 port map( A1 => n124, A2 => n110, ZN => n93);
   U41 : NOR2_X1 port map( A1 => n25, A2 => n110, ZN => n92);
   U42 : NAND2_X1 port map( A1 => n27, A2 => n29, ZN => n110);
   U43 : AOI21_X1 port map( B1 => n123, B2 => n108, A => n114, ZN => n131);
   U44 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => n101);
   U45 : INV_X1 port map( A => n134, ZN => n31);
   U46 : NOR2_X1 port map( A1 => n97, A2 => n137, ZN => n116);
   U47 : NOR4_X1 port map( A1 => n101, A2 => n43, A3 => n55, A4 => n56, ZN => 
                           n137);
   U48 : OAI21_X1 port map( B1 => n112, B2 => n123, A => n91, ZN => n122);
   U49 : NAND2_X1 port map( A1 => n140, A2 => n56, ZN => n100);
   U50 : OAI21_X1 port map( B1 => n112, B2 => n90, A => n91, ZN => n132);
   U51 : OAI21_X1 port map( B1 => n108, B2 => n92, A => n109, ZN => n104);
   U52 : INV_X1 port map( A => n103, ZN => n39);
   U53 : OR2_X1 port map( A1 => n90, A2 => n109, ZN => n123);
   U54 : NAND2_X1 port map( A1 => n141, A2 => n55, ZN => n136);
   U55 : INV_X1 port map( A => n107, ZN => n19);
   U56 : INV_X1 port map( A => n95, ZN => n57);
   U57 : INV_X1 port map( A => n89, ZN => n23);
   U58 : BUF_X1 port map( A => n17, Z => n15);
   U59 : BUF_X1 port map( A => n13, Z => n11);
   U60 : BUF_X1 port map( A => n17, Z => n13);
   U61 : INV_X1 port map( A => n80, ZN => n6);
   U62 : AOI22_X1 port map( A1 => aluOpcode1_0_port, A2 => n76, B1 => 
                           ALU_OPCODE_0_port, B2 => n7, ZN => n80);
   U63 : INV_X1 port map( A => n128, ZN => n49);
   U64 : OAI211_X1 port map( C1 => n85, C2 => n130, A => n131, B => n132, ZN =>
                           n129);
   U65 : INV_X1 port map( A => n77, ZN => n3);
   U66 : OAI21_X1 port map( B1 => N86, B2 => n52, A => n81, ZN => n189);
   U67 : OAI21_X1 port map( B1 => n82, B2 => n83, A => N86, ZN => n81);
   U68 : NAND4_X1 port map( A1 => n104, A2 => n105, A3 => n19, A4 => n106, ZN 
                           => n82);
   U69 : OAI221_X1 port map( B1 => n84, B2 => n85, C1 => n86_port, C2 => n87, A
                           => n88, ZN => n83);
   U70 : INV_X1 port map( A => n78, ZN => n4);
   U71 : OAI22_X1 port map( A1 => N86, A2 => n48, B1 => n7, B2 => n106, ZN => 
                           n192);
   U72 : OAI22_X1 port map( A1 => N86, A2 => n51, B1 => n7, B2 => n111, ZN => 
                           n190);
   U73 : AOI211_X1 port map( C1 => n107, C2 => n112, A => n113, B => n114, ZN 
                           => n111);
   U74 : OAI221_X1 port map( B1 => n35, B2 => n85, C1 => n86_port, C2 => n23, A
                           => n106, ZN => n113);
   U75 : INV_X1 port map( A => n115, ZN => n35);
   U76 : OAI22_X1 port map( A1 => N86, A2 => n50, B1 => n7, B2 => n118, ZN => 
                           n191);
   U77 : AOI211_X1 port map( C1 => n107, C2 => n31, A => n119, B => n21, ZN => 
                           n118);
   U78 : INV_X1 port map( A => n120, ZN => n21);
   U79 : OAI221_X1 port map( B1 => n121, B2 => n85, C1 => n86_port, C2 => n23, 
                           A => n122, ZN => n119);
   U80 : INV_X1 port map( A => n158, ZN => n30);
   U81 : INV_X1 port map( A => n167, ZN => n12);
   U82 : INV_X1 port map( A => n147, ZN => n47);
   U83 : AOI22_X1 port map( A1 => n5, A2 => cw4_0_port, B1 => n53, B2 => 
                           RF_MUX_SEL1_port, ZN => n147);
   U84 : INV_X1 port map( A => n149, ZN => n46);
   U85 : AOI22_X1 port map( A1 => n5, A2 => cw4_1_port, B1 => n53, B2 => 
                           RF_MUX_SEL0_port, ZN => n149);
   U86 : INV_X1 port map( A => n150, ZN => n45);
   U87 : AOI22_X1 port map( A1 => n148, A2 => cw4_2_port, B1 => n53, B2 => 
                           RF_WR_port, ZN => n150);
   U88 : INV_X1 port map( A => n152, ZN => n42);
   U89 : INV_X1 port map( A => n153, ZN => n40);
   U90 : INV_X1 port map( A => n154, ZN => n38);
   U91 : INV_X1 port map( A => n155, ZN => n36);
   U92 : INV_X1 port map( A => n156, ZN => n34);
   U93 : INV_X1 port map( A => n157, ZN => n32);
   U94 : INV_X1 port map( A => n159, ZN => n28);
   U95 : INV_X1 port map( A => n160, ZN => n26);
   U96 : INV_X1 port map( A => n161, ZN => n24);
   U97 : INV_X1 port map( A => n162, ZN => n22);
   U98 : INV_X1 port map( A => n163, ZN => n20);
   U99 : INV_X1 port map( A => n164, ZN => n18);
   U100 : INV_X1 port map( A => n165, ZN => n16);
   U101 : INV_X1 port map( A => n166, ZN => n14);
   U102 : INV_X1 port map( A => n168, ZN => n10);
   U103 : INV_X1 port map( A => n151, ZN => n44);
   U104 : NOR3_X1 port map( A1 => n124, A2 => IR_IN(30), A3 => n29, ZN => n107)
                           ;
   U105 : NOR4_X1 port map( A1 => n43, A2 => n55, A3 => IR_IN(2), A4 => 
                           IR_IN(4), ZN => n103);
   U106 : NOR2_X1 port map( A1 => IR_IN(27), A2 => IR_IN(26), ZN => n112);
   U107 : NOR2_X1 port map( A1 => n58, A2 => IR_IN(0), ZN => n95);
   U108 : NOR3_X1 port map( A1 => n110, A2 => IR_IN(31), A3 => IR_IN(29), ZN =>
                           n143);
   U109 : NOR3_X1 port map( A1 => n124, A2 => IR_IN(28), A3 => n27, ZN => n89);
   U110 : NOR3_X1 port map( A1 => n55, A2 => IR_IN(2), A3 => n43, ZN => n102);
   U111 : NOR3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(4), A3 => n43, ZN => 
                           n140);
   U112 : AOI211_X1 port map( C1 => n54, C2 => n95, A => n96, B => n97, ZN => 
                           n84);
   U113 : OAI222_X1 port map( A1 => IR_IN(1), A2 => n98, B1 => n99, B2 => n59, 
                           C1 => n100, C2 => n101, ZN => n96);
   U114 : AOI21_X1 port map( B1 => n102, B2 => IR_IN(1), A => n103, ZN => n99);
   U115 : AOI211_X1 port map( C1 => n54, C2 => IR_IN(1), A => n125, B => n126, 
                           ZN => n121);
   U116 : OAI22_X1 port map( A1 => IR_IN(1), A2 => n39, B1 => n127, B2 => n98, 
                           ZN => n125);
   U117 : AOI21_X1 port map( B1 => IR_IN(0), B2 => n58, A => n95, ZN => n127);
   U118 : NOR2_X1 port map( A1 => n33, A2 => IR_IN(26), ZN => n90);
   U119 : NOR3_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), A3 => n146, ZN => 
                           n142);
   U120 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN 
                           => n146);
   U121 : NOR3_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), A3 => n56, ZN => 
                           n141);
   U122 : NAND4_X1 port map( A1 => IR_IN(3), A2 => n142, A3 => n144, A4 => n145
                           , ZN => n106);
   U123 : AND2_X1 port map( A1 => n95, A2 => n141, ZN => n144);
   U124 : NOR4_X1 port map( A1 => IR_IN(31), A2 => IR_IN(29), A3 => n110, A4 =>
                           n134, ZN => n145);
   U125 : NOR3_X1 port map( A1 => n92, A2 => n93, A3 => n94, ZN => n87);
   U126 : NOR3_X1 port map( A1 => n25, A2 => IR_IN(30), A3 => IR_IN(29), ZN => 
                           n94);
   U127 : OAI21_X1 port map( B1 => n57, B2 => n98, A => n138, ZN => n97);
   U128 : NAND4_X1 port map( A1 => IR_IN(2), A2 => n58, A3 => IR_IN(3), A4 => 
                           n139, ZN => n138);
   U129 : NOR2_X1 port map( A1 => n59, A2 => n43, ZN => n139);
   U130 : INV_X1 port map( A => IR_IN(5), ZN => n43);
   U131 : NAND4_X1 port map( A1 => n112, A2 => IR_IN(30), A3 => IR_IN(28), A4 
                           => IR_IN(29), ZN => n133);
   U132 : INV_X1 port map( A => IR_IN(1), ZN => n58);
   U133 : NAND2_X1 port map( A1 => n140, A2 => IR_IN(2), ZN => n98);
   U134 : OAI211_X1 port map( C1 => n101, C2 => n98, A => n37, B => n116, ZN =>
                           n115);
   U135 : INV_X1 port map( A => n117, ZN => n37);
   U136 : OAI22_X1 port map( A1 => n58, A2 => n100, B1 => IR_IN(1), B2 => n39, 
                           ZN => n117);
   U137 : INV_X1 port map( A => IR_IN(3), ZN => n55);
   U138 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(28), A3 => IR_IN(29),
                           A4 => n31, ZN => n105);
   U139 : INV_X1 port map( A => IR_IN(28), ZN => n29);
   U140 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n25, ZN => n124);
   U141 : INV_X1 port map( A => IR_IN(2), ZN => n56);
   U142 : INV_X1 port map( A => IR_IN(31), ZN => n25);
   U143 : INV_X1 port map( A => IR_IN(30), ZN => n27);
   U144 : INV_X1 port map( A => IR_IN(0), ZN => n59);
   U145 : AND3_X1 port map( A1 => IR_IN(29), A2 => n29, A3 => IR_IN(30), ZN => 
                           n108);
   U146 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n33, ZN => n134);
   U147 : INV_X1 port map( A => IR_IN(27), ZN => n33);
   U148 : AND2_X1 port map( A1 => IR_IN(27), A2 => IR_IN(26), ZN => n109);
   U149 : AND3_X1 port map( A1 => n41, A2 => n116, A3 => n135, ZN => n130);
   U150 : INV_X1 port map( A => n126, ZN => n41);
   U151 : AOI22_X1 port map( A1 => n102, A2 => IR_IN(1), B1 => n54, B2 => n95, 
                           ZN => n135);
   U152 : INV_X1 port map( A => Rst, ZN => n17);
   ALUB_SEL <= '0';
   ALUA_SEL <= '0';
   cw3_16_port <= '0';
   cw3_14_port <= '0';
   cw3_13_port <= '0';
   cw3_12_port <= '0';
   cw3_11_port <= '0';
   cw3_10_port <= '0';
   cw3_9_port <= '0';
   cw3_8_port <= '0';
   cw3_7_port <= '0';
   cw3_0_port <= '0';
   EX_EN <= '0';
   U166 : AOI22_X1 port map( A1 => aluOpcode1_1_port, A2 => n76, B1 => 
                           ALU_OPCODE_1_port, B2 => n7, ZN => n79);
   U167 : AOI22_X1 port map( A1 => n5, A2 => cw4_3_port, B1 => n53, B2 => 
                           WB_SEL_port, ZN => n151);
   U168 : AOI22_X1 port map( A1 => aluOpcode1_3_port, A2 => n76, B1 => 
                           ALU_OPCODE_3_port, B2 => n7, ZN => n77);
   U169 : AOI22_X1 port map( A1 => aluOpcode1_2_port, A2 => n76, B1 => 
                           ALU_OPCODE_2_port, B2 => n7, ZN => n78);
   U170 : OAI21_X1 port map( B1 => STALL(1), B2 => STALL(0), A => n74, ZN => 
                           N86);
   U171 : INV_X1 port map( A => N86, ZN => n7);
   U172 : NAND2_X1 port map( A1 => STALL(1), A2 => n74, ZN => n148);
   U173 : AOI22_X1 port map( A1 => n7, A2 => aluOpcode1_3_port, B1 => N86, B2 
                           => n129, ZN => n128);
   U174 : AOI22_X1 port map( A1 => aluOpcode1_4_port, A2 => n76, B1 => 
                           ALU_OPCODE_4_port, B2 => n7, ZN => n75);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector (31 
         downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out std_logic_vector (31 
         downto 0);  BLC : out std_logic_vector (1 downto 0);  MEM_WR, MEM_RD :
         out std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component Datapath
      port( CLK, RST : in std_logic;  DATA_IN, IRAM_OUT : in std_logic_vector 
            (31 downto 0);  IRAM_ADDR, DATA_OUT, DATA_ADDR : out 
            std_logic_vector (31 downto 0);  BMP : inout std_logic;  STALL : 
            out std_logic_vector (1 downto 0);  ID_EN, RF_RD, SIGND, IMM_SEL, 
            BPR_EN : in std_logic;  ALU_OPCODE : in std_logic_vector (0 to 4); 
            EX_EN, ALUA_SEL, ALUB_SEL, UCB_EN, MEM_EN, MEM_DATA_SEL : in 
            std_logic;  LD_SEL : in std_logic_vector (2 downto 0);  ALR2_SEL : 
            in std_logic;  CWB_SEL : in std_logic_vector (1 downto 0);  WB_SEL,
            RF_WR : in std_logic;  RF_MUX_SEL : in std_logic_vector (1 downto 
            0));
   end component;
   
   component 
      CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26
      port( Clk, Rst : in std_logic;  STALL : in std_logic_vector (1 downto 0);
            IR_IN : in std_logic_vector (31 downto 0);  BMP : in std_logic;  
            ID_EN, RF_RD, SIGND, IMM_SEL, BPR_EN, UCB_EN : out std_logic;  
            ALU_OPCODE : out std_logic_vector (0 to 4);  EX_EN, ALUA_SEL, 
            ALUB_SEL, MEM_EN, MEM_DATA_SEL, MEM_RD, MEM_WR, CS, MEM_BLC0, 
            MEM_BLC1, LD_SEL0, LD_SEL1, LD_SEL2, ALR2_SEL, CWB_SEL0, CWB_SEL1, 
            WB_SEL, RF_WR, RF_MUX_SEL0, RF_MUX_SEL1 : out std_logic);
   end component;
   
   signal STALL_CODE_1_port, STALL_CODE_0_port, BMP_i, ID_EN_i, RF_RD_i, 
      SIGND_i, IMM_SEL_i, BPR_EN_i, UCB_EN_i, ALU_OPCODE_i_0_port, 
      ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_4_port, MEM_EN_i, MEM_DATA_SEL_i, LD_SEL_i_2_port, 
      LD_SEL_i_1_port, LD_SEL_i_0_port, ALR2_SEL_i, CWB_SEL_i_1_port, 
      CWB_SEL_i_0_port, WB_SEL_i, RF_WR_i, RF_MUX_SEL_i_1_port, 
      RF_MUX_SEL_i_0_port, n1, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701 : std_logic;
   
   signal ALU_OPCODE_pin : std_logic_vector (0 to 4);

begin
   
   ( ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port ) <= ALU_OPCODE_pin;
   CU_I : CU_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE26
      port map( Clk => Clk, Rst => Rst, STALL(1) => STALL_CODE_1_port, STALL(0)
      => STALL_CODE_0_port, IR_IN(31) => IRAM_OUT(31), IR_IN(30) => 
      IRAM_OUT(30), IR_IN(29) => IRAM_OUT(29), IR_IN(28) => IRAM_OUT(28), 
      IR_IN(27) => IRAM_OUT(27), IR_IN(26) => IRAM_OUT(26), IR_IN(25) => 
      IRAM_OUT(25), IR_IN(24) => IRAM_OUT(24), IR_IN(23) => IRAM_OUT(23), 
      IR_IN(22) => IRAM_OUT(22), IR_IN(21) => IRAM_OUT(21), IR_IN(20) => 
      IRAM_OUT(20), IR_IN(19) => IRAM_OUT(19), IR_IN(18) => IRAM_OUT(18), 
      IR_IN(17) => IRAM_OUT(17), IR_IN(16) => IRAM_OUT(16), IR_IN(15) => 
      IRAM_OUT(15), IR_IN(14) => IRAM_OUT(14), IR_IN(13) => IRAM_OUT(13), 
      IR_IN(12) => IRAM_OUT(12), IR_IN(11) => IRAM_OUT(11), IR_IN(10) => 
      IRAM_OUT(10), IR_IN(9) => IRAM_OUT(9), IR_IN(8) => IRAM_OUT(8), IR_IN(7) 
      => IRAM_OUT(7), IR_IN(6) => IRAM_OUT(6), IR_IN(5) => IRAM_OUT(5), 
      IR_IN(4) => IRAM_OUT(4), IR_IN(3) => IRAM_OUT(3), IR_IN(2) => IRAM_OUT(2)
      , IR_IN(1) => IRAM_OUT(1), IR_IN(0) => IRAM_OUT(0), BMP => BMP_i, ID_EN 
      => n_1692, RF_RD => n_1693, SIGND => n_1694, IMM_SEL => n_1695, BPR_EN =>
      n_1696, UCB_EN => n_1697, ALU_OPCODE => ALU_OPCODE_pin, EX_EN => n_1698, 
      ALUA_SEL => n_1699, ALUB_SEL => n_1700, MEM_EN => MEM_EN_i, MEM_DATA_SEL 
      => MEM_DATA_SEL_i, MEM_RD => MEM_RD, MEM_WR => MEM_WR, CS => n_1701, 
      MEM_BLC0 => BLC(0), MEM_BLC1 => BLC(1), LD_SEL0 => LD_SEL_i_0_port, 
      LD_SEL1 => LD_SEL_i_1_port, LD_SEL2 => LD_SEL_i_2_port, ALR2_SEL => 
      ALR2_SEL_i, CWB_SEL0 => CWB_SEL_i_0_port, CWB_SEL1 => CWB_SEL_i_1_port, 
      WB_SEL => WB_SEL_i, RF_WR => RF_WR_i, RF_MUX_SEL0 => RF_MUX_SEL_i_0_port,
      RF_MUX_SEL1 => RF_MUX_SEL_i_1_port);
   DATAP : Datapath port map( CLK => Clk, RST => Rst, DATA_IN(31) => 
                           DATA_IN(31), DATA_IN(30) => DATA_IN(30), DATA_IN(29)
                           => DATA_IN(29), DATA_IN(28) => DATA_IN(28), 
                           DATA_IN(27) => DATA_IN(27), DATA_IN(26) => 
                           DATA_IN(26), DATA_IN(25) => DATA_IN(25), DATA_IN(24)
                           => DATA_IN(24), DATA_IN(23) => DATA_IN(23), 
                           DATA_IN(22) => DATA_IN(22), DATA_IN(21) => 
                           DATA_IN(21), DATA_IN(20) => DATA_IN(20), DATA_IN(19)
                           => DATA_IN(19), DATA_IN(18) => DATA_IN(18), 
                           DATA_IN(17) => DATA_IN(17), DATA_IN(16) => 
                           DATA_IN(16), DATA_IN(15) => DATA_IN(15), DATA_IN(14)
                           => DATA_IN(14), DATA_IN(13) => DATA_IN(13), 
                           DATA_IN(12) => DATA_IN(12), DATA_IN(11) => 
                           DATA_IN(11), DATA_IN(10) => DATA_IN(10), DATA_IN(9) 
                           => DATA_IN(9), DATA_IN(8) => DATA_IN(8), DATA_IN(7) 
                           => DATA_IN(7), DATA_IN(6) => DATA_IN(6), DATA_IN(5) 
                           => DATA_IN(5), DATA_IN(4) => DATA_IN(4), DATA_IN(3) 
                           => DATA_IN(3), DATA_IN(2) => DATA_IN(2), DATA_IN(1) 
                           => DATA_IN(1), DATA_IN(0) => DATA_IN(0), 
                           IRAM_OUT(31) => IRAM_OUT(31), IRAM_OUT(30) => 
                           IRAM_OUT(30), IRAM_OUT(29) => IRAM_OUT(29), 
                           IRAM_OUT(28) => IRAM_OUT(28), IRAM_OUT(27) => 
                           IRAM_OUT(27), IRAM_OUT(26) => IRAM_OUT(26), 
                           IRAM_OUT(25) => IRAM_OUT(25), IRAM_OUT(24) => 
                           IRAM_OUT(24), IRAM_OUT(23) => IRAM_OUT(23), 
                           IRAM_OUT(22) => IRAM_OUT(22), IRAM_OUT(21) => 
                           IRAM_OUT(21), IRAM_OUT(20) => IRAM_OUT(20), 
                           IRAM_OUT(19) => IRAM_OUT(19), IRAM_OUT(18) => 
                           IRAM_OUT(18), IRAM_OUT(17) => IRAM_OUT(17), 
                           IRAM_OUT(16) => IRAM_OUT(16), IRAM_OUT(15) => 
                           IRAM_OUT(15), IRAM_OUT(14) => IRAM_OUT(14), 
                           IRAM_OUT(13) => IRAM_OUT(13), IRAM_OUT(12) => 
                           IRAM_OUT(12), IRAM_OUT(11) => IRAM_OUT(11), 
                           IRAM_OUT(10) => IRAM_OUT(10), IRAM_OUT(9) => 
                           IRAM_OUT(9), IRAM_OUT(8) => IRAM_OUT(8), IRAM_OUT(7)
                           => IRAM_OUT(7), IRAM_OUT(6) => IRAM_OUT(6), 
                           IRAM_OUT(5) => IRAM_OUT(5), IRAM_OUT(4) => 
                           IRAM_OUT(4), IRAM_OUT(3) => IRAM_OUT(3), IRAM_OUT(2)
                           => IRAM_OUT(2), IRAM_OUT(1) => IRAM_OUT(1), 
                           IRAM_OUT(0) => IRAM_OUT(0), IRAM_ADDR(31) => 
                           IRAM_ADDR(31), IRAM_ADDR(30) => IRAM_ADDR(30), 
                           IRAM_ADDR(29) => IRAM_ADDR(29), IRAM_ADDR(28) => 
                           IRAM_ADDR(28), IRAM_ADDR(27) => IRAM_ADDR(27), 
                           IRAM_ADDR(26) => IRAM_ADDR(26), IRAM_ADDR(25) => 
                           IRAM_ADDR(25), IRAM_ADDR(24) => IRAM_ADDR(24), 
                           IRAM_ADDR(23) => IRAM_ADDR(23), IRAM_ADDR(22) => 
                           IRAM_ADDR(22), IRAM_ADDR(21) => IRAM_ADDR(21), 
                           IRAM_ADDR(20) => IRAM_ADDR(20), IRAM_ADDR(19) => 
                           IRAM_ADDR(19), IRAM_ADDR(18) => IRAM_ADDR(18), 
                           IRAM_ADDR(17) => IRAM_ADDR(17), IRAM_ADDR(16) => 
                           IRAM_ADDR(16), IRAM_ADDR(15) => IRAM_ADDR(15), 
                           IRAM_ADDR(14) => IRAM_ADDR(14), IRAM_ADDR(13) => 
                           IRAM_ADDR(13), IRAM_ADDR(12) => IRAM_ADDR(12), 
                           IRAM_ADDR(11) => IRAM_ADDR(11), IRAM_ADDR(10) => 
                           IRAM_ADDR(10), IRAM_ADDR(9) => IRAM_ADDR(9), 
                           IRAM_ADDR(8) => IRAM_ADDR(8), IRAM_ADDR(7) => 
                           IRAM_ADDR(7), IRAM_ADDR(6) => IRAM_ADDR(6), 
                           IRAM_ADDR(5) => IRAM_ADDR(5), IRAM_ADDR(4) => 
                           IRAM_ADDR(4), IRAM_ADDR(3) => IRAM_ADDR(3), 
                           IRAM_ADDR(2) => IRAM_ADDR(2), IRAM_ADDR(1) => 
                           IRAM_ADDR(1), IRAM_ADDR(0) => IRAM_ADDR(0), 
                           DATA_OUT(31) => DATA_OUT(31), DATA_OUT(30) => 
                           DATA_OUT(30), DATA_OUT(29) => DATA_OUT(29), 
                           DATA_OUT(28) => DATA_OUT(28), DATA_OUT(27) => 
                           DATA_OUT(27), DATA_OUT(26) => DATA_OUT(26), 
                           DATA_OUT(25) => DATA_OUT(25), DATA_OUT(24) => 
                           DATA_OUT(24), DATA_OUT(23) => DATA_OUT(23), 
                           DATA_OUT(22) => DATA_OUT(22), DATA_OUT(21) => 
                           DATA_OUT(21), DATA_OUT(20) => DATA_OUT(20), 
                           DATA_OUT(19) => DATA_OUT(19), DATA_OUT(18) => 
                           DATA_OUT(18), DATA_OUT(17) => DATA_OUT(17), 
                           DATA_OUT(16) => DATA_OUT(16), DATA_OUT(15) => 
                           DATA_OUT(15), DATA_OUT(14) => DATA_OUT(14), 
                           DATA_OUT(13) => DATA_OUT(13), DATA_OUT(12) => 
                           DATA_OUT(12), DATA_OUT(11) => DATA_OUT(11), 
                           DATA_OUT(10) => DATA_OUT(10), DATA_OUT(9) => 
                           DATA_OUT(9), DATA_OUT(8) => DATA_OUT(8), DATA_OUT(7)
                           => DATA_OUT(7), DATA_OUT(6) => DATA_OUT(6), 
                           DATA_OUT(5) => DATA_OUT(5), DATA_OUT(4) => 
                           DATA_OUT(4), DATA_OUT(3) => DATA_OUT(3), DATA_OUT(2)
                           => DATA_OUT(2), DATA_OUT(1) => DATA_OUT(1), 
                           DATA_OUT(0) => DATA_OUT(0), DATA_ADDR(31) => 
                           DATA_ADDR(31), DATA_ADDR(30) => DATA_ADDR(30), 
                           DATA_ADDR(29) => DATA_ADDR(29), DATA_ADDR(28) => 
                           DATA_ADDR(28), DATA_ADDR(27) => DATA_ADDR(27), 
                           DATA_ADDR(26) => DATA_ADDR(26), DATA_ADDR(25) => 
                           DATA_ADDR(25), DATA_ADDR(24) => DATA_ADDR(24), 
                           DATA_ADDR(23) => DATA_ADDR(23), DATA_ADDR(22) => 
                           DATA_ADDR(22), DATA_ADDR(21) => DATA_ADDR(21), 
                           DATA_ADDR(20) => DATA_ADDR(20), DATA_ADDR(19) => 
                           DATA_ADDR(19), DATA_ADDR(18) => DATA_ADDR(18), 
                           DATA_ADDR(17) => DATA_ADDR(17), DATA_ADDR(16) => 
                           DATA_ADDR(16), DATA_ADDR(15) => DATA_ADDR(15), 
                           DATA_ADDR(14) => DATA_ADDR(14), DATA_ADDR(13) => 
                           DATA_ADDR(13), DATA_ADDR(12) => DATA_ADDR(12), 
                           DATA_ADDR(11) => DATA_ADDR(11), DATA_ADDR(10) => 
                           DATA_ADDR(10), DATA_ADDR(9) => DATA_ADDR(9), 
                           DATA_ADDR(8) => DATA_ADDR(8), DATA_ADDR(7) => 
                           DATA_ADDR(7), DATA_ADDR(6) => DATA_ADDR(6), 
                           DATA_ADDR(5) => DATA_ADDR(5), DATA_ADDR(4) => 
                           DATA_ADDR(4), DATA_ADDR(3) => DATA_ADDR(3), 
                           DATA_ADDR(2) => DATA_ADDR(2), DATA_ADDR(1) => 
                           DATA_ADDR(1), DATA_ADDR(0) => DATA_ADDR(0), BMP => 
                           BMP_i, STALL(1) => STALL_CODE_1_port, STALL(0) => 
                           STALL_CODE_0_port, ID_EN => ID_EN_i, RF_RD => 
                           RF_RD_i, SIGND => SIGND_i, IMM_SEL => IMM_SEL_i, 
                           BPR_EN => BPR_EN_i, ALU_OPCODE(0) => 
                           ALU_OPCODE_i_0_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, EX_EN => n1, ALUA_SEL => n1, 
                           ALUB_SEL => n1, UCB_EN => UCB_EN_i, MEM_EN => 
                           MEM_EN_i, MEM_DATA_SEL => MEM_DATA_SEL_i, LD_SEL(2) 
                           => LD_SEL_i_2_port, LD_SEL(1) => LD_SEL_i_1_port, 
                           LD_SEL(0) => LD_SEL_i_0_port, ALR2_SEL => ALR2_SEL_i
                           , CWB_SEL(1) => CWB_SEL_i_1_port, CWB_SEL(0) => 
                           CWB_SEL_i_0_port, WB_SEL => WB_SEL_i, RF_WR => 
                           RF_WR_i, RF_MUX_SEL(1) => RF_MUX_SEL_i_1_port, 
                           RF_MUX_SEL(0) => RF_MUX_SEL_i_0_port);
   n1 <= '0';
   UCB_EN_i <= '0';
   BPR_EN_i <= '0';
   IMM_SEL_i <= '0';
   SIGND_i <= '0';
   RF_RD_i <= '0';
   ID_EN_i <= '0';

end SYN_dlx_rtl;
