library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.myTypes.all;
use work.constants.all;


entity TB_ALU is
end TB_ALU;

architecture TEST of TB_ALU is

    --component declaration
component ALU is
    generic (
      NBIT : integer := 32
    ); --# of signals the CMP can generate
    port (
      AluOpcode : in aluOp; -- input signals to select the operation to be performed by the ALU block
      A : in std_logic_vector(NBIT - 1 downto 0);
      B : in std_logic_vector(NBIT - 1 downto 0);
      Cin : in std_logic;
      ALU_out : out std_logic_vector(NBIT - 1 downto 0); -- 32-bit result produced from addition, subtraction, logical, etc.
      Cout : out std_logic; -- carry out generated by the adder/subtractor
      COND : out std_logic_vector(5 downto 0)
    );
  end component;

constant NBIT : integer := 32;

signal opcode_alu : aluOp;
signal carryin, carryout: std_logic;
signal psw : std_logic_vector(5 downto 0);
signal A_tb, B_tb, out_alu : std_logic_vector (NBIT-1 downto 0);

begin
	-- ALU instantiation
         DUT: ALU
         generic map (NBIT)
         port map (opcode_alu, A_tb, B_tb, carryin, out_alu, carryout, psw);

         --PROCESS FOR TESTING TEST
         carryin <= '0';
         ptest: process
         begin
             wait for 10 ns;

            
            opcode_alu <= OP_ADD;
            A_tb <= "00000000000000000000000000000101";
            B_tb <= "00000000000000000000000000000111";
            wait for 20 ns;
            
            opcode_alu <= OP_ADD;
            A_tb <= "00000000000000000000000000000101";
            B_tb <= "00000000000000000000000000000111";
            wait for 20 ns;

            opcode_alu <= OP_SUB;
            A_tb <= "00000000000000000000000000001101";
            B_tb <= "00000000000000000000000000010001";
            wait for 20 ns;

            opcode_alu <= OP_SUB;
            A_tb <= "00000000000000000000000000010001";
            B_tb <= "00000000000000000000000000010000";
            wait for 20 ns;

            opcode_alu <= OP_AND;
            A_tb <= "10001000100010001000100010001000";
            B_tb <= "10001000001000000001000000001111";
            wait for 20 ns;

            opcode_alu <= OP_XOR;
            A_tb <= "10001000100010001000100010001000";
            B_tb <= "10001000001000000001000000001111";
            wait for 20 ns;
            
            opcode_alu <= OP_NOR;
            A_tb <= "10001000100010001000100010001000";
            B_tb <= "10001000001000000001000000001111";
            wait for 20 ns;
            
            opcode_alu <= OP_XNOR;
            A_tb <= "10001000100010001000100010001000";
            B_tb <= "10001000001000000001000000001111";
            wait for 20 ns;

            opcode_alu <= OP_OR;
            A_tb <= "10001000100010001000100010001000";
            B_tb <= "10001000001000000001000000001111";
            wait for 20 ns;
            
            opcode_alu <= OP_NAND;
            A_tb <= "10001000100010001000100010001000";
            B_tb <= "10001000001000000001000000001111";
            wait for 20 ns;

            opcode_alu <= OP_SLL;
            A_tb <= "10001000100010001000100010001111";
            B_tb <= "00000000000000000000000000001010"; 
            wait for 20 ns;
         
            opcode_alu <= OP_SRA;
            A_tb <= "10001000100010001000100010001111"; 
            B_tb <= "00000000000000000000000000001010";
            wait for 20 ns;
            
            opcode_alu <= OP_SLL;
            A_tb <= "11111000100010001000100010001111";
            B_tb <= "00000000000000000000000000001010"; 
            wait for 20 ns;

            opcode_alu <= OP_SRL;
            A_tb <= "10001000100010001000100010001111";
            B_tb <= "00000000000000000000000000011000"; 
            wait for 20 ns;

            opcode_alu <= OP_CMP;
            A_tb <= "00000000000000000000000000001111";
            B_tb <= "00000000000000000000000000001011";
            wait for 20 ns;

            opcode_alu <= OP_CMP;
            A_tb <= "00000000000000000000000000000111";
            B_tb <= "00000000000000000000000000001011";
            wait for 20 ns;

            opcode_alu <= OP_CMP;
            A_tb <= "00000000000000000000000000001111";
            B_tb <= "00000000000000000000000000001111";
            wait for 20 ns;

            wait;

        end process ptest;
         
	
end TEST;
    
       