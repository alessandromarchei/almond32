library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.myTypes.all;
use WORK.constants.all;

--THIS MODULE IS THE TOP LEVEL ENTITY OF THE ARITHMETIC LOGIC UNIT

--INTERNALLY, IT CONTAINS AN ADDER (FOLLOWED BY A COMPARATOR), A LOGICAL UNIT THAT IS ABLE TO PERFORM
--OPERATIONS SUCH AS NOR, XOR, AND , NAND ..., A SHIFTER THAT IS EFFICIENTLY ABLE TO PERFORM LOGIC AND ARITHMETIC SHIFTS
--AND A PIPELINED MULTIPLIER BASED ON THE BOOTH'S ALGORITHM.

--IT CAN PERFORM ONE OPERATION AT A TIME BASED ON THE CONTROL SIGNAL RECEIVED BY THE CONTROL UNIT "ALUOPCODE"
--THANKS TO THIS, THE INTERNAL CONTROL UNIT OF THIS MODULE PROPERLY DRIVES THE ENABLE SIGNALS IN ORDER TO 
--TURN ON AND OFF THE EXECUTION UNITS AND HENCE SAVING DYNAMIC POWER WHEN THEY ARE NOT NEEDED.

entity ALU is
  generic (
    NBIT : integer := 32
  ); --# of signals the CMP can generate
  port (
    CLOCK : in std_logic;
    AluOpcode : in aluOp; -- input signals to select the operation to be performed by the ALU block
    A : in std_logic_vector(NBIT - 1 downto 0);
    B : in std_logic_vector(NBIT - 1 downto 0);
    Cin : in std_logic;
    ALU_out : out std_logic_vector(NBIT - 1 downto 0); -- 32-bit result produced from addition, subtraction, logical, etc.
    Cout : out std_logic; -- carry out generated by the adder/subtractor
    COND : out std_logic_vector(5 downto 0)   -- COND : [NE, E, GE, G, LE, L] (MSB left, LSB right)
  );
end ALU;

architecture BEHAVIORAL of ALU is
  component SHIFTER is
    port (
      data_in : in std_logic_vector(31 downto 0); -- Input data to be shifted
      R : in std_logic_vector(4 downto 0);
      conf : in std_logic_vector(1 downto 0);
      data_out : out std_logic_vector(31 downto 0) -- Shifted output data
    );
  end component;


  --OUTPUT MULTIPLEXER ABLE TO SELECT THE RIGHT OPERATION BASED ON THE ALUOPCODE
  component MUX4to1 is
    Generic (NBIT: integer := 32);
    Port (
      A, B, C, D: in std_logic_vector(NBIT-1 downto 0);
      SEL: in std_logic_vector(1 downto 0);
      Y: out std_logic_vector(NBIT-1 downto 0)
    );
  end component;

  component ADDER is
    generic (
      NBIT : integer := 32;
      NBIT_PER_BLOCK : integer := 4
    );
    port (
      A : in std_logic_vector(NBIT - 1 downto 0);
      B : in std_logic_vector(NBIT - 1 downto 0);
      ADD_SUB : in std_logic; -- Bit to select addition/subtraction
      Cin : in std_logic; -- Transparent in addition, fixed to 1 in subtraction
      S : out std_logic_vector(NBIT - 1 downto 0);
      Cout : out std_logic
    );
  end component;

  component LOGIC is
    generic (NBIT: integer := 32;
             N_SELECTOR: integer := 4
    );
    port (
        S   : in std_logic_vector (N_SELECTOR-1 downto 0); --Selector
        A, B: in std_logic_vector (NBIT-1 downto 0); --Operands
        O   : out std_logic_vector (NBIT-1 downto 0)--Logical evaluation
    );
end component;

  component AND2 is
    Port (
      A : in STD_LOGIC;
      B : in STD_LOGIC;
      Y : out STD_LOGIC
    );
  end component;

  component CMP is
    generic (
      NBIT : integer := 32
    );
    port (
      SUM : in std_logic_vector(NBIT - 1 downto 0); -- The adder receives A and B as inputs and generates SUM and Cout as outputs
      Cout : in std_logic;
      A_L_B : out std_logic; -- A < B   
      A_LE_B : out std_logic; -- A <= B
      A_G_B : out std_logic; -- A > B
      A_GE_B : out std_logic; -- A >= B
      A_E_B : out std_logic; -- A = B
      A_NE_B : out std_logic -- A /= B
    );
  end component;

  component MUL is
    Port (	CLOCK : in std_logic;
    A:	In	std_logic_vector(15 downto 0);
    B:	In	std_logic_vector(15 downto 0);
    Y:	Out	std_logic_vector(31 downto 0));
  end component;


  signal add_sub : std_logic := '0';    --ADDITION AS DEFAULT OPERATION
  signal cin_internal:  std_logic := '0'; 

  signal en_adder, en_cmp, en_logic, en_shifter, en_mul, c_out, en_adc: std_logic;
  signal mux_out : std_logic_vector(1 downto 0); -- to select the right output visible at the ALUOUT port
  -- MUX OUT : '0' ==> ADDER, '1' ==> LOGIC, '2' ==> SHIFTER.
  -- THE COMPARATOR IS ALWAYS VISIBLE AS OUTPUT PORT AT THE OUTPUT

  signal B_shifter : std_logic_vector(4 downto 0);
  -- internal signals connecting the input operands ports to the internal ports of the ALU-submodules
  signal A_adder, B_adder, out_adder, A_logic, B_logic, out_logic, A_shifter, out_shifter, in_cmp, out_mul : std_logic_vector(NBIT - 1 downto 0);
  signal conf : std_logic_vector(1 downto 0); -- used to convert the Aluopcode for the shift into valid signals for the SHIFTER SUB-MODULE

  -- signals for the logic
  signal logic_sel : std_logic_vector(3 downto 0);
  
  signal A_mul, B_mul : std_logic_vector(NBIT/2 - 1 downto 0);
begin

  --CONNECTING THE INTERNAL SIGNAL c_out to the EXTERNAL PORT COUT of the entire module
  Cout <= c_out;

  cin_internal <= Cin and en_adc;

  -- BUILDING THE ENABLE SIGNALS WITH THE PARALLEL SET OF 'AND' GATES
  --AS SPECIFIED ABOVE, THE ENABLE SIGNALS ARE NECESSARY IN ORDER TO SAVE POWER AND TURN OFF THE EXECUTION UNITS
  -- THAT ARE NOT USED AT THE MOMENT.

  -- ADDER ENABLE
  ENABLE_ADDER: for i in 0 to NBIT - 1 generate
    ADDER_A_i: AND2 port map(A(i), en_adder, A_adder(i));
    ADDER_B_i: AND2 port map(B(i), en_adder, B_adder(i));
  end generate;

  -- LOGIC ENABLE
  ENABLE_LOGIC: for i in 0 to NBIT - 1 generate
    LOGIC_A_i: AND2 port map(A(i), en_logic, A_logic(i));
    LOGIC_B_i: AND2 port map(B(i), en_logic, B_logic(i));
  end generate;

  -- SHIFTER ENABLE
  ENABLE_SHIFTER_A: for i in 0 to NBIT - 1 generate
    SHIFTER_A_i: AND2 port map(A(i), en_shifter, A_shifter(i));
  end generate;

  -- 5 BIT SELECTION FOR THE 2ND OPERAND OF THE SHIFTER
  ENABLE_SHIFTER_B: for i in 0 to 4 generate
    SHIFTER_B_i: AND2 port map(B(i), en_shifter, B_shifter(i));
  end generate;

  -- COMPARATOR ENABLE
  ENABLE_CMP_SUM: for i in 0 to NBIT - 1 generate
    SUM_i: AND2 port map(out_adder(i), en_cmp, in_cmp(i)); -- in_cmp IS THE INPUT OF THE COMPARATOR, BASED ON THE ENABLE SIGNAL ANDED WITH OUT_ADDER
  end generate;

  -- MULTIPLIER ENABLE
  ENABLE_MUL : for i in 0 to NBIT/2 - 1 generate
    MUL_A_i : AND2 port map(A(i), en_mul, A_mul(i));
    MUL_B_i : AND2 port map(B(i), en_mul, B_mul(i));
    end generate;

  -- INSTANTIATIONS OF THE COMPONENTS

  -- ADDER
  ADD: ADDER port map(A_adder, B_adder, add_sub, cin_internal, out_adder, c_out);

  -- SHIFTER
  SHIFT: SHIFTER port map(A_shifter, B_shifter, conf, out_shifter);

  -- LOGIC
  LOGICALS: LOGIC port map(logic_sel, A_logic, B_logic, out_logic);

  -- CMP
  COMPARATOR: CMP port map(in_cmp, c_out, COND(0), COND(1), COND(2), COND(3), COND(4), COND(5));

  --MUL
  MULTIPLIER : MUL generic map(16) port map(CLOCK, A_mul, B_mul, out_mul);

  -- OUTPUT MULTIPLEXER TO SELECT THE PROPER ALU OUTPUT
  -- MUX OUT : '0' ==> ADDER, '1' ==> LOGIC, '2' ==> SHIFTER, '3' ==> MULTIPLIER
  OUTPUT_SEL : MUX4TO1 generic map(32) port map(out_adder, out_logic, out_shifter, out_mul, mux_out, ALU_out);


  --ALU CONTROL UNIT : DRIVE THE CONTROL SIGNALS TO PROPERLY SELECT THE EXECUTION UNIT BASED ON THE REQUESTED OPERATION
  OPERATION: process(AluOpcode)
  begin
    case AluOpcode is

      when OP_MUL =>
        en_mul <= '1';
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '0';
        add_sub <= '0';
        mux_out <= "11";
        en_adc <= '0';

      when OP_ADD =>
        en_adder <= '1';
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '0';
        add_sub <= '0';
        mux_out <= "00";
        en_mul <= '0';
        en_adc <= '0';

      when OP_SUB =>
        en_adder <= '1';
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '0';
        add_sub <= '1';
        mux_out <= "00";
        en_mul <= '0';
        en_adc <= '0';

      when OP_ADC =>
        en_adder <= '1';
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '0';
        add_sub <= '0';
        mux_out <= "00";
        en_mul <= '0';
        en_adc <= '1';

      when OP_AND =>
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '1';
        en_shifter <= '0';
        add_sub <= '0';
        logic_sel <= "1000";
        mux_out <= "01";
        en_mul <= '0';
        en_adc <= '0';

      when OP_NAND =>
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '1';
        en_shifter <= '0';
        add_sub <= '0';
        logic_sel <= "0111";
        mux_out <= "01";
        en_mul <= '0';
        en_adc <= '0';

      when OP_OR =>
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '1';
        en_shifter <= '0';
        add_sub <= '0';
        logic_sel <= "1110";
        mux_out <= "01";
        en_mul <= '0';
        en_adc <= '0';

      when OP_NOR =>
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '1';
        en_shifter <= '0';
        add_sub <= '0';
        logic_sel <= "0001";
        mux_out <= "01";
        en_mul <= '0';
        en_adc <= '0';

      when OP_XOR =>
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '1';
        en_shifter <= '0';
        add_sub <= '0';
        logic_sel <= "0110";
        mux_out <= "01";
        en_mul <= '0';
        en_adc <= '0';

      when OP_XNOR =>
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '1';
        en_shifter <= '0';
        add_sub <= '0';
        logic_sel <= "1001";
        mux_out <= "01";
        en_mul <= '0';
        en_adc <= '0';

      when OP_SEQ =>
        en_adder <= '1'; -- SET EQUAL => USE COMPARATOR
        en_cmp <= '1';
        en_logic <= '0';
        en_shifter <= '0';
        add_sub <= '1';
        mux_out <= "00";
        en_mul <= '0';
        en_adc <= '0';
      
      when OP_SNE =>
      en_adder <= '1'; -- SET NOT EQUAL => USE COMPARATOR
      en_cmp <= '1';
      en_logic <= '0';
      en_shifter <= '0';
      add_sub <= '1';
      mux_out <= "00";
      en_mul <= '0';
      en_adc <= '0';

      when OP_SLT =>
      en_adder <= '1'; -- SET less than => USE COMPARATOR
      en_cmp <= '1';
      en_logic <= '0';
      en_shifter <= '0';
      add_sub <= '1';
      mux_out <= "00";
      en_mul <= '0';
      en_adc <= '0';

      when OP_SGT =>
      en_adder <= '1'; -- SET GREATER THAN => USE COMPARATOR
      en_cmp <= '1';
      en_logic <= '0';
      en_shifter <= '0';
      add_sub <= '1';
      mux_out <= "00";
      en_mul <= '0';
      en_adc <= '0';

      when OP_SLE =>
      en_adder <= '1'; -- SET LESS EQUAL => USE COMPARATOR
      en_cmp <= '1';
      en_logic <= '0';
      en_shifter <= '0';
      add_sub <= '1';
      mux_out <= "00";
      en_mul <= '0';
      en_adc <= '0';

      when OP_SGE =>
      en_adder <= '1'; -- SET GREATER EQUAL => USE COMPARATOR
      en_cmp <= '1';
      en_logic <= '0';
      en_shifter <= '0';
      add_sub <= '1';
      mux_out <= "00";
      en_mul <= '0';
      en_adc <= '0';

      when OP_SLL =>
        en_adder <= '0'; -- SHIFT LOGIC LEFT
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '1';
        add_sub <= '0';
        conf <= "00";
        mux_out <= "10";
        en_mul <= '0';
        en_adc <= '0';

      when OP_SRL =>
        en_adder <= '0'; -- SHIFT LOGIC RIGHT
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '1';
        add_sub <= '0';
        conf <= "01";
        mux_out <= "10";
        en_mul <= '0';
        en_adc <= '0';

      when OP_SRA =>
        en_adder <= '0'; -- SHIFT ARITHMETIC RIGHT
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '1';
        add_sub <= '0';
        conf <= "10";
        mux_out <= "10";
        en_mul <= '0';
        en_adc <= '0';

      when others => -- NOP case ==> TURN OFF ALL THE POSSIBLE COMPONENTS
        en_adder <= '0';
        en_cmp <= '0';
        en_logic <= '0';
        en_shifter <= '0';
        add_sub <= '0';
        conf <= "00";
        mux_out <= "00";
        en_mul <= '0';
        en_adc <= '0';
    end case;
  end process;

end architecture;
